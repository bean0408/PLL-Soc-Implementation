


timescale 1ns / 1ps
`default_nettype none


(*blackbox*)
module lvl_shifter(

		inout LVPWR,
		inout VGND,
		//inout VNB,
		//inout VPB,
		inout VPWR,
		
    		input A,
    
    		output X

);

