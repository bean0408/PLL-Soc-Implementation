# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  TIME NANOSECONDS 1 ;
  CAPACITANCE PICOFARADS 1 ;
  RESISTANCE OHMS 1 ;
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;

PROPERTYDEFINITIONS
  LAYER LEF58_TYPE STRING ;
END PROPERTYDEFINITIONS

# High voltage, single height
SITE unithv
  SYMMETRY Y ;
  CLASS CORE ;
  SIZE 0.48 BY 4.07 ;
END unithv

# High voltage, double height
SITE unithvdbl
  SYMMETRY Y ;
  CLASS CORE ;
  SIZE 0.48 BY 8.14 ;
END unithvdbl

LAYER nwell
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE NWELL ;" ;
END nwell

LAYER pwell
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE NWELL ;" ;
END pwell

LAYER li1
  TYPE ROUTING ;
  DIRECTION VERTICAL ;

  PITCH 0.48 ;
  MINWIDTH 0.17 ;

  WIDTH 0.17 ;          # LI 1
  # SPACING  0.17 ;     # LI 2
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 0.17 ;
  AREA 0.0561 ;         # LI 6
  THICKNESS 0.1 ;
  EDGECAPACITANCE 40.697E-6 ;
  CAPACITANCE CPERSQDIST 36.9866E-6 ;
  RESISTANCE RPERSQ 12.2 ;

  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 75 ) ( 0.0125 75 ) ( 0.0225 85.125 ) ( 22.5 10200 ) ) ;
END li1

LAYER mcon
  TYPE CUT ;

  WIDTH 0.17 ;                # Mcon 1
  SPACING 0.19 ;              # Mcon 2
  ENCLOSURE BELOW 0 0 ;       # Mcon 4
  ENCLOSURE ABOVE 0.03 0.06 ; # Met1 4 / Met1 5

  ANTENNADIFFAREARATIO PWL ( ( 0 3 ) ( 0.0125 3 ) ( 0.0225 3.405 ) ( 22.5 408 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.36 ; # mA per via Iavg_max at Tj = 90oC

END mcon

LAYER met1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;

  PITCH 0.37 ;
  MINENCLOSEDAREA 0.14 ;
  MINWIDTH 0.14 ;

  WIDTH 0.14 ;                     # Met1 1
  # SPACING 0.14 ;                 # Met1 2
  # SPACING 0.28 RANGE 3.001 100 ; # Met1 3b
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 0.14
     WIDTH 3 0.28 ;
  AREA 0.083 ;                     # Met1 6
  THICKNESS 0.35 ;

  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;

  EDGECAPACITANCE 40.567E-6 ;
  CAPACITANCE CPERSQDIST 25.7784E-6 ;
  DCCURRENTDENSITY AVERAGE 2.8 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 6.1 ; # mA/um Irms_max at Tj = 90oC

  RESISTANCE RPERSQ 0.125 ;
END met1

LAYER via
  TYPE CUT ;
  WIDTH 0.15 ;                  # Via 1a
  SPACING 0.17 ;                # Via 2
  ENCLOSURE BELOW 0.055 0.085 ; # Via 4a / Via 5a
  ENCLOSURE ABOVE 0.055 0.085 ; # Met2 4 / Met2 5

  ANTENNADIFFAREARATIO PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.29 ; # mA per via Iavg_max at Tj = 90oC
END via

LAYER met2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;

  PITCH 0.48 ;
  MINENCLOSEDAREA 0.14 ;
  MINWIDTH 0.14 ;

  WIDTH 0.14 ;                        # Met2 1
  # SPACING  0.14 ;                   # Met2 2
  # SPACING  0.28 RANGE 3.001 100 ;   # Met2 3b
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 0.14
     WIDTH 3 0.28 ;
  AREA 0.0676 ;                       # Met2 6
  THICKNESS 0.35 ;

  EDGECAPACITANCE 37.759E-6 ;
  CAPACITANCE CPERSQDIST 16.9423E-6 ;
  RESISTANCE RPERSQ 0.125 ;
  DCCURRENTDENSITY AVERAGE 2.8 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 6.1 ; # mA/um Irms_max at Tj = 90oC
  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;
END met2

# ******** Layer via2, type routing, number 44 **************
LAYER via2
  TYPE CUT ;
  WIDTH 0.2 ;                   # Via2 1
  SPACING 0.2 ;                 # Via2 2
  ENCLOSURE BELOW 0.04 0.085 ;  # Via2 4
  ENCLOSURE ABOVE 0.065 0.065 ; # Met3 4
  ANTENNADIFFAREARATIO PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.48 ; # mA per via Iavg_max at Tj = 90oC
END via2

LAYER met3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;

  PITCH 0.74 ;
  MINWIDTH 0.3 ;

  WIDTH 0.3 ;              # Met3 1
  # SPACING 0.3 ;          # Met3 2
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 0.3
     WIDTH 3 0.4 ;
  AREA 0.24 ;              # Met3 6
  THICKNESS 0.8 ;

  EDGECAPACITANCE 40.989E-6 ;
  CAPACITANCE CPERSQDIST 12.3729E-6 ;
  RESISTANCE RPERSQ 0.047 ;
  DCCURRENTDENSITY AVERAGE 6.8 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 14.9 ; # mA/um Irms_max at Tj = 90oC

  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;
END met3

LAYER via3
  TYPE CUT ;
  WIDTH 0.2 ;                   # Via3 1
  SPACING 0.2 ;                 # Via3 2
  ENCLOSURE BELOW 0.06 0.09 ;   # Via3 4 / Via3 5
  ENCLOSURE ABOVE 0.065 0.065 ; # Met4 3
  ANTENNADIFFAREARATIO PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
  DCCURRENTDENSITY AVERAGE 0.48 ; # mA per via Iavg_max at Tj = 90oC
END via3

LAYER met4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;

  PITCH 0.96 ;
  MINWIDTH 0.3 ;

  WIDTH 0.3 ;             # Met4 1
  # SPACING  0.3 ;             # Met4 2
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 0.3
     WIDTH 3 0.4 ;
  AREA 0.24 ;              # Met4 4a

  THICKNESS 0.8 ;

  EDGECAPACITANCE 36.676E-6 ;
  CAPACITANCE CPERSQDIST 8.41537E-6 ;
  RESISTANCE RPERSQ 0.047 ;
  DCCURRENTDENSITY AVERAGE 6.8 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 14.9 ; # mA/um Irms_max at Tj = 90oC

  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;
END met4

LAYER via4
  TYPE CUT ;

  WIDTH 0.8 ;                 # Via4 1
  SPACING 0.8 ;               # Via4 2
  ENCLOSURE BELOW 0.19 0.19 ; # Via4 4
  ENCLOSURE ABOVE 0.31 0.31 ; # Met5 3
  ANTENNADIFFAREARATIO PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
  DCCURRENTDENSITY AVERAGE 2.49 ; # mA per via Iavg_max at Tj = 90oC
END via4

LAYER met5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;

  PITCH 3.33 ;
  MINWIDTH 1.6 ;

  WIDTH 1.6 ;            # Met5 1
  #SPACING  1.6 ;        # Met5 2
  SPACINGTABLE
     PARALLELRUNLENGTH 0
     WIDTH 0 1.6 ;
  AREA 4 ;               # Met5 4

  THICKNESS 1.2 ;

  EDGECAPACITANCE 38.851E-6 ;
  CAPACITANCE CPERSQDIST 6.32063E-6 ;
  RESISTANCE RPERSQ 0.0285 ;
  DCCURRENTDENSITY AVERAGE 10.17 ; # mA/um Iavg_max at Tj = 90oC
  ACCURRENTDENSITY RMS 22.34 ; # mA/um Irms_max at Tj = 90oC

  ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;
END met5


### Routing via cells section   ###
# Plus via rule, metals are along the prefered direction
VIA L1M1_PR DEFAULT
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER li1 ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
  RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIARULE L1M1_PR GENERATE
  LAYER li1 ;
  ENCLOSURE 0 0 ;
  LAYER met1 ;
  ENCLOSURE 0.06 0.03 ;
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  SPACING 0.36 BY 0.36 ;
END L1M1_PR

# Plus via rule, metals are along the non prefered direction
VIA L1M1_PR_R DEFAULT
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER li1 ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
  RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIARULE L1M1_PR_R GENERATE
  LAYER li1 ;
  ENCLOSURE 0 0 ;
  LAYER met1 ;
  ENCLOSURE 0.03 0.06 ;
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  SPACING 0.36 BY 0.36 ;
END L1M1_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA L1M1_PR_M DEFAULT
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER li1 ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
  RECT -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIARULE L1M1_PR_M GENERATE
  LAYER li1 ;
  ENCLOSURE 0 0 ;
  LAYER met1 ;
  ENCLOSURE 0.03 0.06 ;
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  SPACING 0.36 BY 0.36 ;
END L1M1_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA L1M1_PR_MR DEFAULT
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER li1 ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
  RECT -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIARULE L1M1_PR_MR GENERATE
  LAYER li1 ;
  ENCLOSURE 0 0 ;
  LAYER met1 ;
  ENCLOSURE 0.06 0.03 ;
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  SPACING 0.36 BY 0.36 ;
END L1M1_PR_MR

# Centered via rule, we really do not want to use it
VIA L1M1_PR_C DEFAULT
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER li1 ;
  RECT -0.085 -0.085 0.085 0.085 ;
  LAYER met1 ;
  RECT -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIARULE L1M1_PR_C GENERATE
  LAYER li1 ;
  ENCLOSURE 0 0 ;
  LAYER met1 ;
  ENCLOSURE 0.06 0.06 ;
  LAYER mcon ;
  RECT -0.085 -0.085 0.085 0.085 ;
  SPACING 0.36 BY 0.36 ;
END L1M1_PR_C

# Plus via rule, metals are along the prefered direction
VIA M1M2_PR DEFAULT
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met1 ;
  RECT -0.16 -0.13 0.16 0.13 ;
  LAYER met2 ;
  RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIARULE M1M2_PR GENERATE
  LAYER met1 ;
  ENCLOSURE 0.085 0.055 ;
  LAYER met2 ;
  ENCLOSURE 0.055 0.085 ;
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  SPACING 0.32 BY 0.32 ;
END M1M2_PR

# Plus via rule, metals are along the non prefered direction
VIA M1M2_PR_R DEFAULT
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met1 ;
  RECT -0.13 -0.16 0.13 0.16 ;
  LAYER met2 ;
  RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIARULE M1M2_PR_R GENERATE
  LAYER met1 ;
  ENCLOSURE 0.055 0.085 ;
  LAYER met2 ;
  ENCLOSURE 0.085 0.055 ;
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  SPACING 0.32 BY 0.32 ;
END M1M2_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA M1M2_PR_M DEFAULT
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met1 ;
  RECT -0.16 -0.13 0.16 0.13 ;
  LAYER met2 ;
  RECT -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIARULE M1M2_PR_M GENERATE
  LAYER met1 ;
  ENCLOSURE 0.085 0.055 ;
  LAYER met2 ;
  ENCLOSURE 0.085 0.055 ;
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  SPACING 0.32 BY 0.32 ;
END M1M2_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA M1M2_PR_MR DEFAULT
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met1 ;
  RECT -0.13 -0.16 0.13 0.16 ;
  LAYER met2 ;
  RECT -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIARULE M1M2_PR_MR GENERATE
  LAYER met1 ;
  ENCLOSURE 0.055 0.085 ;
  LAYER met2 ;
  ENCLOSURE 0.055 0.085 ;
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  SPACING 0.32 BY 0.32 ;
END M1M2_PR_MR

# Centered via rule, we really do not want to use it
VIA M1M2_PR_C DEFAULT
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  LAYER met1 ;
  RECT -0.16 -0.16 0.16 0.16 ;
  LAYER met2 ;
  RECT -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIARULE M1M2_PR_C GENERATE
  LAYER met1 ;
  ENCLOSURE 0.085 0.085 ;
  LAYER met2 ;
  ENCLOSURE 0.085 0.085 ;
  LAYER via ;
  RECT -0.075 -0.075 0.075 0.075 ;
  SPACING 0.32 BY 0.32 ;
END M1M2_PR_C

# Plus via rule, metals are along the prefered direction
VIA M2M3_PR DEFAULT
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met2 ;
  RECT -0.14 -0.185 0.14 0.185 ;
  LAYER met3 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIARULE M2M3_PR GENERATE
  LAYER met2 ;
  ENCLOSURE 0.04 0.085 ;
  LAYER met3 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M2M3_PR

# Plus via rule, metals are along the non prefered direction
VIA M2M3_PR_R DEFAULT
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met2 ;
  RECT -0.185 -0.14 0.185 0.14 ;
  LAYER met3 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIARULE M2M3_PR_R GENERATE
  LAYER met2 ;
  ENCLOSURE 0.085 0.04 ;
  LAYER met3 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M2M3_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA M2M3_PR_M DEFAULT
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met2 ;
  RECT -0.14 -0.185 0.14 0.185 ;
  LAYER met3 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIARULE M2M3_PR_M GENERATE
  LAYER met2 ;
  ENCLOSURE 0.04 0.085 ;
  LAYER met3 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M2M3_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA M2M3_PR_MR DEFAULT
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met2 ;
  RECT -0.185 -0.14 0.185 0.14 ;
  LAYER met3 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIARULE M2M3_PR_MR GENERATE
  LAYER met2 ;
  ENCLOSURE 0.085 0.04 ;
  LAYER met3 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M2M3_PR_MR

# Centered via rule, we really do not want to use it
VIA M2M3_PR_C DEFAULT
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met2 ;
  RECT -0.185 -0.185 0.185 0.185 ;
  LAYER met3 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIARULE M2M3_PR_C GENERATE
  LAYER met2 ;
  ENCLOSURE 0.085 0.085 ;
  LAYER met3 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via2 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M2M3_PR_C

# Plus via rule, metals are along the prefered direction
VIA M3M4_PR DEFAULT
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
  RECT -0.19 -0.16 0.19 0.16 ;
  LAYER met4 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIARULE M3M4_PR GENERATE
  LAYER met3 ;
  ENCLOSURE 0.09 0.06 ;
  LAYER met4 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M3M4_PR

# Plus via rule, metals are along the non prefered direction
VIA M3M4_PR_R DEFAULT
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
  RECT -0.16 -0.19 0.16 0.19 ;
  LAYER met4 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIARULE M3M4_PR_R GENERATE
  LAYER met3 ;
  ENCLOSURE 0.06 0.09 ;
  LAYER met4 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M3M4_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA M3M4_PR_M DEFAULT
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
  RECT -0.19 -0.16 0.19 0.16 ;
  LAYER met4 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIARULE M3M4_PR_M GENERATE
  LAYER met3 ;
  ENCLOSURE 0.09 0.06 ;
  LAYER met4 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M3M4_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA M3M4_PR_MR DEFAULT
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
  RECT -0.16 -0.19 0.16 0.19 ;
  LAYER met4 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIARULE M3M4_PR_MR GENERATE
  LAYER met3 ;
  ENCLOSURE 0.06 0.09 ;
  LAYER met4 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M3M4_PR_MR

# Centered via rule, we really do not want to use it
VIA M3M4_PR_C DEFAULT
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  LAYER met3 ;
  RECT -0.19 -0.19 0.19 0.19 ;
  LAYER met4 ;
  RECT -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIARULE M3M4_PR_C GENERATE
  LAYER met3 ;
  ENCLOSURE 0.09 0.09 ;
  LAYER met4 ;
  ENCLOSURE 0.065 0.065 ;
  LAYER via3 ;
  RECT -0.1 -0.1 0.1 0.1 ;
  SPACING 0.4 BY 0.4 ;
END M3M4_PR_C

# Plus via rule, metals are along the prefered direction
VIA M4M5_PR DEFAULT
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met4 ;
  RECT -0.59 -0.59 0.59 0.59 ;
  LAYER met5 ;
  RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIARULE M4M5_PR GENERATE
  LAYER met4 ;
  ENCLOSURE 0.19 0.19 ;
  LAYER met5 ;
  ENCLOSURE 0.31 0.31 ;
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  SPACING 1.6 BY 1.6 ;
END M4M5_PR

# Plus via rule, metals are along the non prefered direction
VIA M4M5_PR_R DEFAULT
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met4 ;
  RECT -0.59 -0.59 0.59 0.59 ;
  LAYER met5 ;
  RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIARULE M4M5_PR_R GENERATE
  LAYER met4 ;
  ENCLOSURE 0.19 0.19 ;
  LAYER met5 ;
  ENCLOSURE 0.31 0.31 ;
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  SPACING 1.6 BY 1.6 ;
END M4M5_PR_R

# Minus via rule, lower layer metal is along prefered direction
VIA M4M5_PR_M DEFAULT
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met4 ;
  RECT -0.59 -0.59 0.59 0.59 ;
  LAYER met5 ;
  RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIARULE M4M5_PR_M GENERATE
  LAYER met4 ;
  ENCLOSURE 0.19 0.19 ;
  LAYER met5 ;
  ENCLOSURE 0.31 0.31 ;
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  SPACING 1.6 BY 1.6 ;
END M4M5_PR_M

# Minus via rule, upper layer metal is along prefered direction
VIA M4M5_PR_MR DEFAULT
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met4 ;
  RECT -0.59 -0.59 0.59 0.59 ;
  LAYER met5 ;
  RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIARULE M4M5_PR_MR GENERATE
  LAYER met4 ;
  ENCLOSURE 0.19 0.19 ;
  LAYER met5 ;
  ENCLOSURE 0.31 0.31 ;
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  SPACING 1.6 BY 1.6 ;
END M4M5_PR_MR

# Centered via rule, we really do not want to use it
VIA M4M5_PR_C DEFAULT
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  LAYER met4 ;
  RECT -0.59 -0.59 0.59 0.59 ;
  LAYER met5 ;
  RECT -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

VIARULE M4M5_PR_C GENERATE
  LAYER met4 ;
  ENCLOSURE 0.19 0.19 ;
  LAYER met5 ;
  ENCLOSURE 0.31 0.31 ;
  LAYER via4 ;
  RECT -0.4 -0.4 0.4 0.4 ;
  SPACING 1.6 BY 1.6 ;
END M4M5_PR_C
###  end of single via cells   ###


MACRO sky130_fd_sc_hvl__inv_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__inv_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.440000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.550000 0.835000 1.935000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.641250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.960000 2.175000 1.345000 3.755000 ;
        RECT 1.015000 0.495000 1.345000 2.175000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 1.440000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 1.440000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 1.440000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 1.440000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 1.770000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 1.440000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.440000 0.085000 ;
      RECT 0.000000  3.985000 1.440000 4.155000 ;
      RECT 0.090000  0.365000 0.680000 1.325000 ;
      RECT 0.090000  2.175000 0.680000 3.755000 ;
    LAYER mcon ;
      RECT 0.120000  0.395000 0.290000 0.565000 ;
      RECT 0.120000  3.505000 0.290000 3.675000 ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.480000  0.395000 0.650000 0.565000 ;
      RECT 0.480000  3.505000 0.650000 3.675000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
  END
END sky130_fd_sc_hvl__inv_1
MACRO sky130_fd_sc_hvl__inv_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__inv_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  4.500000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.580000 2.835000 1.750000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  1.260000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.040000 0.495000 1.290000 1.230000 ;
        RECT 1.040000 1.230000 3.185000 1.400000 ;
        RECT 1.040000 1.930000 3.715000 2.100000 ;
        RECT 1.040000 2.100000 1.370000 3.755000 ;
        RECT 2.600000 0.495000 3.185000 1.230000 ;
        RECT 2.680000 2.100000 2.930000 3.755000 ;
        RECT 3.015000 1.400000 3.185000 1.550000 ;
        RECT 3.015000 1.550000 3.715000 1.930000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 3.840000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 3.840000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 3.840000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 3.840000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 4.170000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 3.840000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.985000 3.840000 4.155000 ;
      RECT 0.090000  0.365000 0.680000 1.325000 ;
      RECT 0.090000  2.175000 0.680000 3.755000 ;
      RECT 1.470000  0.365000 2.420000 1.050000 ;
      RECT 1.550000  2.280000 2.500000 3.755000 ;
      RECT 3.120000  2.280000 3.710000 3.755000 ;
      RECT 3.380000  0.365000 3.710000 1.325000 ;
    LAYER mcon ;
      RECT 0.120000  0.395000 0.290000 0.565000 ;
      RECT 0.120000  3.505000 0.290000 3.675000 ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.480000  0.395000 0.650000 0.565000 ;
      RECT 0.480000  3.505000 0.650000 3.675000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.500000  0.395000 1.670000 0.565000 ;
      RECT 1.580000  3.505000 1.750000 3.675000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.860000  0.395000 2.030000 0.565000 ;
      RECT 1.940000  3.505000 2.110000 3.675000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.220000  0.395000 2.390000 0.565000 ;
      RECT 2.300000  3.505000 2.470000 3.675000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
      RECT 3.150000  3.505000 3.320000 3.675000 ;
      RECT 3.410000  0.395000 3.580000 0.565000 ;
      RECT 3.510000  3.505000 3.680000 3.675000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.985000 3.685000 4.155000 ;
  END
END sky130_fd_sc_hvl__inv_4
MACRO sky130_fd_sc_hvl__inv_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__inv_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.400000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  2.250000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.550000 1.070000 1.880000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.630000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.200000 0.540000 1.795000 1.370000 ;
        RECT 1.240000 1.610000 1.795000 1.780000 ;
        RECT 1.240000 1.780000 1.490000 3.755000 ;
        RECT 1.565000 1.370000 1.795000 1.610000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 2.400000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 2.400000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 2.400000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 2.400000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 2.730000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 2.400000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.400000 0.085000 ;
      RECT 0.000000  3.985000 2.400000 4.155000 ;
      RECT 0.090000  0.365000 1.020000 1.370000 ;
      RECT 0.110000  2.175000 1.060000 3.755000 ;
      RECT 1.680000  2.175000 2.270000 3.755000 ;
      RECT 1.980000  0.365000 2.310000 1.370000 ;
    LAYER mcon ;
      RECT 0.110000  0.395000 0.280000 0.565000 ;
      RECT 0.140000  3.505000 0.310000 3.675000 ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.470000  0.395000 0.640000 0.565000 ;
      RECT 0.500000  3.505000 0.670000 3.675000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.830000  0.395000 1.000000 0.565000 ;
      RECT 0.860000  3.505000 1.030000 3.675000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.710000  3.505000 1.880000 3.675000 ;
      RECT 2.010000  0.395000 2.180000 0.565000 ;
      RECT 2.070000  3.505000 2.240000 3.675000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
  END
END sky130_fd_sc_hvl__inv_2
MACRO sky130_fd_sc_hvl__inv_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__inv_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.44000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  18.00000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  1.535000 1.550000  2.185000 1.580000 ;
        RECT  1.535000 1.580000 11.535000 1.750000 ;
        RECT  1.535000 1.750000  2.185000 1.780000 ;
        RECT  3.085000 1.550000  3.735000 1.580000 ;
        RECT  3.085000 1.750000  3.735000 1.780000 ;
        RECT  4.645000 1.550000  5.295000 1.580000 ;
        RECT  4.645000 1.750000  5.295000 1.780000 ;
        RECT  6.205000 1.550000  6.855000 1.580000 ;
        RECT  6.205000 1.750000  6.855000 1.780000 ;
        RECT  7.765000 1.550000  8.415000 1.580000 ;
        RECT  7.765000 1.750000  8.415000 1.780000 ;
        RECT  9.325000 1.550000  9.975000 1.580000 ;
        RECT  9.325000 1.750000  9.975000 1.780000 ;
        RECT 10.885000 1.550000 11.535000 1.580000 ;
        RECT 10.885000 1.750000 11.535000 1.780000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  5.040000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  0.925000 2.290000  1.215000 2.320000 ;
        RECT  0.925000 2.320000 12.135000 2.490000 ;
        RECT  0.925000 2.490000  1.215000 2.520000 ;
        RECT  2.485000 2.290000  2.775000 2.320000 ;
        RECT  2.485000 2.490000  2.775000 2.520000 ;
        RECT  4.045000 2.290000  4.335000 2.320000 ;
        RECT  4.045000 2.490000  4.335000 2.520000 ;
        RECT  5.605000 2.290000  5.895000 2.320000 ;
        RECT  5.605000 2.490000  5.895000 2.520000 ;
        RECT  7.165000 2.290000  7.455000 2.320000 ;
        RECT  7.165000 2.490000  7.455000 2.520000 ;
        RECT  8.725000 2.290000  9.015000 2.320000 ;
        RECT  8.725000 2.490000  9.015000 2.520000 ;
        RECT 10.285000 2.290000 10.575000 2.320000 ;
        RECT 10.285000 2.490000 10.575000 2.520000 ;
        RECT 11.845000 2.290000 12.135000 2.320000 ;
        RECT 11.845000 2.490000 12.135000 2.520000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 13.440000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 13.440000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 13.440000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 13.440000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 13.770000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 13.440000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.440000 0.085000 ;
      RECT  0.000000  3.985000 13.440000 4.155000 ;
      RECT  0.095000  0.375000  0.630000 1.475000 ;
      RECT  0.125000  2.175000  0.655000 3.755000 ;
      RECT  0.900000  0.795000  1.230000 3.755000 ;
      RECT  1.400000  0.375000  2.290000 1.395000 ;
      RECT  1.400000  1.565000  2.290000 1.895000 ;
      RECT  1.400000  2.175000  2.290000 3.755000 ;
      RECT  2.460000  0.795000  2.790000 3.755000 ;
      RECT  2.960000  0.375000  3.850000 1.395000 ;
      RECT  2.960000  1.565000  3.850000 1.895000 ;
      RECT  2.960000  2.175000  3.850000 3.755000 ;
      RECT  4.020000  0.795000  4.350000 3.755000 ;
      RECT  4.520000  0.375000  5.410000 1.395000 ;
      RECT  4.520000  1.565000  5.410000 1.895000 ;
      RECT  4.520000  2.175000  5.410000 3.755000 ;
      RECT  5.580000  0.795000  5.910000 3.755000 ;
      RECT  6.080000  0.375000  6.970000 1.395000 ;
      RECT  6.080000  1.565000  6.970000 1.895000 ;
      RECT  6.080000  2.175000  6.970000 3.755000 ;
      RECT  7.140000  0.795000  7.470000 3.755000 ;
      RECT  7.640000  0.375000  8.530000 1.395000 ;
      RECT  7.640000  1.565000  8.530000 1.895000 ;
      RECT  7.640000  2.175000  8.530000 3.755000 ;
      RECT  8.700000  0.795000  9.030000 3.755000 ;
      RECT  9.200000  0.375000 10.090000 1.395000 ;
      RECT  9.200000  1.565000 10.090000 1.895000 ;
      RECT  9.200000  2.175000 10.090000 3.755000 ;
      RECT 10.260000  0.795000 10.590000 3.755000 ;
      RECT 10.760000  0.375000 11.650000 1.395000 ;
      RECT 10.760000  1.565000 11.650000 1.895000 ;
      RECT 10.760000  2.175000 11.650000 3.755000 ;
      RECT 11.820000  0.795000 12.150000 3.755000 ;
      RECT 12.320000  0.375000 12.935000 1.395000 ;
      RECT 12.320000  2.175000 12.935000 3.675000 ;
    LAYER mcon ;
      RECT  0.095000  0.425000  0.265000 0.595000 ;
      RECT  0.125000  3.475000  0.295000 3.645000 ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.985000  0.325000 4.155000 ;
      RECT  0.455000  0.425000  0.625000 0.595000 ;
      RECT  0.485000  3.475000  0.655000 3.645000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.985000  0.805000 4.155000 ;
      RECT  0.985000  2.320000  1.155000 2.490000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.985000  1.285000 4.155000 ;
      RECT  1.400000  0.425000  1.570000 0.595000 ;
      RECT  1.400000  3.475000  1.570000 3.645000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  1.580000  1.765000 1.750000 ;
      RECT  1.595000  3.985000  1.765000 4.155000 ;
      RECT  1.760000  0.425000  1.930000 0.595000 ;
      RECT  1.760000  3.475000  1.930000 3.645000 ;
      RECT  1.955000  1.580000  2.125000 1.750000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.985000  2.245000 4.155000 ;
      RECT  2.120000  0.425000  2.290000 0.595000 ;
      RECT  2.120000  3.475000  2.290000 3.645000 ;
      RECT  2.545000  2.320000  2.715000 2.490000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.985000  2.725000 4.155000 ;
      RECT  2.960000  0.425000  3.130000 0.595000 ;
      RECT  2.960000  3.475000  3.130000 3.645000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.985000  3.205000 4.155000 ;
      RECT  3.145000  1.580000  3.315000 1.750000 ;
      RECT  3.320000  0.425000  3.490000 0.595000 ;
      RECT  3.320000  3.475000  3.490000 3.645000 ;
      RECT  3.505000  1.580000  3.675000 1.750000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.985000  3.685000 4.155000 ;
      RECT  3.680000  0.425000  3.850000 0.595000 ;
      RECT  3.680000  3.475000  3.850000 3.645000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.985000  4.165000 4.155000 ;
      RECT  4.105000  2.320000  4.275000 2.490000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.985000  4.645000 4.155000 ;
      RECT  4.520000  0.425000  4.690000 0.595000 ;
      RECT  4.520000  3.475000  4.690000 3.645000 ;
      RECT  4.705000  1.580000  4.875000 1.750000 ;
      RECT  4.880000  0.425000  5.050000 0.595000 ;
      RECT  4.880000  3.475000  5.050000 3.645000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.985000  5.125000 4.155000 ;
      RECT  5.065000  1.580000  5.235000 1.750000 ;
      RECT  5.240000  0.425000  5.410000 0.595000 ;
      RECT  5.240000  3.475000  5.410000 3.645000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.985000  5.605000 4.155000 ;
      RECT  5.665000  2.320000  5.835000 2.490000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.985000  6.085000 4.155000 ;
      RECT  6.080000  0.425000  6.250000 0.595000 ;
      RECT  6.080000  3.475000  6.250000 3.645000 ;
      RECT  6.265000  1.580000  6.435000 1.750000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.985000  6.565000 4.155000 ;
      RECT  6.440000  0.425000  6.610000 0.595000 ;
      RECT  6.440000  3.475000  6.610000 3.645000 ;
      RECT  6.625000  1.580000  6.795000 1.750000 ;
      RECT  6.800000  0.425000  6.970000 0.595000 ;
      RECT  6.800000  3.475000  6.970000 3.645000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.985000  7.045000 4.155000 ;
      RECT  7.225000  2.320000  7.395000 2.490000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.985000  7.525000 4.155000 ;
      RECT  7.640000  0.425000  7.810000 0.595000 ;
      RECT  7.640000  3.475000  7.810000 3.645000 ;
      RECT  7.825000  1.580000  7.995000 1.750000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.985000  8.005000 4.155000 ;
      RECT  8.000000  0.425000  8.170000 0.595000 ;
      RECT  8.000000  3.475000  8.170000 3.645000 ;
      RECT  8.185000  1.580000  8.355000 1.750000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.985000  8.485000 4.155000 ;
      RECT  8.360000  0.425000  8.530000 0.595000 ;
      RECT  8.360000  3.475000  8.530000 3.645000 ;
      RECT  8.785000  2.320000  8.955000 2.490000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.985000  8.965000 4.155000 ;
      RECT  9.200000  0.425000  9.370000 0.595000 ;
      RECT  9.200000  3.475000  9.370000 3.645000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.985000  9.445000 4.155000 ;
      RECT  9.385000  1.580000  9.555000 1.750000 ;
      RECT  9.560000  0.425000  9.730000 0.595000 ;
      RECT  9.560000  3.475000  9.730000 3.645000 ;
      RECT  9.745000  1.580000  9.915000 1.750000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.985000  9.925000 4.155000 ;
      RECT  9.920000  0.425000 10.090000 0.595000 ;
      RECT  9.920000  3.475000 10.090000 3.645000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.985000 10.405000 4.155000 ;
      RECT 10.345000  2.320000 10.515000 2.490000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.985000 10.885000 4.155000 ;
      RECT 10.760000  0.425000 10.930000 0.595000 ;
      RECT 10.760000  3.475000 10.930000 3.645000 ;
      RECT 10.945000  1.580000 11.115000 1.750000 ;
      RECT 11.120000  0.425000 11.290000 0.595000 ;
      RECT 11.120000  3.475000 11.290000 3.645000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.985000 11.365000 4.155000 ;
      RECT 11.305000  1.580000 11.475000 1.750000 ;
      RECT 11.480000  0.425000 11.650000 0.595000 ;
      RECT 11.480000  3.475000 11.650000 3.645000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.985000 11.845000 4.155000 ;
      RECT 11.905000  2.320000 12.075000 2.490000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.985000 12.325000 4.155000 ;
      RECT 12.365000  0.425000 12.535000 0.595000 ;
      RECT 12.365000  3.475000 12.535000 3.645000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.985000 12.805000 4.155000 ;
      RECT 12.725000  0.425000 12.895000 0.595000 ;
      RECT 12.725000  3.475000 12.895000 3.645000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.985000 13.285000 4.155000 ;
  END
END sky130_fd_sc_hvl__inv_16
MACRO sky130_fd_sc_hvl__inv_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__inv_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.200000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  9.000000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.310000 1.580000 6.760000 1.815000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  2.520000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.195000 0.730000 1.405000 1.230000 ;
        RECT 1.195000 1.230000 7.110000 1.395000 ;
        RECT 1.195000 1.395000 6.225000 1.400000 ;
        RECT 1.275000 2.035000 7.110000 2.205000 ;
        RECT 1.275000 2.205000 1.605000 3.445000 ;
        RECT 2.755000 0.730000 2.965000 1.230000 ;
        RECT 2.835000 2.205000 3.165000 3.445000 ;
        RECT 4.315000 0.730000 4.525000 1.230000 ;
        RECT 4.395000 2.205000 4.725000 3.445000 ;
        RECT 5.915000 0.730000 6.565000 1.225000 ;
        RECT 5.915000 1.225000 7.110000 1.230000 ;
        RECT 5.955000 2.205000 6.285000 3.445000 ;
        RECT 6.940000 1.395000 7.110000 2.035000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 7.200000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 7.200000 0.085000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 7.200000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 7.200000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.985000 7.200000 4.155000 ;
      LAYER mcon ;
        RECT 0.155000 3.985000 0.325000 4.155000 ;
        RECT 0.635000 3.985000 0.805000 4.155000 ;
        RECT 1.115000 3.985000 1.285000 4.155000 ;
        RECT 1.595000 3.985000 1.765000 4.155000 ;
        RECT 2.075000 3.985000 2.245000 4.155000 ;
        RECT 2.555000 3.985000 2.725000 4.155000 ;
        RECT 3.035000 3.985000 3.205000 4.155000 ;
        RECT 3.515000 3.985000 3.685000 4.155000 ;
        RECT 3.995000 3.985000 4.165000 4.155000 ;
        RECT 4.475000 3.985000 4.645000 4.155000 ;
        RECT 4.955000 3.985000 5.125000 4.155000 ;
        RECT 5.435000 3.985000 5.605000 4.155000 ;
        RECT 5.915000 3.985000 6.085000 4.155000 ;
        RECT 6.395000 3.985000 6.565000 4.155000 ;
        RECT 6.875000 3.985000 7.045000 4.155000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 7.200000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 7.530000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 7.200000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095000 0.380000 7.105000 0.550000 ;
      RECT 0.095000 0.550000 0.985000 1.385000 ;
      RECT 0.095000 2.445000 0.985000 3.625000 ;
      RECT 0.095000 3.625000 7.025000 3.795000 ;
      RECT 1.575000 0.550000 2.585000 1.045000 ;
      RECT 1.775000 2.385000 2.665000 3.625000 ;
      RECT 3.135000 0.550000 4.145000 1.045000 ;
      RECT 3.335000 2.385000 4.225000 3.625000 ;
      RECT 4.695000 0.550000 5.745000 1.045000 ;
      RECT 4.895000 2.385000 5.785000 3.625000 ;
      RECT 6.455000 2.385000 7.025000 3.625000 ;
      RECT 6.735000 0.550000 7.105000 1.045000 ;
    LAYER mcon ;
      RECT 0.095000 3.475000 0.265000 3.645000 ;
      RECT 0.455000 0.380000 0.625000 0.550000 ;
      RECT 0.455000 3.475000 0.625000 3.645000 ;
      RECT 0.815000 0.380000 0.985000 0.550000 ;
      RECT 0.815000 3.475000 0.985000 3.645000 ;
      RECT 1.175000 0.380000 1.345000 0.550000 ;
      RECT 1.535000 0.380000 1.705000 0.550000 ;
      RECT 1.775000 3.475000 1.945000 3.645000 ;
      RECT 1.895000 0.380000 2.065000 0.550000 ;
      RECT 2.135000 3.475000 2.305000 3.645000 ;
      RECT 2.255000 0.380000 2.425000 0.550000 ;
      RECT 2.495000 3.475000 2.665000 3.645000 ;
      RECT 2.615000 0.380000 2.785000 0.550000 ;
      RECT 2.975000 0.380000 3.145000 0.550000 ;
      RECT 3.335000 0.380000 3.505000 0.550000 ;
      RECT 3.335000 3.475000 3.505000 3.645000 ;
      RECT 3.695000 0.380000 3.865000 0.550000 ;
      RECT 3.695000 3.475000 3.865000 3.645000 ;
      RECT 4.055000 0.380000 4.225000 0.550000 ;
      RECT 4.055000 3.475000 4.225000 3.645000 ;
      RECT 4.415000 0.380000 4.585000 0.550000 ;
      RECT 4.775000 0.380000 4.945000 0.550000 ;
      RECT 4.895000 3.475000 5.065000 3.645000 ;
      RECT 5.135000 0.380000 5.305000 0.550000 ;
      RECT 5.255000 3.475000 5.425000 3.645000 ;
      RECT 5.495000 0.380000 5.665000 0.550000 ;
      RECT 5.615000 3.475000 5.785000 3.645000 ;
      RECT 5.855000 0.380000 6.025000 0.550000 ;
      RECT 6.215000 0.380000 6.385000 0.550000 ;
      RECT 6.455000 3.475000 6.625000 3.645000 ;
      RECT 6.575000 0.380000 6.745000 0.550000 ;
      RECT 6.855000 3.475000 7.025000 3.645000 ;
      RECT 6.935000 0.380000 7.105000 0.550000 ;
  END
END sky130_fd_sc_hvl__inv_8
MACRO sky130_fd_sc_hvl__fill_4
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hvl__fill_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.920000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 1.920000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 1.920000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 1.920000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 1.920000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 2.250000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 1.920000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.920000 0.085000 ;
      RECT 0.000000  3.985000 1.920000 4.155000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
  END
END sky130_fd_sc_hvl__fill_4
MACRO sky130_fd_sc_hvl__fill_2
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hvl__fill_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.960000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 0.960000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 0.960000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 0.960000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 0.960000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 1.290000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 0.960000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.960000 0.085000 ;
      RECT 0.000000  3.985000 0.960000 4.155000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
  END
END sky130_fd_sc_hvl__fill_2
MACRO sky130_fd_sc_hvl__fill_1
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hvl__fill_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.480000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 0.480000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 0.480000 0.085000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 0.480000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 0.480000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.985000 0.480000 4.155000 ;
      LAYER mcon ;
        RECT 0.155000 3.985000 0.325000 4.155000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 0.480000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 0.810000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 0.480000 3.815000 ;
    END
  END VPWR
END sky130_fd_sc_hvl__fill_1
MACRO sky130_fd_sc_hvl__fill_8
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hvl__fill_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 3.840000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 3.840000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 3.840000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 3.840000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 4.170000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 3.840000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.985000 3.840000 4.155000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.985000 3.685000 4.155000 ;
  END
END sky130_fd_sc_hvl__fill_8
MACRO sky130_fd_sc_hvl__schmittbuf_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__schmittbuf_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  1.170000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.015000 1.855000 3.305000 2.150000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.596250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.860000 0.515000 5.195000 3.715000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 5.280000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.280000 0.085000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 5.280000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 5.280000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.985000 5.280000 4.155000 ;
      LAYER mcon ;
        RECT 0.155000 3.985000 0.325000 4.155000 ;
        RECT 0.635000 3.985000 0.805000 4.155000 ;
        RECT 1.115000 3.985000 1.285000 4.155000 ;
        RECT 1.595000 3.985000 1.765000 4.155000 ;
        RECT 2.075000 3.985000 2.245000 4.155000 ;
        RECT 2.555000 3.985000 2.725000 4.155000 ;
        RECT 3.035000 3.985000 3.205000 4.155000 ;
        RECT 3.515000 3.985000 3.685000 4.155000 ;
        RECT 3.995000 3.985000 4.165000 4.155000 ;
        RECT 4.475000 3.985000 4.645000 4.155000 ;
        RECT 4.955000 3.985000 5.125000 4.155000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 5.280000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 1.340000 1.975000 ;
        RECT -0.330000 1.975000 5.610000 4.485000 ;
        RECT  3.885000 1.885000 5.610000 1.975000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 5.280000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 1.805000 0.530000 1.975000 ;
      RECT 0.085000 1.975000 0.255000 3.485000 ;
      RECT 0.085000 3.485000 1.030000 3.655000 ;
      RECT 0.280000 1.090000 0.530000 1.805000 ;
      RECT 0.430000 2.165000 0.875000 2.335000 ;
      RECT 0.430000 2.335000 0.680000 3.085000 ;
      RECT 0.705000 0.570000 2.010000 0.795000 ;
      RECT 0.705000 0.795000 0.875000 2.165000 ;
      RECT 0.740000 3.405000 1.030000 3.485000 ;
      RECT 0.740000 3.655000 1.030000 3.735000 ;
      RECT 1.045000 1.655000 4.690000 1.685000 ;
      RECT 1.045000 1.685000 1.835000 1.985000 ;
      RECT 1.060000 0.975000 2.720000 1.145000 ;
      RECT 1.060000 1.145000 1.390000 1.410000 ;
      RECT 1.200000 2.295000 1.460000 3.235000 ;
      RECT 1.200000 3.235000 2.790000 3.405000 ;
      RECT 1.600000 1.315000 1.940000 1.505000 ;
      RECT 1.600000 1.505000 4.210000 1.645000 ;
      RECT 1.600000 1.645000 4.690000 1.655000 ;
      RECT 1.655000 1.985000 1.835000 2.330000 ;
      RECT 1.655000 2.330000 2.010000 3.065000 ;
      RECT 2.390000 1.145000 2.720000 1.335000 ;
      RECT 2.460000 2.320000 2.790000 3.235000 ;
      RECT 3.120000 0.375000 4.630000 1.285000 ;
      RECT 3.130000 3.405000 4.570000 3.735000 ;
      RECT 3.235000 2.320000 4.570000 3.405000 ;
      RECT 3.855000 1.685000 4.690000 2.055000 ;
    LAYER mcon ;
      RECT 3.210000 0.425000 3.380000 0.595000 ;
      RECT 3.225000 3.475000 3.395000 3.645000 ;
      RECT 3.570000 0.425000 3.740000 0.595000 ;
      RECT 3.585000 3.475000 3.755000 3.645000 ;
      RECT 3.945000 3.475000 4.115000 3.645000 ;
      RECT 3.980000 0.425000 4.150000 0.595000 ;
      RECT 4.305000 3.475000 4.475000 3.645000 ;
      RECT 4.410000 0.425000 4.580000 0.595000 ;
  END
END sky130_fd_sc_hvl__schmittbuf_1
MACRO sky130_fd_sc_hvl__lsbufhv2lv_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__lsbufhv2lv_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  8.140000 ;
  SYMMETRY X Y ;
  SITE unithvdbl ;
  PIN A
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.630000 4.870000 1.300000 5.200000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.492900 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 0.735000 3.960000 3.245000 ;
    END
  END X
  PIN LVPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.070000 3.020000 8.090000 3.305000 ;
      LAYER nwell ;
        RECT 3.530000 1.925000 5.000000 5.575000 ;
    END
  END LVPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 7.515000 8.160000 7.885000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 8.025000 8.160000 8.255000 ;
      LAYER pwell ;
        RECT 0.000000 8.055000 8.160000 8.225000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 8.160000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 1.530000 6.255000 ;
        RECT  7.000000 1.885000 8.490000 6.255000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 4.325000 8.160000 4.695000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.985000 0.885000 4.155000 ;
      RECT 0.000000  8.055000 8.160000 8.225000 ;
      RECT 0.130000  2.260000 0.460000 3.445000 ;
      RECT 0.130000  3.445000 0.720000 3.675000 ;
      RECT 0.130000  4.465000 0.720000 4.695000 ;
      RECT 0.130000  4.695000 0.460000 5.880000 ;
      RECT 0.170000  1.080000 0.420000 1.565000 ;
      RECT 0.170000  1.565000 1.750000 1.895000 ;
      RECT 0.170000  6.220000 1.750000 6.575000 ;
      RECT 0.170000  6.575000 0.420000 7.060000 ;
      RECT 0.630000  2.835000 1.750000 3.085000 ;
      RECT 0.895000  0.395000 1.485000 1.395000 ;
      RECT 0.895000  6.745000 1.485000 7.745000 ;
      RECT 0.950000  1.895000 1.200000 2.590000 ;
      RECT 0.950000  5.550000 1.750000 6.220000 ;
      RECT 1.445000  1.895000 1.750000 2.235000 ;
      RECT 1.470000  3.085000 1.750000 5.550000 ;
      RECT 1.920000  0.685000 2.250000 4.255000 ;
      RECT 1.920000  4.255000 3.960000 4.595000 ;
      RECT 1.920000  5.195000 3.540000 5.445000 ;
      RECT 1.920000  5.445000 2.250000 7.455000 ;
      RECT 2.530000  5.615000 3.120000 7.745000 ;
      RECT 2.570000  0.395000 3.160000 3.910000 ;
      RECT 3.290000  5.445000 3.540000 5.595000 ;
      RECT 3.290000  5.595000 5.170000 5.845000 ;
      RECT 3.480000  5.845000 3.810000 7.455000 ;
      RECT 3.710000  4.595000 3.960000 5.415000 ;
      RECT 3.780000  3.415000 4.750000 4.085000 ;
      RECT 4.130000  0.395000 4.720000 1.515000 ;
      RECT 4.130000  2.085000 4.400000 3.075000 ;
      RECT 4.130000  3.075000 4.750000 3.415000 ;
      RECT 4.130000  4.085000 4.400000 5.415000 ;
      RECT 4.570000  2.085000 4.820000 2.655000 ;
      RECT 4.570000  2.655000 5.170000 2.905000 ;
      RECT 4.920000  2.905000 5.170000 5.595000 ;
      RECT 7.275000  3.985000 8.160000 4.155000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.155000  8.055000 0.325000 8.225000 ;
      RECT 0.160000  3.475000 0.330000 3.645000 ;
      RECT 0.160000  4.495000 0.330000 4.665000 ;
      RECT 0.520000  3.475000 0.690000 3.645000 ;
      RECT 0.520000  4.495000 0.690000 4.665000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.635000  8.055000 0.805000 8.225000 ;
      RECT 0.925000  0.425000 1.095000 0.595000 ;
      RECT 0.925000  7.545000 1.095000 7.715000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  8.055000 1.285000 8.225000 ;
      RECT 1.285000  0.425000 1.455000 0.595000 ;
      RECT 1.285000  7.545000 1.455000 7.715000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  8.055000 1.765000 8.225000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  8.055000 2.245000 8.225000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  8.055000 2.725000 8.225000 ;
      RECT 2.560000  7.545000 2.730000 7.715000 ;
      RECT 2.600000  0.425000 2.770000 0.595000 ;
      RECT 2.920000  7.545000 3.090000 7.715000 ;
      RECT 2.960000  0.425000 3.130000 0.595000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  8.055000 3.205000 8.225000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  8.055000 3.685000 8.225000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  8.055000 4.165000 8.225000 ;
      RECT 4.160000  0.425000 4.330000 0.595000 ;
      RECT 4.160000  3.105000 4.330000 3.275000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  8.055000 4.645000 8.225000 ;
      RECT 4.520000  0.425000 4.690000 0.595000 ;
      RECT 4.520000  3.105000 4.690000 3.275000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  8.055000 5.125000 8.225000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  8.055000 5.605000 8.225000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  8.055000 6.085000 8.225000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  8.055000 6.565000 8.225000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  8.055000 7.045000 8.225000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.985000 7.525000 4.155000 ;
      RECT 7.355000  8.055000 7.525000 8.225000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.985000 8.005000 4.155000 ;
      RECT 7.835000  8.055000 8.005000 8.225000 ;
    LAYER met1 ;
      RECT 0.000000 -0.115000 8.160000 0.115000 ;
      RECT 0.000000  0.255000 8.160000 0.625000 ;
      RECT 0.000000  3.445000 8.160000 3.815000 ;
    LAYER pwell ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
  END
END sky130_fd_sc_hvl__lsbufhv2lv_1
MACRO sky130_fd_sc_hvl__sdfxbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__sdfxbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  19.68000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN D
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.165000 1.175000 4.675000 2.150000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.611250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.955000 0.495000 16.285000 2.025000 ;
        RECT 15.955000 2.025000 16.545000 2.515000 ;
        RECT 16.215000 2.515000 16.545000 3.455000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.641250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 19.220000 0.495000 19.555000 3.755000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.930000 1.975000 2.440000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.840000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.565000 1.550000 2.755000 1.750000 ;
        RECT 0.565000 1.750000 0.895000 2.220000 ;
        RECT 2.425000 1.750000 2.755000 2.745000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 10.685000 1.895000 11.395000 2.120000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 19.680000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 19.680000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 19.680000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 19.680000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 20.010000 4.485000 ;
        RECT 15.925000 1.715000 18.490000 1.885000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 19.680000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 19.680000 0.085000 ;
      RECT  0.000000  3.985000 19.680000 4.155000 ;
      RECT  0.110000  1.175000  3.330000 1.345000 ;
      RECT  0.110000  1.345000  0.280000 2.555000 ;
      RECT  0.110000  2.555000  0.440000 3.015000 ;
      RECT  0.540000  0.495000  0.870000 1.175000 ;
      RECT  0.630000  2.620000  1.220000 3.705000 ;
      RECT  1.050000  0.365000  2.000000 0.995000 ;
      RECT  1.400000  2.925000  3.680000 3.095000 ;
      RECT  1.400000  3.095000  1.570000 3.755000 ;
      RECT  1.750000  3.335000  2.700000 3.755000 ;
      RECT  2.810000  0.495000  3.140000 0.825000 ;
      RECT  2.810000  0.825000  3.680000 0.995000 ;
      RECT  2.880000  3.275000  3.210000 3.610000 ;
      RECT  2.880000  3.610000  4.030000 3.780000 ;
      RECT  3.065000  1.345000  3.330000 1.845000 ;
      RECT  3.430000  3.095000  3.680000 3.430000 ;
      RECT  3.510000  0.995000  3.680000 2.330000 ;
      RECT  3.510000  2.330000  5.135000 2.500000 ;
      RECT  3.860000  0.365000  4.785000 0.995000 ;
      RECT  3.860000  2.680000  5.240000 2.850000 ;
      RECT  3.860000  2.850000  4.030000 3.610000 ;
      RECT  4.210000  3.030000  4.540000 3.635000 ;
      RECT  4.210000  3.635000  6.140000 3.805000 ;
      RECT  4.965000  0.265000  5.995000 0.435000 ;
      RECT  4.965000  0.435000  5.135000 2.330000 ;
      RECT  4.990000  2.850000  5.240000 3.430000 ;
      RECT  5.315000  0.615000  5.645000 1.605000 ;
      RECT  5.315000  1.605000  7.120000 1.775000 ;
      RECT  5.420000  1.775000  5.790000 3.455000 ;
      RECT  5.825000  0.435000  5.995000 1.255000 ;
      RECT  5.825000  1.255000  8.165000 1.425000 ;
      RECT  5.970000  1.955000  7.470000 2.125000 ;
      RECT  5.970000  2.125000  6.140000 3.115000 ;
      RECT  5.970000  3.115000  7.560000 3.285000 ;
      RECT  5.970000  3.285000  6.140000 3.635000 ;
      RECT  6.175000  0.365000  7.065000 1.075000 ;
      RECT  6.320000  2.305000  7.910000 2.555000 ;
      RECT  6.320000  3.465000  7.210000 3.755000 ;
      RECT  7.245000  0.590000  9.725000 0.760000 ;
      RECT  7.245000  0.760000  7.575000 1.075000 ;
      RECT  7.300000  1.425000  7.470000 1.955000 ;
      RECT  7.390000  3.285000  9.435000 3.455000 ;
      RECT  7.740000  2.135000  8.785000 2.305000 ;
      RECT  7.740000  2.555000  7.910000 2.855000 ;
      RECT  7.740000  2.855000  8.655000 3.105000 ;
      RECT  7.835000  0.940000  8.165000 1.255000 ;
      RECT  8.090000  2.485000  9.005000 2.675000 ;
      RECT  8.615000  0.940000  8.945000 1.360000 ;
      RECT  8.615000  1.360000  8.785000 2.135000 ;
      RECT  8.835000  2.675000  9.005000 2.750000 ;
      RECT  8.835000  2.750000 10.355000 2.920000 ;
      RECT  9.070000  1.545000 12.130000 1.715000 ;
      RECT  9.070000  1.715000  9.400000 2.215000 ;
      RECT  9.105000  3.100000  9.435000 3.285000 ;
      RECT  9.395000  0.760000  9.725000 1.360000 ;
      RECT  9.675000  1.715000  9.845000 2.320000 ;
      RECT  9.675000  2.320000 10.005000 2.570000 ;
      RECT  9.985000  0.495000 10.315000 1.545000 ;
      RECT 10.025000  1.895000 10.355000 2.140000 ;
      RECT 10.185000  2.140000 10.355000 2.300000 ;
      RECT 10.185000  2.300000 11.565000 2.470000 ;
      RECT 10.185000  2.470000 10.355000 2.750000 ;
      RECT 10.495000  0.365000 11.445000 0.915000 ;
      RECT 10.495000  1.095000 11.875000 1.265000 ;
      RECT 10.495000  1.265000 10.825000 1.365000 ;
      RECT 10.535000  2.650000 11.125000 3.705000 ;
      RECT 11.315000  2.470000 11.565000 3.110000 ;
      RECT 11.625000  0.475000 13.610000 0.645000 ;
      RECT 11.625000  0.645000 11.875000 1.095000 ;
      RECT 11.785000  2.205000 12.115000 3.635000 ;
      RECT 11.785000  3.635000 14.340000 3.805000 ;
      RECT 11.800000  1.445000 12.130000 1.545000 ;
      RECT 11.800000  1.715000 12.130000 2.025000 ;
      RECT 12.150000  0.825000 12.480000 1.245000 ;
      RECT 12.310000  1.245000 12.480000 3.285000 ;
      RECT 12.310000  3.285000 13.795000 3.455000 ;
      RECT 12.660000  2.205000 12.990000 3.105000 ;
      RECT 12.820000  0.825000 13.260000 1.325000 ;
      RECT 12.820000  1.325000 12.990000 1.915000 ;
      RECT 12.820000  1.915000 15.135000 2.085000 ;
      RECT 12.820000  2.085000 12.990000 2.205000 ;
      RECT 13.280000  1.505000 13.610000 1.735000 ;
      RECT 13.440000  0.645000 13.610000 1.505000 ;
      RECT 13.440000  2.265000 13.795000 3.285000 ;
      RECT 13.915000  0.365000 14.865000 1.325000 ;
      RECT 14.010000  2.695000 14.340000 3.635000 ;
      RECT 14.465000  2.265000 15.775000 2.515000 ;
      RECT 14.520000  2.695000 15.425000 3.735000 ;
      RECT 14.805000  1.545000 15.135000 1.915000 ;
      RECT 15.315000  0.495000 15.775000 2.265000 ;
      RECT 15.605000  2.515000 15.775000 2.695000 ;
      RECT 15.605000  2.695000 15.995000 3.635000 ;
      RECT 15.605000  3.635000 16.895000 3.805000 ;
      RECT 16.465000  0.365000 17.415000 1.325000 ;
      RECT 16.725000  1.505000 17.055000 1.835000 ;
      RECT 16.725000  1.835000 16.895000 3.635000 ;
      RECT 17.075000  2.025000 17.665000 3.705000 ;
      RECT 17.630000  0.495000 17.960000 1.505000 ;
      RECT 17.630000  1.505000 19.040000 1.675000 ;
      RECT 17.870000  2.025000 18.200000 2.815000 ;
      RECT 18.030000  1.675000 19.040000 1.835000 ;
      RECT 18.030000  1.835000 18.200000 2.025000 ;
      RECT 18.140000  0.365000 19.040000 1.325000 ;
      RECT 18.380000  2.175000 18.970000 3.755000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.985000  0.325000 4.155000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.985000  0.805000 4.155000 ;
      RECT  0.660000  3.505000  0.830000 3.675000 ;
      RECT  1.020000  3.505000  1.190000 3.675000 ;
      RECT  1.080000  0.395000  1.250000 0.565000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.985000  1.285000 4.155000 ;
      RECT  1.440000  0.395000  1.610000 0.565000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.985000  1.765000 4.155000 ;
      RECT  1.780000  3.505000  1.950000 3.675000 ;
      RECT  1.800000  0.395000  1.970000 0.565000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.985000  2.245000 4.155000 ;
      RECT  2.140000  3.505000  2.310000 3.675000 ;
      RECT  2.500000  3.505000  2.670000 3.675000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.985000  2.725000 4.155000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.985000  3.205000 4.155000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.985000  3.685000 4.155000 ;
      RECT  3.875000  0.395000  4.045000 0.565000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.985000  4.165000 4.155000 ;
      RECT  4.235000  0.395000  4.405000 0.565000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.985000  4.645000 4.155000 ;
      RECT  4.595000  0.395000  4.765000 0.565000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.985000  5.125000 4.155000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.060000  5.605000 3.230000 ;
      RECT  5.435000  3.985000  5.605000 4.155000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.985000  6.085000 4.155000 ;
      RECT  6.175000  0.395000  6.345000 0.565000 ;
      RECT  6.320000  3.505000  6.490000 3.675000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.985000  6.565000 4.155000 ;
      RECT  6.535000  0.395000  6.705000 0.565000 ;
      RECT  6.680000  3.505000  6.850000 3.675000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.985000  7.045000 4.155000 ;
      RECT  6.895000  0.395000  7.065000 0.565000 ;
      RECT  7.040000  3.505000  7.210000 3.675000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.985000  7.525000 4.155000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.985000  8.005000 4.155000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.985000  8.485000 4.155000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.985000  8.965000 4.155000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.985000  9.445000 4.155000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.985000  9.925000 4.155000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.985000 10.405000 4.155000 ;
      RECT 10.525000  0.395000 10.695000 0.565000 ;
      RECT 10.565000  3.505000 10.735000 3.675000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.985000 10.885000 4.155000 ;
      RECT 10.885000  0.395000 11.055000 0.565000 ;
      RECT 10.925000  3.505000 11.095000 3.675000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.985000 11.365000 4.155000 ;
      RECT 11.245000  0.395000 11.415000 0.565000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.985000 11.845000 4.155000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.985000 12.325000 4.155000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.985000 12.805000 4.155000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.985000 13.285000 4.155000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.060000 13.765000 3.230000 ;
      RECT 13.595000  3.985000 13.765000 4.155000 ;
      RECT 13.945000  0.395000 14.115000 0.565000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.985000 14.245000 4.155000 ;
      RECT 14.305000  0.395000 14.475000 0.565000 ;
      RECT 14.525000  3.505000 14.695000 3.675000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.985000 14.725000 4.155000 ;
      RECT 14.665000  0.395000 14.835000 0.565000 ;
      RECT 14.885000  3.505000 15.055000 3.675000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.985000 15.205000 4.155000 ;
      RECT 15.245000  3.505000 15.415000 3.675000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.985000 15.685000 4.155000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000  3.985000 16.165000 4.155000 ;
      RECT 16.475000 -0.085000 16.645000 0.085000 ;
      RECT 16.475000  3.985000 16.645000 4.155000 ;
      RECT 16.495000  0.395000 16.665000 0.565000 ;
      RECT 16.855000  0.395000 17.025000 0.565000 ;
      RECT 16.955000 -0.085000 17.125000 0.085000 ;
      RECT 16.955000  3.985000 17.125000 4.155000 ;
      RECT 17.105000  3.505000 17.275000 3.675000 ;
      RECT 17.215000  0.395000 17.385000 0.565000 ;
      RECT 17.435000 -0.085000 17.605000 0.085000 ;
      RECT 17.435000  3.985000 17.605000 4.155000 ;
      RECT 17.465000  3.505000 17.635000 3.675000 ;
      RECT 17.915000 -0.085000 18.085000 0.085000 ;
      RECT 17.915000  3.985000 18.085000 4.155000 ;
      RECT 18.145000  0.395000 18.315000 0.565000 ;
      RECT 18.395000 -0.085000 18.565000 0.085000 ;
      RECT 18.395000  3.985000 18.565000 4.155000 ;
      RECT 18.410000  3.505000 18.580000 3.675000 ;
      RECT 18.505000  0.395000 18.675000 0.565000 ;
      RECT 18.770000  3.505000 18.940000 3.675000 ;
      RECT 18.865000  0.395000 19.035000 0.565000 ;
      RECT 18.875000 -0.085000 19.045000 0.085000 ;
      RECT 18.875000  3.985000 19.045000 4.155000 ;
      RECT 19.355000 -0.085000 19.525000 0.085000 ;
      RECT 19.355000  3.985000 19.525000 4.155000 ;
    LAYER met1 ;
      RECT  5.375000 3.030000  5.665000 3.075000 ;
      RECT  5.375000 3.075000 13.825000 3.215000 ;
      RECT  5.375000 3.215000  5.665000 3.260000 ;
      RECT 13.535000 3.030000 13.825000 3.075000 ;
      RECT 13.535000 3.215000 13.825000 3.260000 ;
  END
END sky130_fd_sc_hvl__sdfxbp_1
MACRO sky130_fd_sc_hvl__dfrbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__dfrbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  16.80000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN D
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.850000 0.810000 4.165000 2.105000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.626250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 16.340000 0.515000 16.690000 3.755000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.641250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.045000 0.665000 14.425000 1.495000 ;
        RECT 14.045000 1.495000 14.380000 1.780000 ;
        RECT 14.130000 1.780000 14.380000 3.755000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  2.980000 1.505000  3.665000 2.120000 ;
        RECT  3.495000 0.460000  6.625000 0.630000 ;
        RECT  3.495000 0.630000  3.665000 1.505000 ;
        RECT  6.455000 0.630000  6.625000 1.125000 ;
        RECT  6.455000 1.125000  8.515000 1.295000 ;
        RECT  7.165000 1.825000  8.515000 1.995000 ;
        RECT  8.345000 0.265000 11.075000 0.435000 ;
        RECT  8.345000 0.435000  8.515000 1.125000 ;
        RECT  8.345000 1.295000  8.515000 1.825000 ;
        RECT 10.905000 0.435000 11.075000 0.960000 ;
        RECT 10.905000 0.960000 11.840000 1.130000 ;
        RECT 11.510000 1.130000 11.840000 1.350000 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.595000 1.175000 0.925000 1.720000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 16.800000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 16.800000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 16.800000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 16.800000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 17.130000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 16.800000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 16.800000 0.085000 ;
      RECT  0.000000  3.985000 16.800000 4.155000 ;
      RECT  0.165000  0.495000  0.495000 0.995000 ;
      RECT  0.165000  0.995000  0.415000 2.275000 ;
      RECT  0.165000  2.275000  1.835000 2.445000 ;
      RECT  0.165000  2.445000  0.415000 3.455000 ;
      RECT  0.595000  2.625000  1.485000 3.705000 ;
      RECT  0.675000  0.365000  1.625000 0.995000 ;
      RECT  1.505000  1.900000  1.835000 2.275000 ;
      RECT  1.665000  2.445000  1.835000 3.635000 ;
      RECT  1.665000  3.635000  3.205000 3.805000 ;
      RECT  1.805000  0.495000  2.185000 0.995000 ;
      RECT  2.015000  0.995000  2.185000 1.550000 ;
      RECT  2.015000  1.550000  2.275000 3.455000 ;
      RECT  2.365000  0.365000  3.315000 1.325000 ;
      RECT  2.525000  2.300000  4.515000 2.470000 ;
      RECT  2.525000  2.470000  2.855000 3.420000 ;
      RECT  3.035000  2.650000  3.905000 2.820000 ;
      RECT  3.035000  2.820000  3.205000 3.635000 ;
      RECT  3.385000  3.000000  3.555000 3.705000 ;
      RECT  3.735000  2.820000  3.905000 3.600000 ;
      RECT  3.735000  3.600000  5.565000 3.770000 ;
      RECT  4.085000  3.000000  4.515000 3.420000 ;
      RECT  4.345000  0.825000  4.655000 1.325000 ;
      RECT  4.345000  1.325000  4.515000 2.300000 ;
      RECT  4.345000  2.470000  4.515000 3.000000 ;
      RECT  4.695000  1.505000  5.925000 1.780000 ;
      RECT  4.695000  1.780000  4.865000 2.820000 ;
      RECT  4.865000  3.000000  5.215000 3.420000 ;
      RECT  5.045000  2.200000  6.275000 2.370000 ;
      RECT  5.045000  2.370000  5.215000 3.000000 ;
      RECT  5.270000  0.825000  5.600000 1.155000 ;
      RECT  5.270000  1.155000  6.275000 1.325000 ;
      RECT  5.395000  2.550000  5.650000 2.875000 ;
      RECT  5.395000  2.875000  7.035000 3.045000 ;
      RECT  5.395000  3.045000  5.565000 3.600000 ;
      RECT  5.595000  1.780000  5.925000 2.020000 ;
      RECT  5.745000  3.225000  6.685000 3.705000 ;
      RECT  6.105000  1.325000  6.275000 1.475000 ;
      RECT  6.105000  1.475000  8.165000 1.645000 ;
      RECT  6.105000  1.645000  6.275000 2.200000 ;
      RECT  6.105000  2.370000  6.275000 2.525000 ;
      RECT  6.105000  2.525000  7.385000 2.695000 ;
      RECT  6.455000  1.825000  6.785000 2.175000 ;
      RECT  6.455000  2.175000  9.025000 2.345000 ;
      RECT  6.865000  3.045000  7.035000 3.635000 ;
      RECT  6.865000  3.635000  7.735000 3.805000 ;
      RECT  7.215000  0.365000  8.165000 0.945000 ;
      RECT  7.215000  2.695000  7.385000 3.455000 ;
      RECT  7.565000  2.700000  9.375000 2.870000 ;
      RECT  7.565000  2.870000  7.735000 3.635000 ;
      RECT  7.915000  3.050000  8.865000 3.705000 ;
      RECT  8.695000  0.615000  9.025000 2.175000 ;
      RECT  8.695000  2.345000  9.025000 2.520000 ;
      RECT  9.205000  1.230000 10.375000 1.400000 ;
      RECT  9.205000  1.400000  9.375000 2.700000 ;
      RECT  9.555000  2.270000 10.410000 2.440000 ;
      RECT  9.555000  2.440000  9.805000 3.350000 ;
      RECT  9.580000  0.615000 10.725000 0.785000 ;
      RECT  9.580000  0.785000  9.910000 0.995000 ;
      RECT  9.725000  1.580000 10.060000 2.090000 ;
      RECT 10.090000  1.070000 10.375000 1.230000 ;
      RECT 10.240000  2.000000 12.530000 2.170000 ;
      RECT 10.240000  2.170000 10.410000 2.270000 ;
      RECT 10.555000  0.785000 10.725000 2.000000 ;
      RECT 10.590000  2.350000 11.540000 3.705000 ;
      RECT 10.930000  1.310000 11.260000 1.530000 ;
      RECT 10.930000  1.530000 12.880000 1.700000 ;
      RECT 10.930000  1.700000 11.260000 1.820000 ;
      RECT 11.255000  0.365000 12.205000 0.780000 ;
      RECT 11.965000  2.350000 12.880000 2.520000 ;
      RECT 11.965000  2.520000 12.295000 2.770000 ;
      RECT 12.200000  1.880000 12.530000 2.000000 ;
      RECT 12.710000  0.515000 13.075000 0.975000 ;
      RECT 12.710000  0.975000 12.880000 1.530000 ;
      RECT 12.710000  1.700000 12.880000 2.350000 ;
      RECT 13.060000  2.175000 13.950000 3.755000 ;
      RECT 13.255000  0.365000 13.845000 1.495000 ;
      RECT 14.665000  0.825000 15.015000 1.505000 ;
      RECT 14.665000  1.505000 16.160000 1.835000 ;
      RECT 14.665000  1.835000 14.995000 3.005000 ;
      RECT 15.175000  2.175000 16.125000 3.755000 ;
      RECT 15.195000  0.365000 16.145000 1.325000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.985000  0.325000 4.155000 ;
      RECT  0.595000  3.505000  0.765000 3.675000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.985000  0.805000 4.155000 ;
      RECT  0.705000  0.395000  0.875000 0.565000 ;
      RECT  0.955000  3.505000  1.125000 3.675000 ;
      RECT  1.065000  0.395000  1.235000 0.565000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.985000  1.285000 4.155000 ;
      RECT  1.315000  3.505000  1.485000 3.675000 ;
      RECT  1.425000  0.395000  1.595000 0.565000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.985000  1.765000 4.155000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  1.580000  2.245000 1.750000 ;
      RECT  2.075000  3.985000  2.245000 4.155000 ;
      RECT  2.395000  0.395000  2.565000 0.565000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.985000  2.725000 4.155000 ;
      RECT  2.755000  0.395000  2.925000 0.565000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.985000  3.205000 4.155000 ;
      RECT  3.115000  0.395000  3.285000 0.565000 ;
      RECT  3.385000  3.505000  3.555000 3.675000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.985000  3.685000 4.155000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.985000  4.165000 4.155000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.985000  4.645000 4.155000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  1.580000  5.125000 1.750000 ;
      RECT  4.955000  3.985000  5.125000 4.155000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.985000  5.605000 4.155000 ;
      RECT  5.770000  3.505000  5.940000 3.675000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.985000  6.085000 4.155000 ;
      RECT  6.130000  3.505000  6.300000 3.675000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.985000  6.565000 4.155000 ;
      RECT  6.490000  3.505000  6.660000 3.675000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.985000  7.045000 4.155000 ;
      RECT  7.245000  0.395000  7.415000 0.565000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.985000  7.525000 4.155000 ;
      RECT  7.605000  0.395000  7.775000 0.565000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.985000  8.005000 4.155000 ;
      RECT  7.945000  3.505000  8.115000 3.675000 ;
      RECT  7.965000  0.395000  8.135000 0.565000 ;
      RECT  8.305000  3.505000  8.475000 3.675000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.985000  8.485000 4.155000 ;
      RECT  8.665000  3.505000  8.835000 3.675000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.985000  8.965000 4.155000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.985000  9.445000 4.155000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  1.580000  9.925000 1.750000 ;
      RECT  9.755000  3.985000  9.925000 4.155000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.985000 10.405000 4.155000 ;
      RECT 10.620000  3.505000 10.790000 3.675000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.985000 10.885000 4.155000 ;
      RECT 10.980000  3.505000 11.150000 3.675000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.985000 11.365000 4.155000 ;
      RECT 11.285000  0.395000 11.455000 0.565000 ;
      RECT 11.340000  3.505000 11.510000 3.675000 ;
      RECT 11.645000  0.395000 11.815000 0.565000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.985000 11.845000 4.155000 ;
      RECT 12.005000  0.395000 12.175000 0.565000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.985000 12.325000 4.155000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.985000 12.805000 4.155000 ;
      RECT 13.060000  3.505000 13.230000 3.675000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.985000 13.285000 4.155000 ;
      RECT 13.285000  0.395000 13.455000 0.565000 ;
      RECT 13.420000  3.505000 13.590000 3.675000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.985000 13.765000 4.155000 ;
      RECT 13.645000  0.395000 13.815000 0.565000 ;
      RECT 13.780000  3.505000 13.950000 3.675000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.985000 14.245000 4.155000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.985000 14.725000 4.155000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.985000 15.205000 4.155000 ;
      RECT 15.205000  3.505000 15.375000 3.675000 ;
      RECT 15.225000  0.395000 15.395000 0.565000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.985000 15.685000 4.155000 ;
      RECT 15.565000  3.505000 15.735000 3.675000 ;
      RECT 15.585000  0.395000 15.755000 0.565000 ;
      RECT 15.925000  3.505000 16.095000 3.675000 ;
      RECT 15.945000  0.395000 16.115000 0.565000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000  3.985000 16.165000 4.155000 ;
      RECT 16.475000 -0.085000 16.645000 0.085000 ;
      RECT 16.475000  3.985000 16.645000 4.155000 ;
    LAYER met1 ;
      RECT 2.015000 1.550000 2.305000 1.595000 ;
      RECT 2.015000 1.595000 9.985000 1.735000 ;
      RECT 2.015000 1.735000 2.305000 1.780000 ;
      RECT 4.895000 1.550000 5.185000 1.595000 ;
      RECT 4.895000 1.735000 5.185000 1.780000 ;
      RECT 9.695000 1.550000 9.985000 1.595000 ;
      RECT 9.695000 1.735000 9.985000 1.780000 ;
  END
END sky130_fd_sc_hvl__dfrbp_1
MACRO sky130_fd_sc_hvl__dlxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__dlxtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN D
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.795000 3.100000 2.465000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.626250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.700000 0.515000 8.050000 3.755000 ;
    END
  END Q
  PIN GATE
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.540000 1.175000 0.870000 1.725000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 8.160000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 8.160000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 8.160000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 8.160000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 8.490000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 8.160000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.985000 8.160000 4.155000 ;
      RECT 0.110000  0.495000 0.665000 0.995000 ;
      RECT 0.110000  0.995000 0.360000 1.905000 ;
      RECT 0.110000  1.905000 1.795000 2.015000 ;
      RECT 0.110000  2.015000 1.780000 2.075000 ;
      RECT 0.110000  2.075000 0.360000 2.985000 ;
      RECT 0.540000  2.255000 1.430000 3.705000 ;
      RECT 0.845000  0.365000 1.795000 0.995000 ;
      RECT 1.540000  1.345000 1.795000 1.905000 ;
      RECT 1.610000  2.075000 1.780000 2.645000 ;
      RECT 1.610000  2.645000 3.190000 2.815000 ;
      RECT 1.890000  2.995000 2.840000 3.705000 ;
      RECT 1.960000  2.195000 2.290000 2.465000 ;
      RECT 1.975000  0.515000 2.225000 1.445000 ;
      RECT 1.975000  1.445000 3.880000 1.615000 ;
      RECT 1.975000  1.615000 2.290000 2.195000 ;
      RECT 2.405000  0.365000 2.995000 0.975000 ;
      RECT 3.020000  2.815000 3.190000 3.635000 ;
      RECT 3.020000  3.635000 4.050000 3.805000 ;
      RECT 3.225000  0.495000 3.555000 0.995000 ;
      RECT 3.370000  2.165000 4.230000 2.335000 ;
      RECT 3.370000  2.335000 3.540000 2.895000 ;
      RECT 3.370000  2.895000 3.700000 3.455000 ;
      RECT 3.385000  0.995000 3.555000 1.095000 ;
      RECT 3.385000  1.095000 4.230000 1.265000 ;
      RECT 3.550000  1.615000 3.880000 1.985000 ;
      RECT 3.720000  2.515000 4.740000 2.715000 ;
      RECT 3.880000  2.715000 4.050000 3.635000 ;
      RECT 4.005000  0.495000 4.335000 0.745000 ;
      RECT 4.005000  0.745000 5.090000 0.915000 ;
      RECT 4.060000  1.265000 4.230000 2.165000 ;
      RECT 4.230000  2.895000 5.090000 3.065000 ;
      RECT 4.230000  3.065000 4.480000 3.725000 ;
      RECT 4.410000  1.095000 4.740000 2.515000 ;
      RECT 4.920000  0.915000 5.090000 1.835000 ;
      RECT 4.920000  1.835000 6.680000 2.005000 ;
      RECT 4.920000  2.005000 5.090000 2.895000 ;
      RECT 5.270000  0.365000 5.860000 0.895000 ;
      RECT 5.270000  2.895000 6.220000 3.705000 ;
      RECT 5.430000  1.075000 5.760000 1.425000 ;
      RECT 5.430000  1.425000 7.030000 1.595000 ;
      RECT 5.430000  1.595000 5.760000 1.655000 ;
      RECT 6.025000  2.185000 7.030000 2.355000 ;
      RECT 6.025000  2.355000 6.355000 2.675000 ;
      RECT 6.045000  0.845000 6.375000 1.425000 ;
      RECT 6.350000  1.775000 6.680000 1.835000 ;
      RECT 6.535000  2.535000 7.485000 3.755000 ;
      RECT 6.555000  0.365000 7.505000 1.245000 ;
      RECT 6.860000  1.595000 7.030000 2.185000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.540000  3.505000 0.710000 3.675000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.875000  0.395000 1.045000 0.565000 ;
      RECT 0.900000  3.505000 1.070000 3.675000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.235000  0.395000 1.405000 0.565000 ;
      RECT 1.260000  3.505000 1.430000 3.675000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  0.395000 1.765000 0.565000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.920000  3.505000 2.090000 3.675000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.280000  3.505000 2.450000 3.675000 ;
      RECT 2.435000  0.395000 2.605000 0.565000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 2.640000  3.505000 2.810000 3.675000 ;
      RECT 2.795000  0.395000 2.965000 0.565000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.985000 3.685000 4.155000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.985000 4.165000 4.155000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.985000 4.645000 4.155000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.985000 5.125000 4.155000 ;
      RECT 5.300000  0.395000 5.470000 0.565000 ;
      RECT 5.300000  3.505000 5.470000 3.675000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.985000 5.605000 4.155000 ;
      RECT 5.660000  0.395000 5.830000 0.565000 ;
      RECT 5.660000  3.505000 5.830000 3.675000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.985000 6.085000 4.155000 ;
      RECT 6.020000  3.505000 6.190000 3.675000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.985000 6.565000 4.155000 ;
      RECT 6.565000  3.505000 6.735000 3.675000 ;
      RECT 6.585000  0.395000 6.755000 0.565000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.985000 7.045000 4.155000 ;
      RECT 6.925000  3.505000 7.095000 3.675000 ;
      RECT 6.945000  0.395000 7.115000 0.565000 ;
      RECT 7.285000  3.505000 7.455000 3.675000 ;
      RECT 7.305000  0.395000 7.475000 0.565000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.985000 7.525000 4.155000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.985000 8.005000 4.155000 ;
  END
END sky130_fd_sc_hvl__dlxtp_1
MACRO sky130_fd_sc_hvl__or3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__or3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.915000 1.080000 2.450000 1.390000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.910000 1.535000 3.260000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.530000 1.080000 1.315000 1.390000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.626250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.460000 0.495000 3.715000 3.755000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 3.840000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 3.840000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 3.840000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 3.840000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 4.170000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 3.840000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.985000 3.840000 4.155000 ;
      RECT 0.145000  0.495000 0.360000 1.560000 ;
      RECT 0.145000  1.560000 3.255000 1.730000 ;
      RECT 0.145000  1.730000 0.395000 2.780000 ;
      RECT 0.530000  0.365000 1.385000 0.910000 ;
      RECT 1.565000  0.495000 1.965000 0.910000 ;
      RECT 1.565000  0.910000 1.735000 1.560000 ;
      RECT 1.620000  3.430000 3.280000 3.755000 ;
      RECT 1.705000  2.175000 3.280000 3.430000 ;
      RECT 2.620000  0.365000 3.290000 1.325000 ;
      RECT 2.925000  1.730000 3.255000 1.935000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.580000  0.395000 0.750000 0.565000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.165000  0.395000 1.335000 0.565000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.670000  3.505000 1.840000 3.675000 ;
      RECT 2.030000  3.505000 2.200000 3.675000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.390000  3.505000 2.560000 3.675000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 2.690000  0.395000 2.860000 0.565000 ;
      RECT 2.750000  3.505000 2.920000 3.675000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
      RECT 3.050000  0.395000 3.220000 0.565000 ;
      RECT 3.110000  3.505000 3.280000 3.675000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.985000 3.685000 4.155000 ;
  END
END sky130_fd_sc_hvl__or3_1
MACRO sky130_fd_sc_hvl__xor2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__xor2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  2.250000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.775000 3.235000 2.150000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  2.250000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.560000 1.775000 1.510000 2.055000 ;
        RECT 1.340000 1.425000 3.585000 1.505000 ;
        RECT 1.340000 1.505000 3.715000 1.595000 ;
        RECT 1.340000 1.595000 1.510000 1.775000 ;
        RECT 3.415000 1.595000 3.715000 1.835000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.637500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.850000 0.495000 4.370000 1.325000 ;
        RECT 3.965000 1.325000 4.370000 2.425000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 5.280000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 5.280000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 5.280000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 5.280000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 5.610000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 5.280000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.280000 0.085000 ;
      RECT 0.000000  3.985000 5.280000 4.155000 ;
      RECT 0.090000  0.365000 0.680000 1.245000 ;
      RECT 0.130000  1.425000 1.160000 1.595000 ;
      RECT 0.130000  1.595000 0.380000 2.435000 ;
      RECT 0.130000  2.435000 3.230000 2.605000 ;
      RECT 0.130000  2.605000 0.380000 3.755000 ;
      RECT 0.560000  2.785000 2.530000 3.755000 ;
      RECT 0.910000  0.495000 1.160000 1.425000 ;
      RECT 1.340000  0.365000 3.670000 1.245000 ;
      RECT 2.710000  2.785000 2.880000 2.955000 ;
      RECT 2.710000  2.955000 5.150000 3.125000 ;
      RECT 2.710000  3.125000 2.880000 3.755000 ;
      RECT 3.060000  2.605000 4.720000 2.775000 ;
      RECT 3.060000  3.305000 4.720000 3.755000 ;
      RECT 4.550000  0.365000 5.140000 1.325000 ;
      RECT 4.550000  1.665000 4.880000 1.995000 ;
      RECT 4.550000  1.995000 4.720000 2.605000 ;
      RECT 4.900000  2.175000 5.150000 2.955000 ;
      RECT 4.900000  3.125000 5.150000 3.755000 ;
    LAYER mcon ;
      RECT 0.120000  0.395000 0.290000 0.565000 ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.480000  0.395000 0.650000 0.565000 ;
      RECT 0.560000  3.505000 0.730000 3.675000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.920000  3.505000 1.090000 3.675000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.280000  3.505000 1.450000 3.675000 ;
      RECT 1.340000  0.395000 1.510000 0.565000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.640000  3.505000 1.810000 3.675000 ;
      RECT 1.700000  0.395000 1.870000 0.565000 ;
      RECT 2.000000  3.505000 2.170000 3.675000 ;
      RECT 2.060000  0.395000 2.230000 0.565000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.360000  3.505000 2.530000 3.675000 ;
      RECT 2.420000  0.395000 2.590000 0.565000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 2.780000  0.395000 2.950000 0.565000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
      RECT 3.085000  3.505000 3.255000 3.675000 ;
      RECT 3.140000  0.395000 3.310000 0.565000 ;
      RECT 3.445000  3.505000 3.615000 3.675000 ;
      RECT 3.500000  0.395000 3.670000 0.565000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.985000 3.685000 4.155000 ;
      RECT 3.805000  3.505000 3.975000 3.675000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.985000 4.165000 4.155000 ;
      RECT 4.165000  3.505000 4.335000 3.675000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.985000 4.645000 4.155000 ;
      RECT 4.525000  3.505000 4.695000 3.675000 ;
      RECT 4.580000  0.395000 4.750000 0.565000 ;
      RECT 4.940000  0.395000 5.110000 0.565000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.985000 5.125000 4.155000 ;
  END
END sky130_fd_sc_hvl__xor2_1
MACRO sky130_fd_sc_hvl__lsbufhv2lv_simple_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__lsbufhv2lv_simple_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  8.140000 ;
  SYMMETRY X Y ;
  SITE unithvdbl ;
  PIN A
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.355000 1.465000 4.685000 3.260000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.626250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.995000 0.495000 3.255000 2.175000 ;
        RECT 2.995000 2.175000 3.440000 3.755000 ;
    END
  END X
  PIN LVPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.070000 3.020000 8.570000 3.305000 ;
      LAYER nwell ;
        RECT 2.800000 1.885000 5.425000 4.825000 ;
    END
  END LVPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 7.515000 8.640000 7.885000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 8.025000 8.640000 8.255000 ;
      LAYER pwell ;
        RECT 0.000000 8.055000 8.640000 8.225000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 8.640000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 0.800000 6.255000 ;
        RECT  7.425000 1.885000 8.970000 6.255000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 4.325000 8.640000 4.695000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.640000 0.085000 ;
      RECT 0.000000  3.985000 0.800000 4.155000 ;
      RECT 0.000000  8.055000 8.640000 8.225000 ;
      RECT 3.130000  3.955000 5.095000 4.525000 ;
      RECT 3.435000  0.365000 4.685000 0.935000 ;
      RECT 3.565000  1.115000 5.115000 1.285000 ;
      RECT 3.565000  1.285000 3.895000 1.745000 ;
      RECT 3.620000  2.175000 4.175000 3.955000 ;
      RECT 4.865000  0.495000 5.115000 1.115000 ;
      RECT 4.865000  1.285000 5.115000 3.005000 ;
      RECT 7.425000  3.985000 8.640000 4.155000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.155000  8.055000 0.325000 8.225000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  8.055000 0.805000 8.225000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  8.055000 1.285000 8.225000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  8.055000 1.765000 8.225000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  8.055000 2.245000 8.225000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  8.055000 2.725000 8.225000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  8.055000 3.205000 8.225000 ;
      RECT 3.435000  0.395000 3.605000 0.565000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  8.055000 3.685000 8.225000 ;
      RECT 3.630000  3.075000 3.800000 3.245000 ;
      RECT 3.795000  0.395000 3.965000 0.565000 ;
      RECT 3.990000  3.075000 4.160000 3.245000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  8.055000 4.165000 8.225000 ;
      RECT 4.155000  0.395000 4.325000 0.565000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  8.055000 4.645000 8.225000 ;
      RECT 4.515000  0.395000 4.685000 0.565000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  8.055000 5.125000 8.225000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  8.055000 5.605000 8.225000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  8.055000 6.085000 8.225000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  8.055000 6.565000 8.225000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  8.055000 7.045000 8.225000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  8.055000 7.525000 8.225000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.985000 8.005000 4.155000 ;
      RECT 7.835000  8.055000 8.005000 8.225000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.985000 8.485000 4.155000 ;
      RECT 8.315000  8.055000 8.485000 8.225000 ;
    LAYER met1 ;
      RECT 0.000000 -0.115000 8.640000 0.115000 ;
      RECT 0.000000  0.255000 8.640000 0.625000 ;
      RECT 0.000000  3.445000 8.640000 3.815000 ;
    LAYER pwell ;
      RECT 0.000000 -0.085000 8.640000 0.085000 ;
  END
END sky130_fd_sc_hvl__lsbufhv2lv_simple_1
MACRO sky130_fd_sc_hvl__a21oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__a21oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A1
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.505000 1.915000 1.750000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.505000 1.315000 1.750000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.470000 1.805000 2.800000 3.260000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.832500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.220000 0.495000 2.470000 1.455000 ;
        RECT 2.220000 1.455000 3.235000 1.625000 ;
        RECT 2.980000 1.625000 3.235000 3.755000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 3.360000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 3.360000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 3.360000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 3.360000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 3.690000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 3.360000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.985000 3.360000 4.155000 ;
      RECT 0.260000  1.930000 2.290000 2.100000 ;
      RECT 0.260000  2.100000 0.510000 3.755000 ;
      RECT 0.330000  0.365000 2.040000 1.325000 ;
      RECT 0.690000  2.280000 1.940000 3.755000 ;
      RECT 2.120000  2.100000 2.290000 3.755000 ;
      RECT 2.675000  0.365000 3.265000 1.275000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.380000  0.395000 0.550000 0.565000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.690000  3.505000 0.860000 3.675000 ;
      RECT 0.740000  0.395000 0.910000 0.565000 ;
      RECT 1.050000  3.505000 1.220000 3.675000 ;
      RECT 1.100000  0.395000 1.270000 0.565000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.410000  3.505000 1.580000 3.675000 ;
      RECT 1.460000  0.395000 1.630000 0.565000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.770000  3.505000 1.940000 3.675000 ;
      RECT 1.820000  0.395000 1.990000 0.565000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 2.705000  0.395000 2.875000 0.565000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
      RECT 3.065000  0.395000 3.235000 0.565000 ;
  END
END sky130_fd_sc_hvl__a21oi_1
MACRO sky130_fd_sc_hvl__buf_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__buf_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.400000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 1.465000 1.795000 3.260000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.626250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.495000 0.365000 2.175000 ;
        RECT 0.115000 2.175000 0.550000 3.755000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 2.400000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 2.400000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 2.400000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 2.400000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 2.730000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 2.400000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.400000 0.085000 ;
      RECT 0.000000  3.985000 2.400000 4.155000 ;
      RECT 0.545000  0.365000 1.795000 0.935000 ;
      RECT 0.675000  1.115000 2.225000 1.285000 ;
      RECT 0.675000  1.285000 1.005000 1.745000 ;
      RECT 0.730000  2.175000 1.285000 3.755000 ;
      RECT 1.975000  0.495000 2.225000 1.115000 ;
      RECT 1.975000  1.285000 2.225000 3.005000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.545000  0.395000 0.715000 0.565000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.740000  3.505000 0.910000 3.675000 ;
      RECT 0.905000  0.395000 1.075000 0.565000 ;
      RECT 1.100000  3.505000 1.270000 3.675000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.265000  0.395000 1.435000 0.565000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.625000  0.395000 1.795000 0.565000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
  END
END sky130_fd_sc_hvl__buf_1
MACRO sky130_fd_sc_hvl__buf_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__buf_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.885000 1.775000 4.215000 2.120000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.260000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.550000 1.390000 1.780000 ;
        RECT 1.220000 0.495000 1.470000 1.205000 ;
        RECT 1.220000 1.205000 3.030000 1.375000 ;
        RECT 1.220000 1.375000 1.390000 1.550000 ;
        RECT 1.220000 1.780000 1.390000 1.905000 ;
        RECT 1.220000 1.905000 3.110000 2.075000 ;
        RECT 1.220000 2.075000 1.470000 3.755000 ;
        RECT 2.780000 0.495000 3.030000 1.205000 ;
        RECT 2.780000 2.075000 3.110000 3.755000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 4.800000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 4.800000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 4.800000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 4.800000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 5.130000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 4.800000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.985000 4.800000 4.155000 ;
      RECT 0.090000  0.365000 1.040000 1.325000 ;
      RECT 0.090000  2.175000 1.040000 3.755000 ;
      RECT 1.570000  1.555000 4.670000 1.595000 ;
      RECT 1.570000  1.595000 3.600000 1.725000 ;
      RECT 1.650000  0.365000 2.600000 1.025000 ;
      RECT 1.650000  2.255000 2.600000 3.755000 ;
      RECT 3.210000  0.365000 4.160000 1.245000 ;
      RECT 3.290000  2.300000 4.240000 3.755000 ;
      RECT 3.430000  1.425000 4.670000 1.555000 ;
      RECT 4.340000  0.495000 4.670000 1.425000 ;
      RECT 4.420000  1.595000 4.670000 3.755000 ;
    LAYER mcon ;
      RECT 0.120000  0.395000 0.290000 0.565000 ;
      RECT 0.120000  3.505000 0.290000 3.675000 ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.480000  0.395000 0.650000 0.565000 ;
      RECT 0.480000  3.505000 0.650000 3.675000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.840000  0.395000 1.010000 0.565000 ;
      RECT 0.840000  3.505000 1.010000 3.675000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.680000  0.395000 1.850000 0.565000 ;
      RECT 1.680000  3.505000 1.850000 3.675000 ;
      RECT 2.040000  0.395000 2.210000 0.565000 ;
      RECT 2.040000  3.505000 2.210000 3.675000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.400000  0.395000 2.570000 0.565000 ;
      RECT 2.400000  3.505000 2.570000 3.675000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
      RECT 3.240000  0.395000 3.410000 0.565000 ;
      RECT 3.320000  3.505000 3.490000 3.675000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.985000 3.685000 4.155000 ;
      RECT 3.600000  0.395000 3.770000 0.565000 ;
      RECT 3.680000  3.505000 3.850000 3.675000 ;
      RECT 3.960000  0.395000 4.130000 0.565000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.985000 4.165000 4.155000 ;
      RECT 4.040000  3.505000 4.210000 3.675000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.985000 4.645000 4.155000 ;
  END
END sky130_fd_sc_hvl__buf_4
MACRO sky130_fd_sc_hvl__buf_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__buf_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.600000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  3.375000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.635000 1.580000 2.245000 1.815000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  2.520000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.605000 2.035000 8.965000 2.205000 ;
        RECT 3.605000 2.205000 3.935000 3.445000 ;
        RECT 3.665000 0.805000 3.875000 1.625000 ;
        RECT 3.665000 1.625000 8.555000 1.795000 ;
        RECT 5.165000 2.205000 5.495000 3.445000 ;
        RECT 5.225000 0.805000 5.435000 1.625000 ;
        RECT 6.725000 2.205000 7.055000 3.445000 ;
        RECT 6.785000 0.805000 6.995000 1.625000 ;
        RECT 8.285000 2.205000 8.965000 3.230000 ;
        RECT 8.285000 3.230000 8.735000 3.445000 ;
        RECT 8.345000 0.805000 8.965000 0.975000 ;
        RECT 8.345000 0.975000 8.555000 1.625000 ;
        RECT 8.735000 0.975000 8.965000 2.035000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 9.600000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 9.600000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 9.600000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 9.600000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 9.930000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 9.600000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.600000 0.085000 ;
      RECT 0.000000  3.985000 9.600000 4.155000 ;
      RECT 0.245000  0.805000 0.455000 1.475000 ;
      RECT 0.245000  1.475000 0.435000 2.095000 ;
      RECT 0.245000  2.095000 2.595000 2.265000 ;
      RECT 0.245000  2.265000 0.435000 3.545000 ;
      RECT 0.615000  2.445000 1.865000 3.625000 ;
      RECT 0.615000  3.625000 9.505000 3.795000 ;
      RECT 0.675000  0.380000 9.505000 0.550000 ;
      RECT 0.675000  0.550000 1.925000 1.385000 ;
      RECT 2.045000  2.265000 2.595000 3.445000 ;
      RECT 2.105000  0.730000 2.315000 1.230000 ;
      RECT 2.105000  1.230000 2.595000 1.400000 ;
      RECT 2.425000  1.400000 2.595000 1.625000 ;
      RECT 2.425000  1.625000 3.380000 1.955000 ;
      RECT 2.425000  1.955000 2.595000 2.095000 ;
      RECT 2.605000  0.550000 3.495000 0.760000 ;
      RECT 2.765000  0.760000 3.495000 1.445000 ;
      RECT 2.765000  2.385000 3.435000 3.625000 ;
      RECT 4.045000  0.550000 5.055000 1.445000 ;
      RECT 4.105000  2.385000 4.995000 3.625000 ;
      RECT 5.605000  0.550000 6.615000 1.445000 ;
      RECT 5.665000  2.385000 6.555000 3.625000 ;
      RECT 7.165000  0.550000 8.175000 1.445000 ;
      RECT 7.225000  2.385000 8.115000 3.625000 ;
      RECT 8.905000  3.475000 9.505000 3.625000 ;
      RECT 8.975000  0.550000 9.505000 0.600000 ;
      RECT 9.135000  0.600000 9.505000 1.445000 ;
      RECT 9.135000  2.385000 9.505000 3.475000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.615000  3.475000 0.785000 3.645000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.975000  3.475000 1.145000 3.645000 ;
      RECT 1.035000  0.380000 1.205000 0.550000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.335000  3.475000 1.505000 3.645000 ;
      RECT 1.395000  0.380000 1.565000 0.550000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.695000  3.475000 1.865000 3.645000 ;
      RECT 1.755000  0.380000 1.925000 0.550000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 2.605000  0.380000 2.775000 0.550000 ;
      RECT 2.770000  3.475000 2.940000 3.645000 ;
      RECT 2.965000  0.380000 3.135000 0.550000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
      RECT 3.130000  3.475000 3.300000 3.645000 ;
      RECT 3.325000  0.380000 3.495000 0.550000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.985000 3.685000 4.155000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.985000 4.165000 4.155000 ;
      RECT 4.070000  0.380000 4.240000 0.550000 ;
      RECT 4.105000  3.475000 4.275000 3.645000 ;
      RECT 4.430000  0.380000 4.600000 0.550000 ;
      RECT 4.465000  3.475000 4.635000 3.645000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.985000 4.645000 4.155000 ;
      RECT 4.790000  0.380000 4.960000 0.550000 ;
      RECT 4.825000  3.475000 4.995000 3.645000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.985000 5.125000 4.155000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.985000 5.605000 4.155000 ;
      RECT 5.665000  3.475000 5.835000 3.645000 ;
      RECT 5.670000  0.380000 5.840000 0.550000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.985000 6.085000 4.155000 ;
      RECT 6.025000  3.475000 6.195000 3.645000 ;
      RECT 6.030000  0.380000 6.200000 0.550000 ;
      RECT 6.385000  3.475000 6.555000 3.645000 ;
      RECT 6.390000  0.380000 6.560000 0.550000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.985000 6.565000 4.155000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.985000 7.045000 4.155000 ;
      RECT 7.230000  3.475000 7.400000 3.645000 ;
      RECT 7.235000  0.380000 7.405000 0.550000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.985000 7.525000 4.155000 ;
      RECT 7.595000  0.380000 7.765000 0.550000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.985000 8.005000 4.155000 ;
      RECT 7.945000  3.475000 8.115000 3.645000 ;
      RECT 7.955000  0.380000 8.125000 0.550000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.985000 8.485000 4.155000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.985000 8.965000 4.155000 ;
      RECT 8.975000  0.380000 9.145000 0.550000 ;
      RECT 9.265000  3.475000 9.435000 3.645000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.985000 9.445000 4.155000 ;
      RECT 9.335000  0.380000 9.505000 0.550000 ;
  END
END sky130_fd_sc_hvl__buf_8
MACRO sky130_fd_sc_hvl__buf_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__buf_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  17.76000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  6.750000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.220000 1.580000 4.630000 1.815000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  5.040000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  5.590000 2.290000  5.880000 2.320000 ;
        RECT  5.590000 2.320000 16.800000 2.490000 ;
        RECT  5.590000 2.490000  5.880000 2.520000 ;
        RECT  7.150000 2.290000  7.440000 2.320000 ;
        RECT  7.150000 2.490000  7.440000 2.520000 ;
        RECT  8.710000 2.290000  9.000000 2.320000 ;
        RECT  8.710000 2.490000  9.000000 2.520000 ;
        RECT 10.270000 2.290000 10.560000 2.320000 ;
        RECT 10.270000 2.490000 10.560000 2.520000 ;
        RECT 11.830000 2.290000 12.120000 2.320000 ;
        RECT 11.830000 2.490000 12.120000 2.520000 ;
        RECT 13.390000 2.290000 13.680000 2.320000 ;
        RECT 13.390000 2.490000 13.680000 2.520000 ;
        RECT 14.950000 2.290000 15.240000 2.320000 ;
        RECT 14.950000 2.490000 15.240000 2.520000 ;
        RECT 16.510000 2.290000 16.800000 2.320000 ;
        RECT 16.510000 2.490000 16.800000 2.520000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 17.760000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 17.760000 0.085000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
        RECT 13.595000 -0.085000 13.765000 0.085000 ;
        RECT 14.075000 -0.085000 14.245000 0.085000 ;
        RECT 14.555000 -0.085000 14.725000 0.085000 ;
        RECT 15.035000 -0.085000 15.205000 0.085000 ;
        RECT 15.515000 -0.085000 15.685000 0.085000 ;
        RECT 15.995000 -0.085000 16.165000 0.085000 ;
        RECT 16.475000 -0.085000 16.645000 0.085000 ;
        RECT 16.955000 -0.085000 17.125000 0.085000 ;
        RECT 17.435000 -0.085000 17.605000 0.085000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 17.760000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 17.760000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.985000 17.760000 4.155000 ;
      LAYER mcon ;
        RECT  0.155000 3.985000  0.325000 4.155000 ;
        RECT  0.635000 3.985000  0.805000 4.155000 ;
        RECT  1.115000 3.985000  1.285000 4.155000 ;
        RECT  1.595000 3.985000  1.765000 4.155000 ;
        RECT  2.075000 3.985000  2.245000 4.155000 ;
        RECT  2.555000 3.985000  2.725000 4.155000 ;
        RECT  3.035000 3.985000  3.205000 4.155000 ;
        RECT  3.515000 3.985000  3.685000 4.155000 ;
        RECT  3.995000 3.985000  4.165000 4.155000 ;
        RECT  4.475000 3.985000  4.645000 4.155000 ;
        RECT  4.955000 3.985000  5.125000 4.155000 ;
        RECT  5.435000 3.985000  5.605000 4.155000 ;
        RECT  5.915000 3.985000  6.085000 4.155000 ;
        RECT  6.395000 3.985000  6.565000 4.155000 ;
        RECT  6.875000 3.985000  7.045000 4.155000 ;
        RECT  7.355000 3.985000  7.525000 4.155000 ;
        RECT  7.835000 3.985000  8.005000 4.155000 ;
        RECT  8.315000 3.985000  8.485000 4.155000 ;
        RECT  8.795000 3.985000  8.965000 4.155000 ;
        RECT  9.275000 3.985000  9.445000 4.155000 ;
        RECT  9.755000 3.985000  9.925000 4.155000 ;
        RECT 10.235000 3.985000 10.405000 4.155000 ;
        RECT 10.715000 3.985000 10.885000 4.155000 ;
        RECT 11.195000 3.985000 11.365000 4.155000 ;
        RECT 11.675000 3.985000 11.845000 4.155000 ;
        RECT 12.155000 3.985000 12.325000 4.155000 ;
        RECT 12.635000 3.985000 12.805000 4.155000 ;
        RECT 13.115000 3.985000 13.285000 4.155000 ;
        RECT 13.595000 3.985000 13.765000 4.155000 ;
        RECT 14.075000 3.985000 14.245000 4.155000 ;
        RECT 14.555000 3.985000 14.725000 4.155000 ;
        RECT 15.035000 3.985000 15.205000 4.155000 ;
        RECT 15.515000 3.985000 15.685000 4.155000 ;
        RECT 15.995000 3.985000 16.165000 4.155000 ;
        RECT 16.475000 3.985000 16.645000 4.155000 ;
        RECT 16.955000 3.985000 17.125000 4.155000 ;
        RECT 17.435000 3.985000 17.605000 4.155000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 17.760000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 18.090000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 17.760000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.110000 0.425000  0.645000 1.410000 ;
      RECT  0.110000 2.175000  0.680000 3.755000 ;
      RECT  0.815000 0.755000  1.170000 1.195000 ;
      RECT  0.815000 1.195000  5.350000 1.410000 ;
      RECT  0.850000 1.985000  5.350000 2.265000 ;
      RECT  0.850000 2.265000  1.160000 3.755000 ;
      RECT  1.340000 0.415000  2.230000 1.025000 ;
      RECT  1.340000 2.445000  2.230000 3.675000 ;
      RECT  2.400000 0.730000  2.790000 1.195000 ;
      RECT  2.400000 2.265000  2.710000 3.755000 ;
      RECT  2.880000 2.445000  3.770000 3.675000 ;
      RECT  2.960000 0.425000  3.855000 1.025000 ;
      RECT  3.940000 2.265000  4.290000 3.755000 ;
      RECT  4.025000 0.730000  4.270000 1.195000 ;
      RECT  4.440000 0.425000  5.330000 1.025000 ;
      RECT  4.460000 2.445000  5.350000 3.675000 ;
      RECT  4.800000 1.410000  5.350000 1.985000 ;
      RECT  5.570000 0.790000  5.900000 3.755000 ;
      RECT  6.070000 0.425000  6.960000 1.395000 ;
      RECT  6.070000 2.175000  6.960000 3.755000 ;
      RECT  6.160000 1.565000  6.830000 1.895000 ;
      RECT  7.130000 0.790000  7.460000 3.755000 ;
      RECT  7.630000 0.425000  8.520000 1.395000 ;
      RECT  7.630000 2.175000  8.520000 3.755000 ;
      RECT  7.720000 1.565000  8.390000 1.895000 ;
      RECT  8.690000 0.790000  9.020000 3.755000 ;
      RECT  9.190000 0.425000 10.080000 1.395000 ;
      RECT  9.190000 2.175000 10.080000 3.755000 ;
      RECT  9.280000 1.565000  9.950000 1.895000 ;
      RECT 10.250000 0.790000 10.580000 3.755000 ;
      RECT 10.750000 0.425000 11.640000 1.395000 ;
      RECT 10.750000 2.175000 11.640000 3.755000 ;
      RECT 10.840000 1.565000 11.510000 1.895000 ;
      RECT 11.810000 0.790000 12.140000 3.755000 ;
      RECT 12.310000 0.425000 13.200000 1.395000 ;
      RECT 12.310000 2.175000 13.200000 3.755000 ;
      RECT 12.400000 1.565000 13.070000 1.895000 ;
      RECT 13.370000 0.790000 13.700000 3.755000 ;
      RECT 13.870000 0.425000 14.760000 1.395000 ;
      RECT 13.870000 2.175000 14.760000 3.755000 ;
      RECT 13.960000 1.565000 14.630000 1.895000 ;
      RECT 14.930000 0.790000 15.260000 3.755000 ;
      RECT 15.430000 0.425000 16.320000 1.395000 ;
      RECT 15.430000 2.175000 16.320000 3.755000 ;
      RECT 15.520000 1.565000 16.190000 1.895000 ;
      RECT 16.490000 0.790000 16.900000 3.755000 ;
      RECT 17.070000 0.425000 17.600000 1.495000 ;
      RECT 17.070000 2.175000 17.600000 3.755000 ;
    LAYER mcon ;
      RECT  0.115000 0.425000  0.285000 0.595000 ;
      RECT  0.150000 3.475000  0.320000 3.645000 ;
      RECT  0.475000 0.425000  0.645000 0.595000 ;
      RECT  0.510000 3.475000  0.680000 3.645000 ;
      RECT  1.340000 0.425000  1.510000 0.595000 ;
      RECT  1.340000 3.475000  1.510000 3.645000 ;
      RECT  1.700000 0.425000  1.870000 0.595000 ;
      RECT  1.700000 3.475000  1.870000 3.645000 ;
      RECT  2.060000 0.425000  2.230000 0.595000 ;
      RECT  2.060000 3.475000  2.230000 3.645000 ;
      RECT  2.880000 3.475000  3.050000 3.645000 ;
      RECT  3.240000 3.475000  3.410000 3.645000 ;
      RECT  3.320000 0.425000  3.490000 0.595000 ;
      RECT  3.600000 3.475000  3.770000 3.645000 ;
      RECT  3.680000 0.425000  3.850000 0.595000 ;
      RECT  4.460000 3.475000  4.630000 3.645000 ;
      RECT  4.800000 0.425000  4.970000 0.595000 ;
      RECT  4.800000 1.580000  4.970000 1.750000 ;
      RECT  4.820000 3.475000  4.990000 3.645000 ;
      RECT  5.160000 0.425000  5.330000 0.595000 ;
      RECT  5.160000 1.580000  5.330000 1.750000 ;
      RECT  5.180000 3.475000  5.350000 3.645000 ;
      RECT  5.650000 2.320000  5.820000 2.490000 ;
      RECT  6.070000 3.475000  6.240000 3.645000 ;
      RECT  6.230000 1.580000  6.400000 1.750000 ;
      RECT  6.430000 0.425000  6.600000 0.595000 ;
      RECT  6.430000 3.475000  6.600000 3.645000 ;
      RECT  6.590000 1.580000  6.760000 1.750000 ;
      RECT  6.790000 0.425000  6.960000 0.595000 ;
      RECT  6.790000 3.475000  6.960000 3.645000 ;
      RECT  7.210000 2.320000  7.380000 2.490000 ;
      RECT  7.630000 3.475000  7.800000 3.645000 ;
      RECT  7.790000 1.580000  7.960000 1.750000 ;
      RECT  7.990000 0.425000  8.160000 0.595000 ;
      RECT  7.990000 3.475000  8.160000 3.645000 ;
      RECT  8.150000 1.580000  8.320000 1.750000 ;
      RECT  8.350000 0.425000  8.520000 0.595000 ;
      RECT  8.350000 3.475000  8.520000 3.645000 ;
      RECT  8.770000 2.320000  8.940000 2.490000 ;
      RECT  9.190000 3.475000  9.360000 3.645000 ;
      RECT  9.350000 1.580000  9.520000 1.750000 ;
      RECT  9.550000 0.425000  9.720000 0.595000 ;
      RECT  9.550000 3.475000  9.720000 3.645000 ;
      RECT  9.710000 1.580000  9.880000 1.750000 ;
      RECT  9.910000 0.425000 10.080000 0.595000 ;
      RECT  9.910000 3.475000 10.080000 3.645000 ;
      RECT 10.330000 2.320000 10.500000 2.490000 ;
      RECT 10.750000 3.475000 10.920000 3.645000 ;
      RECT 10.910000 1.580000 11.080000 1.750000 ;
      RECT 11.110000 0.425000 11.280000 0.595000 ;
      RECT 11.110000 3.475000 11.280000 3.645000 ;
      RECT 11.270000 1.580000 11.440000 1.750000 ;
      RECT 11.470000 0.425000 11.640000 0.595000 ;
      RECT 11.470000 3.475000 11.640000 3.645000 ;
      RECT 11.890000 2.320000 12.060000 2.490000 ;
      RECT 12.310000 3.475000 12.480000 3.645000 ;
      RECT 12.470000 1.580000 12.640000 1.750000 ;
      RECT 12.670000 0.425000 12.840000 0.595000 ;
      RECT 12.670000 3.475000 12.840000 3.645000 ;
      RECT 12.830000 1.580000 13.000000 1.750000 ;
      RECT 13.030000 0.425000 13.200000 0.595000 ;
      RECT 13.030000 3.475000 13.200000 3.645000 ;
      RECT 13.450000 2.320000 13.620000 2.490000 ;
      RECT 13.870000 3.475000 14.040000 3.645000 ;
      RECT 14.030000 1.580000 14.200000 1.750000 ;
      RECT 14.230000 0.425000 14.400000 0.595000 ;
      RECT 14.230000 3.475000 14.400000 3.645000 ;
      RECT 14.390000 1.580000 14.560000 1.750000 ;
      RECT 14.590000 0.425000 14.760000 0.595000 ;
      RECT 14.590000 3.475000 14.760000 3.645000 ;
      RECT 15.010000 2.320000 15.180000 2.490000 ;
      RECT 15.430000 3.475000 15.600000 3.645000 ;
      RECT 15.590000 1.580000 15.760000 1.750000 ;
      RECT 15.790000 0.425000 15.960000 0.595000 ;
      RECT 15.790000 3.475000 15.960000 3.645000 ;
      RECT 15.950000 1.580000 16.120000 1.750000 ;
      RECT 16.150000 0.425000 16.320000 0.595000 ;
      RECT 16.150000 3.475000 16.320000 3.645000 ;
      RECT 16.570000 2.320000 16.740000 2.490000 ;
      RECT 17.070000 3.475000 17.240000 3.645000 ;
      RECT 17.430000 0.425000 17.600000 0.595000 ;
      RECT 17.430000 3.475000 17.600000 3.645000 ;
    LAYER met1 ;
      RECT  4.740000 1.550000  5.360000 1.580000 ;
      RECT  4.740000 1.580000 16.250000 1.750000 ;
      RECT  4.740000 1.750000  5.360000 1.780000 ;
      RECT  6.170000 1.550000  6.820000 1.580000 ;
      RECT  6.170000 1.750000  6.820000 1.780000 ;
      RECT  7.730000 1.550000  8.380000 1.580000 ;
      RECT  7.730000 1.750000  8.380000 1.780000 ;
      RECT  9.290000 1.550000  9.940000 1.580000 ;
      RECT  9.290000 1.750000  9.940000 1.780000 ;
      RECT 10.850000 1.550000 11.500000 1.580000 ;
      RECT 10.850000 1.750000 11.500000 1.780000 ;
      RECT 12.410000 1.550000 13.060000 1.580000 ;
      RECT 12.410000 1.750000 13.060000 1.780000 ;
      RECT 13.970000 1.550000 14.620000 1.580000 ;
      RECT 13.970000 1.750000 14.620000 1.780000 ;
      RECT 15.530000 1.550000 16.180000 1.580000 ;
      RECT 15.530000 1.750000 16.180000 1.780000 ;
  END
END sky130_fd_sc_hvl__buf_16
MACRO sky130_fd_sc_hvl__buf_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__buf_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.775000 2.775000 2.120000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.630000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.550000 1.390000 1.720000 ;
        RECT 0.125000 1.720000 1.370000 1.780000 ;
        RECT 1.200000 1.780000 1.370000 3.755000 ;
        RECT 1.220000 0.495000 1.390000 1.550000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 3.360000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 3.360000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 3.360000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 3.360000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 3.690000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 3.360000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.985000 3.360000 4.155000 ;
      RECT 0.090000  0.365000 1.040000 1.325000 ;
      RECT 0.090000  2.175000 1.020000 3.755000 ;
      RECT 1.550000  2.300000 2.800000 3.755000 ;
      RECT 1.570000  0.365000 2.820000 1.245000 ;
      RECT 1.570000  1.425000 3.250000 1.595000 ;
      RECT 1.570000  1.595000 1.865000 1.755000 ;
      RECT 2.980000  1.595000 3.250000 3.005000 ;
      RECT 3.000000  0.825000 3.250000 1.425000 ;
    LAYER mcon ;
      RECT 0.110000  3.505000 0.280000 3.675000 ;
      RECT 0.120000  0.395000 0.290000 0.565000 ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.470000  3.505000 0.640000 3.675000 ;
      RECT 0.480000  0.395000 0.650000 0.565000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.830000  3.505000 1.000000 3.675000 ;
      RECT 0.840000  0.395000 1.010000 0.565000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.550000  3.505000 1.720000 3.675000 ;
      RECT 1.570000  0.395000 1.740000 0.565000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.910000  3.505000 2.080000 3.675000 ;
      RECT 1.930000  0.395000 2.100000 0.565000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.270000  3.505000 2.440000 3.675000 ;
      RECT 2.290000  0.395000 2.460000 0.565000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 2.630000  3.505000 2.800000 3.675000 ;
      RECT 2.650000  0.395000 2.820000 0.565000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
  END
END sky130_fd_sc_hvl__buf_2
MACRO sky130_fd_sc_hvl__buf_32
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__buf_32 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  33.60000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  11.25000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.220000 1.580000 4.630000 1.815000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  10.08000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 8.950000 2.290000 32.640000 2.520000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 33.600000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 33.600000 0.085000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
        RECT 13.595000 -0.085000 13.765000 0.085000 ;
        RECT 14.075000 -0.085000 14.245000 0.085000 ;
        RECT 14.555000 -0.085000 14.725000 0.085000 ;
        RECT 15.035000 -0.085000 15.205000 0.085000 ;
        RECT 15.515000 -0.085000 15.685000 0.085000 ;
        RECT 15.995000 -0.085000 16.165000 0.085000 ;
        RECT 16.475000 -0.085000 16.645000 0.085000 ;
        RECT 16.955000 -0.085000 17.125000 0.085000 ;
        RECT 17.435000 -0.085000 17.605000 0.085000 ;
        RECT 17.915000 -0.085000 18.085000 0.085000 ;
        RECT 18.395000 -0.085000 18.565000 0.085000 ;
        RECT 18.875000 -0.085000 19.045000 0.085000 ;
        RECT 19.355000 -0.085000 19.525000 0.085000 ;
        RECT 19.835000 -0.085000 20.005000 0.085000 ;
        RECT 20.315000 -0.085000 20.485000 0.085000 ;
        RECT 20.795000 -0.085000 20.965000 0.085000 ;
        RECT 21.275000 -0.085000 21.445000 0.085000 ;
        RECT 21.755000 -0.085000 21.925000 0.085000 ;
        RECT 22.235000 -0.085000 22.405000 0.085000 ;
        RECT 22.715000 -0.085000 22.885000 0.085000 ;
        RECT 23.195000 -0.085000 23.365000 0.085000 ;
        RECT 23.675000 -0.085000 23.845000 0.085000 ;
        RECT 24.155000 -0.085000 24.325000 0.085000 ;
        RECT 24.635000 -0.085000 24.805000 0.085000 ;
        RECT 25.115000 -0.085000 25.285000 0.085000 ;
        RECT 25.595000 -0.085000 25.765000 0.085000 ;
        RECT 26.075000 -0.085000 26.245000 0.085000 ;
        RECT 26.555000 -0.085000 26.725000 0.085000 ;
        RECT 27.035000 -0.085000 27.205000 0.085000 ;
        RECT 27.515000 -0.085000 27.685000 0.085000 ;
        RECT 27.995000 -0.085000 28.165000 0.085000 ;
        RECT 28.475000 -0.085000 28.645000 0.085000 ;
        RECT 28.955000 -0.085000 29.125000 0.085000 ;
        RECT 29.435000 -0.085000 29.605000 0.085000 ;
        RECT 29.915000 -0.085000 30.085000 0.085000 ;
        RECT 30.395000 -0.085000 30.565000 0.085000 ;
        RECT 30.875000 -0.085000 31.045000 0.085000 ;
        RECT 31.355000 -0.085000 31.525000 0.085000 ;
        RECT 31.835000 -0.085000 32.005000 0.085000 ;
        RECT 32.315000 -0.085000 32.485000 0.085000 ;
        RECT 32.795000 -0.085000 32.965000 0.085000 ;
        RECT 33.275000 -0.085000 33.445000 0.085000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 33.600000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 33.600000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.985000 33.600000 4.155000 ;
      LAYER mcon ;
        RECT  0.155000 3.985000  0.325000 4.155000 ;
        RECT  0.635000 3.985000  0.805000 4.155000 ;
        RECT  1.115000 3.985000  1.285000 4.155000 ;
        RECT  1.595000 3.985000  1.765000 4.155000 ;
        RECT  2.075000 3.985000  2.245000 4.155000 ;
        RECT  2.555000 3.985000  2.725000 4.155000 ;
        RECT  3.035000 3.985000  3.205000 4.155000 ;
        RECT  3.515000 3.985000  3.685000 4.155000 ;
        RECT  3.995000 3.985000  4.165000 4.155000 ;
        RECT  4.475000 3.985000  4.645000 4.155000 ;
        RECT  4.955000 3.985000  5.125000 4.155000 ;
        RECT  5.435000 3.985000  5.605000 4.155000 ;
        RECT  5.915000 3.985000  6.085000 4.155000 ;
        RECT  6.395000 3.985000  6.565000 4.155000 ;
        RECT  6.875000 3.985000  7.045000 4.155000 ;
        RECT  7.355000 3.985000  7.525000 4.155000 ;
        RECT  7.835000 3.985000  8.005000 4.155000 ;
        RECT  8.315000 3.985000  8.485000 4.155000 ;
        RECT  8.795000 3.985000  8.965000 4.155000 ;
        RECT  9.275000 3.985000  9.445000 4.155000 ;
        RECT  9.755000 3.985000  9.925000 4.155000 ;
        RECT 10.235000 3.985000 10.405000 4.155000 ;
        RECT 10.715000 3.985000 10.885000 4.155000 ;
        RECT 11.195000 3.985000 11.365000 4.155000 ;
        RECT 11.675000 3.985000 11.845000 4.155000 ;
        RECT 12.155000 3.985000 12.325000 4.155000 ;
        RECT 12.635000 3.985000 12.805000 4.155000 ;
        RECT 13.115000 3.985000 13.285000 4.155000 ;
        RECT 13.595000 3.985000 13.765000 4.155000 ;
        RECT 14.075000 3.985000 14.245000 4.155000 ;
        RECT 14.555000 3.985000 14.725000 4.155000 ;
        RECT 15.035000 3.985000 15.205000 4.155000 ;
        RECT 15.515000 3.985000 15.685000 4.155000 ;
        RECT 15.995000 3.985000 16.165000 4.155000 ;
        RECT 16.475000 3.985000 16.645000 4.155000 ;
        RECT 16.955000 3.985000 17.125000 4.155000 ;
        RECT 17.435000 3.985000 17.605000 4.155000 ;
        RECT 17.915000 3.985000 18.085000 4.155000 ;
        RECT 18.395000 3.985000 18.565000 4.155000 ;
        RECT 18.875000 3.985000 19.045000 4.155000 ;
        RECT 19.355000 3.985000 19.525000 4.155000 ;
        RECT 19.835000 3.985000 20.005000 4.155000 ;
        RECT 20.315000 3.985000 20.485000 4.155000 ;
        RECT 20.795000 3.985000 20.965000 4.155000 ;
        RECT 21.275000 3.985000 21.445000 4.155000 ;
        RECT 21.755000 3.985000 21.925000 4.155000 ;
        RECT 22.235000 3.985000 22.405000 4.155000 ;
        RECT 22.715000 3.985000 22.885000 4.155000 ;
        RECT 23.195000 3.985000 23.365000 4.155000 ;
        RECT 23.675000 3.985000 23.845000 4.155000 ;
        RECT 24.155000 3.985000 24.325000 4.155000 ;
        RECT 24.635000 3.985000 24.805000 4.155000 ;
        RECT 25.115000 3.985000 25.285000 4.155000 ;
        RECT 25.595000 3.985000 25.765000 4.155000 ;
        RECT 26.075000 3.985000 26.245000 4.155000 ;
        RECT 26.555000 3.985000 26.725000 4.155000 ;
        RECT 27.035000 3.985000 27.205000 4.155000 ;
        RECT 27.515000 3.985000 27.685000 4.155000 ;
        RECT 27.995000 3.985000 28.165000 4.155000 ;
        RECT 28.475000 3.985000 28.645000 4.155000 ;
        RECT 28.955000 3.985000 29.125000 4.155000 ;
        RECT 29.435000 3.985000 29.605000 4.155000 ;
        RECT 29.915000 3.985000 30.085000 4.155000 ;
        RECT 30.395000 3.985000 30.565000 4.155000 ;
        RECT 30.875000 3.985000 31.045000 4.155000 ;
        RECT 31.355000 3.985000 31.525000 4.155000 ;
        RECT 31.835000 3.985000 32.005000 4.155000 ;
        RECT 32.315000 3.985000 32.485000 4.155000 ;
        RECT 32.795000 3.985000 32.965000 4.155000 ;
        RECT 33.275000 3.985000 33.445000 4.155000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 33.600000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 33.930000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 33.600000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.110000 0.425000  0.645000 1.410000 ;
      RECT  0.110000 2.175000  0.680000 3.755000 ;
      RECT  0.815000 0.755000  1.170000 1.195000 ;
      RECT  0.815000 1.195000  7.410000 1.410000 ;
      RECT  0.850000 1.985000  7.410000 2.265000 ;
      RECT  0.850000 2.265000  1.160000 3.755000 ;
      RECT  1.340000 0.415000  2.230000 1.025000 ;
      RECT  1.340000 2.445000  2.230000 3.675000 ;
      RECT  2.400000 0.730000  2.790000 1.195000 ;
      RECT  2.400000 2.265000  2.710000 3.755000 ;
      RECT  2.880000 2.445000  3.770000 3.675000 ;
      RECT  2.960000 0.425000  3.855000 1.025000 ;
      RECT  3.940000 2.265000  4.290000 3.755000 ;
      RECT  4.025000 0.730000  4.270000 1.195000 ;
      RECT  4.440000 0.425000  5.330000 1.025000 ;
      RECT  4.460000 2.445000  5.350000 3.675000 ;
      RECT  4.800000 1.410000  7.410000 1.985000 ;
      RECT  5.520000 0.730000  5.910000 1.195000 ;
      RECT  5.520000 2.265000  5.830000 3.755000 ;
      RECT  6.000000 2.445000  6.890000 3.675000 ;
      RECT  6.080000 0.425000  6.975000 1.025000 ;
      RECT  7.060000 2.265000  7.410000 3.755000 ;
      RECT  7.145000 0.730000  7.390000 1.195000 ;
      RECT  7.560000 0.425000  8.480000 1.025000 ;
      RECT  7.580000 1.025000  8.480000 1.395000 ;
      RECT  7.580000 2.235000  8.480000 3.675000 ;
      RECT  8.930000 0.790000  9.260000 3.755000 ;
      RECT  9.430000 0.425000 10.320000 1.395000 ;
      RECT  9.430000 2.175000 10.320000 3.755000 ;
      RECT  9.520000 1.565000 10.190000 1.895000 ;
      RECT 10.490000 0.790000 10.820000 3.755000 ;
      RECT 10.990000 0.425000 11.880000 1.395000 ;
      RECT 10.990000 2.175000 11.880000 3.755000 ;
      RECT 11.080000 1.565000 11.750000 1.895000 ;
      RECT 12.050000 0.790000 12.380000 3.755000 ;
      RECT 12.550000 0.425000 13.440000 1.395000 ;
      RECT 12.550000 2.175000 13.440000 3.755000 ;
      RECT 12.640000 1.565000 13.310000 1.895000 ;
      RECT 13.610000 0.790000 13.940000 3.755000 ;
      RECT 14.110000 0.425000 15.000000 1.395000 ;
      RECT 14.110000 2.175000 15.000000 3.755000 ;
      RECT 14.200000 1.565000 14.870000 1.895000 ;
      RECT 15.170000 0.790000 15.500000 3.755000 ;
      RECT 15.670000 0.425000 16.560000 1.395000 ;
      RECT 15.670000 2.175000 16.560000 3.755000 ;
      RECT 15.760000 1.565000 16.430000 1.895000 ;
      RECT 16.730000 0.790000 17.060000 3.755000 ;
      RECT 17.230000 0.425000 18.120000 1.395000 ;
      RECT 17.230000 2.175000 18.120000 3.755000 ;
      RECT 17.320000 1.565000 17.990000 1.895000 ;
      RECT 18.290000 0.790000 18.620000 3.755000 ;
      RECT 18.790000 0.425000 19.680000 1.395000 ;
      RECT 18.790000 2.175000 19.680000 3.755000 ;
      RECT 18.880000 1.565000 19.550000 1.895000 ;
      RECT 19.850000 0.790000 20.260000 3.755000 ;
      RECT 20.430000 0.425000 20.960000 1.395000 ;
      RECT 20.430000 1.565000 21.100000 1.895000 ;
      RECT 20.430000 2.175000 20.960000 3.755000 ;
      RECT 21.410000 0.790000 21.740000 3.755000 ;
      RECT 21.910000 0.425000 22.800000 1.395000 ;
      RECT 21.910000 2.175000 22.800000 3.755000 ;
      RECT 22.000000 1.565000 22.670000 1.895000 ;
      RECT 22.970000 0.790000 23.300000 3.755000 ;
      RECT 23.470000 0.425000 24.360000 1.395000 ;
      RECT 23.470000 2.175000 24.360000 3.755000 ;
      RECT 23.560000 1.565000 24.230000 1.895000 ;
      RECT 24.530000 0.790000 24.860000 3.755000 ;
      RECT 25.030000 0.425000 25.920000 1.395000 ;
      RECT 25.030000 2.175000 25.920000 3.755000 ;
      RECT 25.120000 1.565000 25.790000 1.895000 ;
      RECT 26.090000 0.790000 26.420000 3.755000 ;
      RECT 26.590000 0.425000 27.480000 1.395000 ;
      RECT 26.590000 2.175000 27.480000 3.755000 ;
      RECT 26.680000 1.565000 27.350000 1.895000 ;
      RECT 27.650000 0.790000 27.980000 3.755000 ;
      RECT 28.150000 0.425000 29.040000 1.395000 ;
      RECT 28.150000 2.175000 29.040000 3.755000 ;
      RECT 28.240000 1.565000 28.910000 1.895000 ;
      RECT 29.210000 0.790000 29.540000 3.755000 ;
      RECT 29.710000 0.425000 30.600000 1.395000 ;
      RECT 29.710000 2.175000 30.600000 3.755000 ;
      RECT 29.800000 1.565000 30.470000 1.895000 ;
      RECT 30.770000 0.790000 31.100000 3.755000 ;
      RECT 31.270000 0.425000 32.160000 1.395000 ;
      RECT 31.270000 2.175000 32.160000 3.755000 ;
      RECT 31.360000 1.565000 32.030000 1.895000 ;
      RECT 32.330000 0.790000 32.740000 3.755000 ;
      RECT 32.910000 0.425000 33.440000 1.495000 ;
      RECT 32.910000 2.175000 33.440000 3.755000 ;
    LAYER mcon ;
      RECT  0.115000 0.425000  0.285000 0.595000 ;
      RECT  0.150000 3.475000  0.320000 3.645000 ;
      RECT  0.475000 0.425000  0.645000 0.595000 ;
      RECT  0.510000 3.475000  0.680000 3.645000 ;
      RECT  1.340000 0.425000  1.510000 0.595000 ;
      RECT  1.340000 3.475000  1.510000 3.645000 ;
      RECT  1.700000 0.425000  1.870000 0.595000 ;
      RECT  1.700000 3.475000  1.870000 3.645000 ;
      RECT  2.060000 0.425000  2.230000 0.595000 ;
      RECT  2.060000 3.475000  2.230000 3.645000 ;
      RECT  2.880000 3.475000  3.050000 3.645000 ;
      RECT  3.240000 3.475000  3.410000 3.645000 ;
      RECT  3.320000 0.425000  3.490000 0.595000 ;
      RECT  3.600000 3.475000  3.770000 3.645000 ;
      RECT  3.680000 0.425000  3.850000 0.595000 ;
      RECT  4.460000 3.475000  4.630000 3.645000 ;
      RECT  4.800000 0.425000  4.970000 0.595000 ;
      RECT  4.820000 3.475000  4.990000 3.645000 ;
      RECT  5.020000 1.580000  5.190000 1.750000 ;
      RECT  5.160000 0.425000  5.330000 0.595000 ;
      RECT  5.180000 3.475000  5.350000 3.645000 ;
      RECT  5.380000 1.580000  5.550000 1.750000 ;
      RECT  5.740000 1.580000  5.910000 1.750000 ;
      RECT  6.000000 3.475000  6.170000 3.645000 ;
      RECT  6.100000 1.580000  6.270000 1.750000 ;
      RECT  6.360000 3.475000  6.530000 3.645000 ;
      RECT  6.440000 0.425000  6.610000 0.595000 ;
      RECT  6.460000 1.580000  6.630000 1.750000 ;
      RECT  6.720000 3.475000  6.890000 3.645000 ;
      RECT  6.800000 0.425000  6.970000 0.595000 ;
      RECT  6.820000 1.580000  6.990000 1.750000 ;
      RECT  7.180000 1.580000  7.350000 1.750000 ;
      RECT  7.580000 3.475000  7.750000 3.645000 ;
      RECT  7.920000 0.425000  8.090000 0.595000 ;
      RECT  7.940000 3.475000  8.110000 3.645000 ;
      RECT  8.280000 0.425000  8.450000 0.595000 ;
      RECT  8.300000 3.475000  8.470000 3.645000 ;
      RECT  9.010000 2.320000  9.180000 2.490000 ;
      RECT  9.430000 3.475000  9.600000 3.645000 ;
      RECT  9.590000 1.580000  9.760000 1.750000 ;
      RECT  9.790000 0.425000  9.960000 0.595000 ;
      RECT  9.790000 3.475000  9.960000 3.645000 ;
      RECT  9.950000 1.580000 10.120000 1.750000 ;
      RECT 10.150000 0.425000 10.320000 0.595000 ;
      RECT 10.150000 3.475000 10.320000 3.645000 ;
      RECT 10.570000 2.320000 10.740000 2.490000 ;
      RECT 10.990000 3.475000 11.160000 3.645000 ;
      RECT 11.150000 1.580000 11.320000 1.750000 ;
      RECT 11.350000 0.425000 11.520000 0.595000 ;
      RECT 11.350000 3.475000 11.520000 3.645000 ;
      RECT 11.510000 1.580000 11.680000 1.750000 ;
      RECT 11.710000 0.425000 11.880000 0.595000 ;
      RECT 11.710000 3.475000 11.880000 3.645000 ;
      RECT 12.130000 2.320000 12.300000 2.490000 ;
      RECT 12.550000 3.475000 12.720000 3.645000 ;
      RECT 12.710000 1.580000 12.880000 1.750000 ;
      RECT 12.910000 0.425000 13.080000 0.595000 ;
      RECT 12.910000 3.475000 13.080000 3.645000 ;
      RECT 13.070000 1.580000 13.240000 1.750000 ;
      RECT 13.270000 0.425000 13.440000 0.595000 ;
      RECT 13.270000 3.475000 13.440000 3.645000 ;
      RECT 13.690000 2.320000 13.860000 2.490000 ;
      RECT 14.110000 3.475000 14.280000 3.645000 ;
      RECT 14.270000 1.580000 14.440000 1.750000 ;
      RECT 14.470000 0.425000 14.640000 0.595000 ;
      RECT 14.470000 3.475000 14.640000 3.645000 ;
      RECT 14.630000 1.580000 14.800000 1.750000 ;
      RECT 14.830000 0.425000 15.000000 0.595000 ;
      RECT 14.830000 3.475000 15.000000 3.645000 ;
      RECT 15.250000 2.320000 15.420000 2.490000 ;
      RECT 15.670000 3.475000 15.840000 3.645000 ;
      RECT 15.830000 1.580000 16.000000 1.750000 ;
      RECT 16.030000 0.425000 16.200000 0.595000 ;
      RECT 16.030000 3.475000 16.200000 3.645000 ;
      RECT 16.190000 1.580000 16.360000 1.750000 ;
      RECT 16.390000 0.425000 16.560000 0.595000 ;
      RECT 16.390000 3.475000 16.560000 3.645000 ;
      RECT 16.810000 2.320000 16.980000 2.490000 ;
      RECT 17.230000 3.475000 17.400000 3.645000 ;
      RECT 17.390000 1.580000 17.560000 1.750000 ;
      RECT 17.590000 0.425000 17.760000 0.595000 ;
      RECT 17.590000 3.475000 17.760000 3.645000 ;
      RECT 17.750000 1.580000 17.920000 1.750000 ;
      RECT 17.950000 0.425000 18.120000 0.595000 ;
      RECT 17.950000 3.475000 18.120000 3.645000 ;
      RECT 18.370000 2.320000 18.540000 2.490000 ;
      RECT 18.790000 3.475000 18.960000 3.645000 ;
      RECT 18.950000 1.580000 19.120000 1.750000 ;
      RECT 19.150000 0.425000 19.320000 0.595000 ;
      RECT 19.150000 3.475000 19.320000 3.645000 ;
      RECT 19.310000 1.580000 19.480000 1.750000 ;
      RECT 19.510000 0.425000 19.680000 0.595000 ;
      RECT 19.510000 3.475000 19.680000 3.645000 ;
      RECT 19.930000 2.320000 20.100000 2.490000 ;
      RECT 20.430000 3.475000 20.600000 3.645000 ;
      RECT 20.500000 1.580000 20.670000 1.750000 ;
      RECT 20.790000 0.425000 20.960000 0.595000 ;
      RECT 20.790000 3.475000 20.960000 3.645000 ;
      RECT 20.860000 1.580000 21.030000 1.750000 ;
      RECT 21.490000 2.320000 21.660000 2.490000 ;
      RECT 21.910000 3.475000 22.080000 3.645000 ;
      RECT 22.070000 1.580000 22.240000 1.750000 ;
      RECT 22.270000 0.425000 22.440000 0.595000 ;
      RECT 22.270000 3.475000 22.440000 3.645000 ;
      RECT 22.430000 1.580000 22.600000 1.750000 ;
      RECT 22.630000 0.425000 22.800000 0.595000 ;
      RECT 22.630000 3.475000 22.800000 3.645000 ;
      RECT 23.050000 2.320000 23.220000 2.490000 ;
      RECT 23.470000 3.475000 23.640000 3.645000 ;
      RECT 23.630000 1.580000 23.800000 1.750000 ;
      RECT 23.830000 0.425000 24.000000 0.595000 ;
      RECT 23.830000 3.475000 24.000000 3.645000 ;
      RECT 23.990000 1.580000 24.160000 1.750000 ;
      RECT 24.190000 0.425000 24.360000 0.595000 ;
      RECT 24.190000 3.475000 24.360000 3.645000 ;
      RECT 24.610000 2.320000 24.780000 2.490000 ;
      RECT 25.030000 3.475000 25.200000 3.645000 ;
      RECT 25.190000 1.580000 25.360000 1.750000 ;
      RECT 25.390000 0.425000 25.560000 0.595000 ;
      RECT 25.390000 3.475000 25.560000 3.645000 ;
      RECT 25.550000 1.580000 25.720000 1.750000 ;
      RECT 25.750000 0.425000 25.920000 0.595000 ;
      RECT 25.750000 3.475000 25.920000 3.645000 ;
      RECT 26.170000 2.320000 26.340000 2.490000 ;
      RECT 26.590000 3.475000 26.760000 3.645000 ;
      RECT 26.750000 1.580000 26.920000 1.750000 ;
      RECT 26.950000 0.425000 27.120000 0.595000 ;
      RECT 26.950000 3.475000 27.120000 3.645000 ;
      RECT 27.110000 1.580000 27.280000 1.750000 ;
      RECT 27.310000 0.425000 27.480000 0.595000 ;
      RECT 27.310000 3.475000 27.480000 3.645000 ;
      RECT 27.730000 2.320000 27.900000 2.490000 ;
      RECT 28.150000 3.475000 28.320000 3.645000 ;
      RECT 28.310000 1.580000 28.480000 1.750000 ;
      RECT 28.510000 0.425000 28.680000 0.595000 ;
      RECT 28.510000 3.475000 28.680000 3.645000 ;
      RECT 28.670000 1.580000 28.840000 1.750000 ;
      RECT 28.870000 0.425000 29.040000 0.595000 ;
      RECT 28.870000 3.475000 29.040000 3.645000 ;
      RECT 29.290000 2.320000 29.460000 2.490000 ;
      RECT 29.710000 3.475000 29.880000 3.645000 ;
      RECT 29.870000 1.580000 30.040000 1.750000 ;
      RECT 30.070000 0.425000 30.240000 0.595000 ;
      RECT 30.070000 3.475000 30.240000 3.645000 ;
      RECT 30.230000 1.580000 30.400000 1.750000 ;
      RECT 30.430000 0.425000 30.600000 0.595000 ;
      RECT 30.430000 3.475000 30.600000 3.645000 ;
      RECT 30.850000 2.320000 31.020000 2.490000 ;
      RECT 31.270000 3.475000 31.440000 3.645000 ;
      RECT 31.430000 1.580000 31.600000 1.750000 ;
      RECT 31.630000 0.425000 31.800000 0.595000 ;
      RECT 31.630000 3.475000 31.800000 3.645000 ;
      RECT 31.790000 1.580000 31.960000 1.750000 ;
      RECT 31.990000 0.425000 32.160000 0.595000 ;
      RECT 31.990000 3.475000 32.160000 3.645000 ;
      RECT 32.410000 2.320000 32.580000 2.490000 ;
      RECT 32.910000 3.475000 33.080000 3.645000 ;
      RECT 33.270000 0.425000 33.440000 0.595000 ;
      RECT 33.270000 3.475000 33.440000 3.645000 ;
    LAYER met1 ;
      RECT 4.960000 1.550000 32.090000 1.780000 ;
  END
END sky130_fd_sc_hvl__buf_32
MACRO sky130_fd_sc_hvl__sdfsbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__sdfsbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  20.16000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN D
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.975000 1.845000 2.305000 2.355000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.498750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 19.700000 0.495000 20.035000 1.325000 ;
        RECT 19.700000 2.355000 20.035000 3.435000 ;
        RECT 19.805000 1.325000 20.035000 2.355000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.611250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 17.405000 0.495000 17.785000 3.735000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 0.810000 3.690000 2.150000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.840000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.495000 2.955000 1.665000 ;
        RECT 0.605000 1.665000 1.795000 2.165000 ;
        RECT 2.680000 1.095000 2.955000 1.495000 ;
        RECT 2.680000 1.665000 2.955000 1.765000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.840000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.205000 1.210000 12.355000 1.380000 ;
        RECT 12.185000 0.265000 14.170000 0.435000 ;
        RECT 12.185000 0.435000 12.355000 1.210000 ;
        RECT 14.000000 0.435000 14.170000 1.425000 ;
        RECT 14.000000 1.425000 14.845000 1.645000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.380000 1.180000 4.710000 2.150000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 20.160000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 20.160000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 20.160000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 20.160000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 20.490000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 20.160000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 20.160000 0.085000 ;
      RECT  0.000000  3.985000 20.160000 4.155000 ;
      RECT  0.130000  0.495000  0.485000 1.095000 ;
      RECT  0.130000  1.095000  2.300000 1.315000 ;
      RECT  0.130000  1.315000  0.300000 2.535000 ;
      RECT  0.130000  2.535000  2.885000 2.705000 ;
      RECT  0.130000  2.705000  0.460000 3.305000 ;
      RECT  0.640000  2.885000  1.590000 3.705000 ;
      RECT  0.665000  0.365000  1.615000 0.915000 ;
      RECT  2.400000  2.885000  3.235000 3.055000 ;
      RECT  2.400000  3.055000  2.730000 3.305000 ;
      RECT  2.425000  0.495000  2.755000 0.745000 ;
      RECT  2.425000  0.745000  3.305000 0.915000 ;
      RECT  2.635000  2.015000  2.885000 2.535000 ;
      RECT  3.065000  2.455000  4.655000 2.625000 ;
      RECT  3.065000  2.625000  3.235000 2.885000 ;
      RECT  3.135000  0.915000  3.305000 2.455000 ;
      RECT  3.415000  2.805000  4.305000 3.705000 ;
      RECT  3.870000  0.365000  4.760000 0.995000 ;
      RECT  4.485000  2.625000  4.655000 3.635000 ;
      RECT  4.485000  3.635000  5.515000 3.805000 ;
      RECT  4.835000  2.805000  5.165000 3.455000 ;
      RECT  4.940000  0.515000  5.190000 1.700000 ;
      RECT  4.940000  1.700000  6.065000 1.870000 ;
      RECT  4.940000  1.870000  5.165000 2.805000 ;
      RECT  5.345000  2.050000  6.215000 2.220000 ;
      RECT  5.345000  2.220000  5.515000 3.635000 ;
      RECT  5.370000  0.365000  5.960000 1.020000 ;
      RECT  5.695000  2.400000  5.865000 3.705000 ;
      RECT  5.735000  1.200000  6.065000 1.700000 ;
      RECT  6.045000  2.220000  6.215000 3.390000 ;
      RECT  6.045000  3.390000  7.295000 3.560000 ;
      RECT  6.190000  0.265000  8.220000 0.435000 ;
      RECT  6.190000  0.435000  6.565000 1.020000 ;
      RECT  6.395000  1.020000  6.565000 2.290000 ;
      RECT  6.395000  2.290000  6.645000 3.210000 ;
      RECT  6.760000  0.615000  7.010000 1.060000 ;
      RECT  6.840000  1.060000  7.010000 2.740000 ;
      RECT  6.840000  2.740000  7.295000 3.390000 ;
      RECT  7.190000  0.435000  7.360000 2.290000 ;
      RECT  7.190000  2.290000  7.520000 2.560000 ;
      RECT  7.540000  0.640000  7.870000 1.060000 ;
      RECT  7.700000  1.060000  7.870000 1.910000 ;
      RECT  7.700000  1.910000 11.645000 2.080000 ;
      RECT  7.700000  2.080000  7.995000 3.240000 ;
      RECT  8.050000  0.435000  8.220000 1.150000 ;
      RECT  8.050000  1.150000  8.325000 1.560000 ;
      RECT  8.050000  1.560000 12.530000 1.730000 ;
      RECT  8.200000  2.290000  8.530000 2.610000 ;
      RECT  8.200000  2.610000  9.915000 2.780000 ;
      RECT  8.410000  0.365000  9.360000 0.960000 ;
      RECT  8.615000  2.960000  9.565000 3.705000 ;
      RECT  8.910000  1.140000  9.910000 1.380000 ;
      RECT  8.910000  2.260000 10.425000 2.430000 ;
      RECT  9.580000  0.515000  9.910000 1.140000 ;
      RECT  9.745000  2.780000  9.915000 3.170000 ;
      RECT  9.745000  3.170000 10.775000 3.340000 ;
      RECT 10.095000  2.430000 10.425000 2.990000 ;
      RECT 10.545000  0.365000 11.495000 1.030000 ;
      RECT 10.605000  3.000000 12.335000 3.170000 ;
      RECT 10.955000  3.350000 11.905000 3.755000 ;
      RECT 11.315000  2.080000 11.645000 2.555000 ;
      RECT 12.025000  2.125000 13.405000 2.295000 ;
      RECT 12.025000  2.295000 12.335000 3.000000 ;
      RECT 12.200000  1.730000 12.530000 1.875000 ;
      RECT 12.515000  2.525000 15.300000 2.695000 ;
      RECT 12.515000  2.695000 12.845000 3.755000 ;
      RECT 12.655000  0.615000 13.755000 0.785000 ;
      RECT 12.655000  0.785000 12.985000 1.325000 ;
      RECT 13.165000  1.415000 13.405000 2.125000 ;
      RECT 13.500000  2.875000 14.450000 3.705000 ;
      RECT 13.585000  0.785000 13.755000 1.825000 ;
      RECT 13.585000  1.825000 15.545000 1.995000 ;
      RECT 13.585000  1.995000 13.755000 2.525000 ;
      RECT 13.935000  2.175000 16.060000 2.345000 ;
      RECT 14.350000  0.365000 15.300000 1.245000 ;
      RECT 14.970000  2.695000 15.300000 3.175000 ;
      RECT 15.215000  1.425000 15.545000 1.825000 ;
      RECT 15.685000  2.345000 16.060000 2.675000 ;
      RECT 15.730000  0.825000 16.060000 2.175000 ;
      RECT 16.240000  0.365000 17.190000 1.325000 ;
      RECT 16.240000  2.195000 17.190000 3.735000 ;
      RECT 18.025000  0.825000 18.355000 1.505000 ;
      RECT 18.025000  1.505000 19.575000 1.675000 ;
      RECT 18.025000  1.675000 18.355000 3.185000 ;
      RECT 18.535000  0.365000 19.485000 1.325000 ;
      RECT 18.535000  2.355000 19.485000 3.705000 ;
      RECT 19.245000  1.675000 19.575000 2.175000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.985000  0.325000 4.155000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.985000  0.805000 4.155000 ;
      RECT  0.670000  3.505000  0.840000 3.675000 ;
      RECT  0.695000  0.395000  0.865000 0.565000 ;
      RECT  1.030000  3.505000  1.200000 3.675000 ;
      RECT  1.055000  0.395000  1.225000 0.565000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.985000  1.285000 4.155000 ;
      RECT  1.390000  3.505000  1.560000 3.675000 ;
      RECT  1.415000  0.395000  1.585000 0.565000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.985000  1.765000 4.155000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.985000  2.245000 4.155000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.985000  2.725000 4.155000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.985000  3.205000 4.155000 ;
      RECT  3.415000  3.505000  3.585000 3.675000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.985000  3.685000 4.155000 ;
      RECT  3.775000  3.505000  3.945000 3.675000 ;
      RECT  3.870000  0.395000  4.040000 0.565000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.985000  4.165000 4.155000 ;
      RECT  4.135000  3.505000  4.305000 3.675000 ;
      RECT  4.230000  0.395000  4.400000 0.565000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.985000  4.645000 4.155000 ;
      RECT  4.590000  0.395000  4.760000 0.565000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.985000  5.125000 4.155000 ;
      RECT  5.400000  0.395000  5.570000 0.565000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.985000  5.605000 4.155000 ;
      RECT  5.695000  3.505000  5.865000 3.675000 ;
      RECT  5.760000  0.395000  5.930000 0.565000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.985000  6.085000 4.155000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.985000  6.565000 4.155000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.985000  7.045000 4.155000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.985000  7.525000 4.155000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.985000  8.005000 4.155000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.985000  8.485000 4.155000 ;
      RECT  8.440000  0.395000  8.610000 0.565000 ;
      RECT  8.645000  3.505000  8.815000 3.675000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.985000  8.965000 4.155000 ;
      RECT  8.800000  0.395000  8.970000 0.565000 ;
      RECT  9.005000  3.505000  9.175000 3.675000 ;
      RECT  9.160000  0.395000  9.330000 0.565000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.985000  9.445000 4.155000 ;
      RECT  9.365000  3.505000  9.535000 3.675000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.985000  9.925000 4.155000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.985000 10.405000 4.155000 ;
      RECT 10.575000  0.395000 10.745000 0.565000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.985000 10.885000 4.155000 ;
      RECT 10.935000  0.395000 11.105000 0.565000 ;
      RECT 10.985000  3.505000 11.155000 3.675000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.985000 11.365000 4.155000 ;
      RECT 11.295000  0.395000 11.465000 0.565000 ;
      RECT 11.345000  3.505000 11.515000 3.675000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.985000 11.845000 4.155000 ;
      RECT 11.705000  3.505000 11.875000 3.675000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.985000 12.325000 4.155000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.985000 12.805000 4.155000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.985000 13.285000 4.155000 ;
      RECT 13.530000  3.505000 13.700000 3.675000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.985000 13.765000 4.155000 ;
      RECT 13.890000  3.505000 14.060000 3.675000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.985000 14.245000 4.155000 ;
      RECT 14.250000  3.505000 14.420000 3.675000 ;
      RECT 14.380000  0.395000 14.550000 0.565000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.985000 14.725000 4.155000 ;
      RECT 14.740000  0.395000 14.910000 0.565000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.985000 15.205000 4.155000 ;
      RECT 15.100000  0.395000 15.270000 0.565000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.985000 15.685000 4.155000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000  3.985000 16.165000 4.155000 ;
      RECT 16.270000  0.395000 16.440000 0.565000 ;
      RECT 16.270000  3.505000 16.440000 3.675000 ;
      RECT 16.475000 -0.085000 16.645000 0.085000 ;
      RECT 16.475000  3.985000 16.645000 4.155000 ;
      RECT 16.630000  0.395000 16.800000 0.565000 ;
      RECT 16.630000  3.505000 16.800000 3.675000 ;
      RECT 16.955000 -0.085000 17.125000 0.085000 ;
      RECT 16.955000  3.985000 17.125000 4.155000 ;
      RECT 16.990000  0.395000 17.160000 0.565000 ;
      RECT 16.990000  3.505000 17.160000 3.675000 ;
      RECT 17.435000 -0.085000 17.605000 0.085000 ;
      RECT 17.435000  3.985000 17.605000 4.155000 ;
      RECT 17.915000 -0.085000 18.085000 0.085000 ;
      RECT 17.915000  3.985000 18.085000 4.155000 ;
      RECT 18.395000 -0.085000 18.565000 0.085000 ;
      RECT 18.395000  3.985000 18.565000 4.155000 ;
      RECT 18.565000  0.395000 18.735000 0.565000 ;
      RECT 18.565000  3.505000 18.735000 3.675000 ;
      RECT 18.875000 -0.085000 19.045000 0.085000 ;
      RECT 18.875000  3.985000 19.045000 4.155000 ;
      RECT 18.925000  0.395000 19.095000 0.565000 ;
      RECT 18.925000  3.505000 19.095000 3.675000 ;
      RECT 19.285000  0.395000 19.455000 0.565000 ;
      RECT 19.285000  3.505000 19.455000 3.675000 ;
      RECT 19.355000 -0.085000 19.525000 0.085000 ;
      RECT 19.355000  3.985000 19.525000 4.155000 ;
      RECT 19.835000 -0.085000 20.005000 0.085000 ;
      RECT 19.835000  3.985000 20.005000 4.155000 ;
  END
END sky130_fd_sc_hvl__sdfsbp_1
MACRO sky130_fd_sc_hvl__a22oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__a22oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A1
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.505000 2.755000 1.750000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.940000 1.505000 3.715000 1.750000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 1.505000 1.795000 1.750000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.505000 0.835000 1.835000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.630000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.925000 2.175000 1.285000 3.455000 ;
        RECT 1.085000 0.810000 1.955000 0.980000 ;
        RECT 1.085000 0.980000 1.285000 2.175000 ;
        RECT 1.705000 0.495000 1.955000 0.810000 ;
        RECT 1.705000 0.980000 1.955000 1.325000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 3.840000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 3.840000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 3.840000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 3.840000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 4.170000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 3.840000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.985000 3.840000 4.155000 ;
      RECT 0.090000  0.365000 0.680000 1.325000 ;
      RECT 0.145000  2.175000 0.475000 3.635000 ;
      RECT 0.145000  3.635000 1.955000 3.805000 ;
      RECT 1.705000  1.930000 3.595000 2.100000 ;
      RECT 1.705000  2.100000 1.955000 3.635000 ;
      RECT 2.135000  0.365000 3.750000 1.325000 ;
      RECT 2.135000  2.280000 3.085000 3.755000 ;
      RECT 3.265000  2.100000 3.595000 3.755000 ;
    LAYER mcon ;
      RECT 0.120000  0.395000 0.290000 0.565000 ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.480000  0.395000 0.650000 0.565000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.135000  0.395000 2.305000 0.565000 ;
      RECT 2.165000  3.505000 2.335000 3.675000 ;
      RECT 2.495000  0.395000 2.665000 0.565000 ;
      RECT 2.525000  3.505000 2.695000 3.675000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 2.855000  0.395000 3.025000 0.565000 ;
      RECT 2.885000  3.505000 3.055000 3.675000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
      RECT 3.215000  0.395000 3.385000 0.565000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.985000 3.685000 4.155000 ;
      RECT 3.575000  0.395000 3.745000 0.565000 ;
  END
END sky130_fd_sc_hvl__a22oi_1
MACRO sky130_fd_sc_hvl__sdfstp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__sdfstp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  18.72000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN D
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.945000 1.845000 2.275000 2.355000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.478750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 18.260000 0.495000 18.610000 3.395000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.420000 1.175000 3.750000 2.150000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.840000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.565000 1.495000 2.890000 1.665000 ;
        RECT 0.565000 1.665000 0.895000 2.165000 ;
        RECT 2.525000 1.095000 2.890000 1.495000 ;
        RECT 2.525000 1.665000 2.890000 1.780000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.840000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.535000 1.175000 11.635000 1.345000 ;
        RECT 11.465000 0.265000 14.215000 0.435000 ;
        RECT 11.465000 0.435000 11.635000 1.175000 ;
        RECT 14.045000 0.435000 14.215000 0.810000 ;
        RECT 14.045000 0.810000 14.520000 1.760000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.175000 4.525000 2.150000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 18.720000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 18.720000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 18.720000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 18.720000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 19.050000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 18.720000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 18.720000 0.085000 ;
      RECT  0.000000  3.985000 18.720000 4.155000 ;
      RECT  0.110000  0.515000  0.440000 1.095000 ;
      RECT  0.110000  1.095000  2.255000 1.315000 ;
      RECT  0.110000  1.315000  0.280000 2.535000 ;
      RECT  0.110000  2.535000  2.890000 2.705000 ;
      RECT  0.110000  2.705000  0.440000 3.285000 ;
      RECT  0.620000  0.365000  1.570000 0.915000 ;
      RECT  0.620000  2.885000  1.570000 3.705000 ;
      RECT  2.380000  0.495000  2.710000 0.745000 ;
      RECT  2.380000  0.745000  3.240000 0.915000 ;
      RECT  2.380000  2.885000  3.240000 3.055000 ;
      RECT  2.380000  3.055000  2.710000 3.305000 ;
      RECT  2.635000  2.015000  2.890000 2.535000 ;
      RECT  3.070000  0.915000  3.240000 2.455000 ;
      RECT  3.070000  2.455000  4.665000 2.625000 ;
      RECT  3.070000  2.625000  3.240000 2.885000 ;
      RECT  3.420000  0.365000  4.370000 0.995000 ;
      RECT  3.420000  2.805000  4.315000 3.705000 ;
      RECT  4.495000  2.625000  4.665000 3.635000 ;
      RECT  4.495000  3.635000  5.365000 3.805000 ;
      RECT  4.650000  0.515000  5.015000 0.975000 ;
      RECT  4.845000  0.975000  5.015000 1.735000 ;
      RECT  4.845000  1.735000  5.835000 1.905000 ;
      RECT  4.845000  1.905000  5.015000 3.455000 ;
      RECT  5.195000  2.275000  6.075000 2.445000 ;
      RECT  5.195000  2.445000  5.365000 3.635000 ;
      RECT  5.200000  0.365000  5.450000 1.055000 ;
      RECT  5.505000  1.235000  5.835000 1.735000 ;
      RECT  5.545000  2.625000  5.725000 3.705000 ;
      RECT  5.630000  0.265000  7.230000 0.435000 ;
      RECT  5.630000  0.435000  5.800000 1.235000 ;
      RECT  5.905000  2.445000  6.075000 3.635000 ;
      RECT  5.905000  3.635000  7.095000 3.805000 ;
      RECT  5.980000  0.675000  6.310000 1.055000 ;
      RECT  6.140000  1.055000  6.310000 1.425000 ;
      RECT  6.140000  1.425000  6.530000 2.095000 ;
      RECT  6.255000  2.095000  6.530000 3.455000 ;
      RECT  6.550000  0.615000  6.880000 1.025000 ;
      RECT  6.710000  1.025000  6.880000 2.675000 ;
      RECT  6.710000  2.675000  7.095000 3.635000 ;
      RECT  7.060000  0.435000  7.230000 1.605000 ;
      RECT  7.060000  1.605000  7.445000 1.775000 ;
      RECT  7.275000  1.775000  7.445000 3.355000 ;
      RECT  7.275000  3.355000  8.305000 3.525000 ;
      RECT  7.410000  0.525000  7.795000 1.025000 ;
      RECT  7.625000  1.025000  7.795000 1.355000 ;
      RECT  7.625000  1.355000  8.655000 1.525000 ;
      RECT  7.625000  1.525000  7.795000 2.675000 ;
      RECT  7.625000  2.675000  7.955000 3.175000 ;
      RECT  7.975000  1.705000  8.305000 1.875000 ;
      RECT  7.975000  1.875000 12.220000 2.045000 ;
      RECT  8.135000  2.225000  8.410000 2.575000 ;
      RECT  8.135000  2.575000  9.795000 2.745000 ;
      RECT  8.135000  2.745000  8.305000 3.355000 ;
      RECT  8.200000  0.365000  9.150000 0.925000 ;
      RECT  8.485000  1.525000 11.525000 1.695000 ;
      RECT  8.495000  2.925000  9.445000 3.705000 ;
      RECT  8.790000  2.225000 10.305000 2.395000 ;
      RECT  8.835000  1.105000  9.700000 1.275000 ;
      RECT  8.835000  1.275000  9.165000 1.345000 ;
      RECT  9.370000  0.515000  9.700000 1.105000 ;
      RECT  9.520000  1.455000  9.850000 1.525000 ;
      RECT  9.625000  2.745000  9.795000 3.105000 ;
      RECT  9.625000  3.105000 10.655000 3.275000 ;
      RECT  9.975000  2.395000 10.305000 2.925000 ;
      RECT 10.335000  0.365000 11.285000 0.995000 ;
      RECT 10.485000  2.935000 12.180000 3.105000 ;
      RECT 10.835000  3.285000 11.785000 3.755000 ;
      RECT 11.905000  2.225000 12.570000 2.395000 ;
      RECT 11.905000  2.395000 12.180000 2.935000 ;
      RECT 11.970000  1.685000 12.220000 1.875000 ;
      RECT 12.095000  0.615000 13.350000 0.785000 ;
      RECT 12.095000  0.785000 12.265000 1.335000 ;
      RECT 12.095000  1.335000 12.570000 1.505000 ;
      RECT 12.360000  2.675000 12.920000 2.845000 ;
      RECT 12.360000  2.845000 12.690000 3.755000 ;
      RECT 12.400000  1.505000 12.570000 2.225000 ;
      RECT 12.445000  0.965000 12.920000 1.155000 ;
      RECT 12.750000  1.155000 12.920000 1.940000 ;
      RECT 12.750000  1.940000 15.585000 2.110000 ;
      RECT 12.750000  2.110000 12.920000 2.675000 ;
      RECT 13.100000  0.785000 13.350000 1.745000 ;
      RECT 13.265000  2.675000 14.215000 3.705000 ;
      RECT 13.710000  2.290000 14.565000 2.495000 ;
      RECT 14.395000  2.495000 14.565000 3.335000 ;
      RECT 14.395000  3.335000 15.625000 3.505000 ;
      RECT 14.700000  0.365000 15.590000 1.325000 ;
      RECT 14.745000  2.110000 15.585000 2.175000 ;
      RECT 14.745000  2.175000 15.075000 3.155000 ;
      RECT 15.255000  1.505000 15.585000 1.940000 ;
      RECT 15.295000  2.695000 16.020000 2.865000 ;
      RECT 15.295000  2.865000 15.625000 3.335000 ;
      RECT 15.770000  0.825000 16.020000 2.695000 ;
      RECT 15.815000  3.045000 16.405000 3.705000 ;
      RECT 16.585000  0.825000 16.915000 1.505000 ;
      RECT 16.585000  1.505000 18.080000 1.675000 ;
      RECT 16.585000  1.675000 16.915000 2.355000 ;
      RECT 16.585000  2.355000 16.955000 3.145000 ;
      RECT 17.095000  0.365000 18.045000 1.325000 ;
      RECT 17.135000  2.355000 18.080000 3.705000 ;
      RECT 17.750000  1.675000 18.080000 2.175000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.985000  0.325000 4.155000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.985000  0.805000 4.155000 ;
      RECT  0.650000  0.395000  0.820000 0.565000 ;
      RECT  0.650000  3.505000  0.820000 3.675000 ;
      RECT  1.010000  0.395000  1.180000 0.565000 ;
      RECT  1.010000  3.505000  1.180000 3.675000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.985000  1.285000 4.155000 ;
      RECT  1.370000  0.395000  1.540000 0.565000 ;
      RECT  1.370000  3.505000  1.540000 3.675000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.985000  1.765000 4.155000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.985000  2.245000 4.155000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.985000  2.725000 4.155000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.985000  3.205000 4.155000 ;
      RECT  3.420000  3.505000  3.590000 3.675000 ;
      RECT  3.450000  0.395000  3.620000 0.565000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.985000  3.685000 4.155000 ;
      RECT  3.780000  3.505000  3.950000 3.675000 ;
      RECT  3.810000  0.395000  3.980000 0.565000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.985000  4.165000 4.155000 ;
      RECT  4.140000  3.505000  4.310000 3.675000 ;
      RECT  4.170000  0.395000  4.340000 0.565000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.985000  4.645000 4.155000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.985000  5.125000 4.155000 ;
      RECT  5.230000  0.395000  5.400000 0.565000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.985000  5.605000 4.155000 ;
      RECT  5.550000  3.505000  5.720000 3.675000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.985000  6.085000 4.155000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.985000  6.565000 4.155000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.985000  7.045000 4.155000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.985000  7.525000 4.155000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.985000  8.005000 4.155000 ;
      RECT  8.230000  0.395000  8.400000 0.565000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.985000  8.485000 4.155000 ;
      RECT  8.525000  3.505000  8.695000 3.675000 ;
      RECT  8.590000  0.395000  8.760000 0.565000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.985000  8.965000 4.155000 ;
      RECT  8.885000  3.505000  9.055000 3.675000 ;
      RECT  8.950000  0.395000  9.120000 0.565000 ;
      RECT  9.245000  3.505000  9.415000 3.675000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.985000  9.445000 4.155000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.985000  9.925000 4.155000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.985000 10.405000 4.155000 ;
      RECT 10.365000  0.395000 10.535000 0.565000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.985000 10.885000 4.155000 ;
      RECT 10.725000  0.395000 10.895000 0.565000 ;
      RECT 10.865000  3.505000 11.035000 3.675000 ;
      RECT 11.085000  0.395000 11.255000 0.565000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.985000 11.365000 4.155000 ;
      RECT 11.225000  3.505000 11.395000 3.675000 ;
      RECT 11.585000  3.505000 11.755000 3.675000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.985000 11.845000 4.155000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.985000 12.325000 4.155000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.985000 12.805000 4.155000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.985000 13.285000 4.155000 ;
      RECT 13.295000  3.505000 13.465000 3.675000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.985000 13.765000 4.155000 ;
      RECT 13.655000  3.505000 13.825000 3.675000 ;
      RECT 14.015000  3.505000 14.185000 3.675000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.985000 14.245000 4.155000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.985000 14.725000 4.155000 ;
      RECT 14.700000  0.395000 14.870000 0.565000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.985000 15.205000 4.155000 ;
      RECT 15.060000  0.395000 15.230000 0.565000 ;
      RECT 15.420000  0.395000 15.590000 0.565000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.985000 15.685000 4.155000 ;
      RECT 15.845000  3.505000 16.015000 3.675000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000  3.985000 16.165000 4.155000 ;
      RECT 16.205000  3.505000 16.375000 3.675000 ;
      RECT 16.475000 -0.085000 16.645000 0.085000 ;
      RECT 16.475000  3.985000 16.645000 4.155000 ;
      RECT 16.955000 -0.085000 17.125000 0.085000 ;
      RECT 16.955000  3.985000 17.125000 4.155000 ;
      RECT 17.125000  0.395000 17.295000 0.565000 ;
      RECT 17.160000  3.505000 17.330000 3.675000 ;
      RECT 17.435000 -0.085000 17.605000 0.085000 ;
      RECT 17.435000  3.985000 17.605000 4.155000 ;
      RECT 17.485000  0.395000 17.655000 0.565000 ;
      RECT 17.520000  3.505000 17.690000 3.675000 ;
      RECT 17.845000  0.395000 18.015000 0.565000 ;
      RECT 17.880000  3.505000 18.050000 3.675000 ;
      RECT 17.915000 -0.085000 18.085000 0.085000 ;
      RECT 17.915000  3.985000 18.085000 4.155000 ;
      RECT 18.395000 -0.085000 18.565000 0.085000 ;
      RECT 18.395000  3.985000 18.565000 4.155000 ;
  END
END sky130_fd_sc_hvl__sdfstp_1
MACRO sky130_fd_sc_hvl__nor2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__nor2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.400000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.775000 1.315000 2.120000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.495000 1.775000 1.825000 2.120000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.637500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.200000 0.495000 1.530000 1.425000 ;
        RECT 1.200000 1.425000 2.275000 1.595000 ;
        RECT 2.020000 1.595000 2.275000 3.755000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 2.400000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 2.400000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 2.400000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 2.400000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 2.730000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 2.400000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.400000 0.085000 ;
      RECT 0.000000  3.985000 2.400000 4.155000 ;
      RECT 0.090000  0.365000 1.020000 1.325000 ;
      RECT 0.090000  2.300000 1.760000 3.755000 ;
      RECT 1.720000  0.365000 2.310000 1.245000 ;
    LAYER mcon ;
      RECT 0.110000  0.395000 0.280000 0.565000 ;
      RECT 0.120000  3.505000 0.290000 3.675000 ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.470000  0.395000 0.640000 0.565000 ;
      RECT 0.480000  3.505000 0.650000 3.675000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.830000  0.395000 1.000000 0.565000 ;
      RECT 0.840000  3.505000 1.010000 3.675000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.200000  3.505000 1.370000 3.675000 ;
      RECT 1.560000  3.505000 1.730000 3.675000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.750000  0.395000 1.920000 0.565000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.110000  0.395000 2.280000 0.565000 ;
  END
END sky130_fd_sc_hvl__nor2_1
MACRO sky130_fd_sc_hvl__probe_p_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__probe_p_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.600000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  3.375000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.635000 1.580000 2.245000 1.815000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  2.520000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT 3.290000 1.235000 6.310000 2.835000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 9.600000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 9.600000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 9.600000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 9.600000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 9.930000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 9.600000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.600000 0.085000 ;
      RECT 0.000000  3.985000 9.600000 4.155000 ;
      RECT 0.245000  0.805000 0.455000 1.475000 ;
      RECT 0.245000  1.475000 0.435000 2.095000 ;
      RECT 0.245000  2.095000 2.595000 2.265000 ;
      RECT 0.245000  2.265000 0.435000 3.545000 ;
      RECT 0.615000  2.445000 1.865000 3.625000 ;
      RECT 0.615000  3.625000 9.505000 3.795000 ;
      RECT 0.675000  0.380000 9.505000 0.550000 ;
      RECT 0.675000  0.550000 1.925000 1.385000 ;
      RECT 2.045000  2.265000 2.595000 3.445000 ;
      RECT 2.105000  0.730000 2.315000 1.230000 ;
      RECT 2.105000  1.230000 2.595000 1.400000 ;
      RECT 2.425000  1.400000 2.595000 1.625000 ;
      RECT 2.425000  1.625000 3.380000 1.955000 ;
      RECT 2.425000  1.955000 2.595000 2.095000 ;
      RECT 2.605000  0.550000 3.495000 0.760000 ;
      RECT 2.765000  0.760000 3.495000 1.445000 ;
      RECT 2.765000  2.385000 3.435000 3.625000 ;
      RECT 3.605000  2.035000 8.965000 2.205000 ;
      RECT 3.605000  2.205000 3.935000 3.445000 ;
      RECT 3.665000  0.805000 3.875000 1.625000 ;
      RECT 3.665000  1.625000 8.555000 1.795000 ;
      RECT 4.045000  0.550000 5.055000 1.445000 ;
      RECT 4.105000  2.385000 4.995000 3.625000 ;
      RECT 5.165000  2.205000 5.495000 3.445000 ;
      RECT 5.225000  0.805000 5.435000 1.625000 ;
      RECT 5.605000  0.550000 6.615000 1.445000 ;
      RECT 5.665000  2.385000 6.555000 3.625000 ;
      RECT 6.725000  2.205000 7.055000 3.445000 ;
      RECT 6.785000  0.805000 6.995000 1.625000 ;
      RECT 7.165000  0.550000 8.175000 1.445000 ;
      RECT 7.225000  2.385000 8.115000 3.625000 ;
      RECT 8.285000  2.205000 8.965000 3.230000 ;
      RECT 8.285000  3.230000 8.735000 3.445000 ;
      RECT 8.345000  0.805000 8.965000 0.975000 ;
      RECT 8.345000  0.975000 8.555000 1.625000 ;
      RECT 8.735000  0.975000 8.965000 2.035000 ;
      RECT 8.905000  3.475000 9.505000 3.625000 ;
      RECT 8.975000  0.550000 9.505000 0.600000 ;
      RECT 9.135000  0.600000 9.505000 1.445000 ;
      RECT 9.135000  2.385000 9.505000 3.475000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.615000  3.475000 0.785000 3.645000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.975000  3.475000 1.145000 3.645000 ;
      RECT 1.035000  0.380000 1.205000 0.550000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.335000  3.475000 1.505000 3.645000 ;
      RECT 1.395000  0.380000 1.565000 0.550000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.695000  3.475000 1.865000 3.645000 ;
      RECT 1.755000  0.380000 1.925000 0.550000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 2.605000  0.380000 2.775000 0.550000 ;
      RECT 2.770000  3.475000 2.940000 3.645000 ;
      RECT 2.965000  0.380000 3.135000 0.550000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
      RECT 3.130000  3.475000 3.300000 3.645000 ;
      RECT 3.325000  0.380000 3.495000 0.550000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.985000 3.685000 4.155000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.985000 4.165000 4.155000 ;
      RECT 4.070000  0.380000 4.240000 0.550000 ;
      RECT 4.105000  3.475000 4.275000 3.645000 ;
      RECT 4.430000  0.380000 4.600000 0.550000 ;
      RECT 4.465000  3.475000 4.635000 3.645000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.985000 4.645000 4.155000 ;
      RECT 4.790000  0.380000 4.960000 0.550000 ;
      RECT 4.825000  3.475000 4.995000 3.645000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.985000 5.125000 4.155000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.985000 5.605000 4.155000 ;
      RECT 5.665000  3.475000 5.835000 3.645000 ;
      RECT 5.670000  0.380000 5.840000 0.550000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.985000 6.085000 4.155000 ;
      RECT 6.025000  3.475000 6.195000 3.645000 ;
      RECT 6.030000  0.380000 6.200000 0.550000 ;
      RECT 6.385000  3.475000 6.555000 3.645000 ;
      RECT 6.390000  0.380000 6.560000 0.550000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.985000 6.565000 4.155000 ;
      RECT 6.725000  2.035000 6.895000 2.205000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.985000 7.045000 4.155000 ;
      RECT 7.085000  2.035000 7.255000 2.205000 ;
      RECT 7.230000  3.475000 7.400000 3.645000 ;
      RECT 7.235000  0.380000 7.405000 0.550000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.985000 7.525000 4.155000 ;
      RECT 7.595000  0.380000 7.765000 0.550000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.985000 8.005000 4.155000 ;
      RECT 7.945000  3.475000 8.115000 3.645000 ;
      RECT 7.955000  0.380000 8.125000 0.550000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.985000 8.485000 4.155000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.985000 8.965000 4.155000 ;
      RECT 8.975000  0.380000 9.145000 0.550000 ;
      RECT 9.265000  3.475000 9.435000 3.645000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.985000 9.445000 4.155000 ;
      RECT 9.335000  0.380000 9.505000 0.550000 ;
    LAYER met1 ;
      RECT 5.505000 1.975000 6.145000 2.005000 ;
      RECT 5.505000 2.005000 7.315000 2.235000 ;
    LAYER met2 ;
      RECT 5.485000 1.865000 6.165000 2.235000 ;
    LAYER met3 ;
      RECT 5.435000 1.885000 6.215000 2.215000 ;
    LAYER met4 ;
      RECT 3.410000 1.355000 6.190000 2.535000 ;
    LAYER via ;
      RECT 5.535000 1.975000 5.795000 2.235000 ;
      RECT 5.855000 1.975000 6.115000 2.235000 ;
    LAYER via2 ;
      RECT 5.485000 1.910000 5.765000 2.190000 ;
      RECT 5.885000 1.910000 6.165000 2.190000 ;
    LAYER via3 ;
      RECT 5.465000 1.890000 5.785000 2.210000 ;
      RECT 5.865000 1.890000 6.185000 2.210000 ;
    LAYER via4 ;
      RECT 5.010000 1.355000 6.190000 2.535000 ;
  END
END sky130_fd_sc_hvl__probe_p_8
MACRO sky130_fd_sc_hvl__a21o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__a21o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A1
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.805000 1.505000 3.715000 1.835000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.895000 1.505000 4.195000 1.835000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.505000 2.275000 1.750000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.611250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 0.495000 0.460000 1.325000 ;
        RECT 0.110000 1.325000 0.360000 3.735000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 4.320000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 4.320000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 4.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 4.320000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 4.650000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 4.320000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.985000 4.320000 4.155000 ;
      RECT 0.540000  2.280000 1.440000 3.755000 ;
      RECT 0.565000  1.725000 0.895000 1.930000 ;
      RECT 0.565000  1.930000 2.625000 2.100000 ;
      RECT 0.640000  0.365000 2.250000 1.325000 ;
      RECT 1.620000  2.100000 1.870000 3.755000 ;
      RECT 2.320000  2.280000 4.210000 2.450000 ;
      RECT 2.320000  2.450000 2.650000 3.755000 ;
      RECT 2.430000  0.495000 2.680000 1.325000 ;
      RECT 2.455000  1.325000 2.625000 1.930000 ;
      RECT 2.830000  2.630000 3.780000 3.755000 ;
      RECT 2.860000  0.365000 4.170000 1.325000 ;
      RECT 3.960000  2.195000 4.210000 2.280000 ;
      RECT 3.960000  2.450000 4.210000 3.735000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.545000  3.505000 0.715000 3.675000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.640000  0.395000 0.810000 0.565000 ;
      RECT 0.905000  3.505000 1.075000 3.675000 ;
      RECT 1.000000  0.395000 1.170000 0.565000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.265000  3.505000 1.435000 3.675000 ;
      RECT 1.360000  0.395000 1.530000 0.565000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.720000  0.395000 1.890000 0.565000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.080000  0.395000 2.250000 0.565000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 2.860000  3.505000 3.030000 3.675000 ;
      RECT 2.890000  0.395000 3.060000 0.565000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
      RECT 3.220000  3.505000 3.390000 3.675000 ;
      RECT 3.250000  0.395000 3.420000 0.565000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.985000 3.685000 4.155000 ;
      RECT 3.580000  3.505000 3.750000 3.675000 ;
      RECT 3.610000  0.395000 3.780000 0.565000 ;
      RECT 3.970000  0.395000 4.140000 0.565000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.985000 4.165000 4.155000 ;
  END
END sky130_fd_sc_hvl__a21o_1
MACRO sky130_fd_sc_hvl__sdfrtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__sdfrtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  19.20000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN D
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.910000 2.660000 3.205000 3.260000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.626250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 18.820000 0.515000 19.075000 3.755000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  4.415000 2.290000  4.705000 2.335000 ;
        RECT  4.415000 2.335000 14.305000 2.475000 ;
        RECT  4.415000 2.475000  4.705000 2.520000 ;
        RECT  8.255000 2.290000  8.545000 2.335000 ;
        RECT  8.255000 2.475000  8.545000 2.520000 ;
        RECT 14.015000 2.290000 14.305000 2.335000 ;
        RECT 14.015000 2.475000 14.305000 2.520000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.180000 1.115000 1.510000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.840000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.995000 1.445000 2.245000 1.835000 ;
        RECT 1.995000 1.835000 3.175000 2.005000 ;
        RECT 1.995000 2.005000 2.380000 2.575000 ;
        RECT 3.005000 1.550000 5.635000 1.835000 ;
        RECT 4.880000 1.835000 5.635000 2.525000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 15.485000 1.955000 16.140000 2.495000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 19.200000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 19.200000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 19.200000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 19.200000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 19.530000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 19.200000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 19.200000 0.085000 ;
      RECT  0.000000  3.985000 19.200000 4.155000 ;
      RECT  0.305000  1.690000  1.465000 1.860000 ;
      RECT  0.305000  1.860000  0.475000 3.105000 ;
      RECT  0.305000  3.105000  2.730000 3.275000 ;
      RECT  0.305000  3.275000  0.635000 3.705000 ;
      RECT  0.665000  0.265000  3.975000 0.435000 ;
      RECT  0.665000  0.435000  0.995000 0.995000 ;
      RECT  0.730000  2.255000  1.060000 2.755000 ;
      RECT  0.730000  2.755000  2.730000 2.925000 ;
      RECT  1.295000  0.615000  2.485000 0.915000 ;
      RECT  1.295000  0.915000  1.465000 1.690000 ;
      RECT  1.420000  3.455000  2.370000 3.705000 ;
      RECT  1.645000  1.095000  2.810000 1.175000 ;
      RECT  1.645000  1.175000  5.535000 1.265000 ;
      RECT  1.645000  1.265000  1.815000 2.755000 ;
      RECT  2.480000  1.265000  5.535000 1.345000 ;
      RECT  2.480000  1.345000  2.810000 1.655000 ;
      RECT  2.560000  2.310000  3.555000 2.480000 ;
      RECT  2.560000  2.480000  2.730000 2.755000 ;
      RECT  2.560000  3.275000  2.730000 3.535000 ;
      RECT  2.560000  3.535000  3.555000 3.705000 ;
      RECT  3.385000  2.480000  3.555000 2.705000 ;
      RECT  3.385000  2.705000  5.485000 2.875000 ;
      RECT  3.385000  3.055000  4.975000 3.225000 ;
      RECT  3.385000  3.225000  3.555000 3.535000 ;
      RECT  3.645000  0.435000  3.975000 0.995000 ;
      RECT  3.735000  3.405000  4.625000 3.705000 ;
      RECT  3.965000  2.015000  4.300000 2.290000 ;
      RECT  3.965000  2.290000  4.675000 2.525000 ;
      RECT  4.155000  0.365000  5.105000 0.995000 ;
      RECT  4.805000  3.225000  4.975000 3.635000 ;
      RECT  4.805000  3.635000  6.005000 3.805000 ;
      RECT  5.155000  2.875000  5.485000 3.455000 ;
      RECT  5.285000  0.515000  5.535000 1.175000 ;
      RECT  5.755000  0.515000  6.005000 1.005000 ;
      RECT  5.755000  3.165000  6.005000 3.635000 ;
      RECT  5.835000  1.005000  6.005000 3.165000 ;
      RECT  6.185000  0.265000  7.255000 0.435000 ;
      RECT  6.185000  0.435000  6.355000 3.635000 ;
      RECT  6.185000  3.635000  7.215000 3.805000 ;
      RECT  6.535000  0.615000  6.865000 0.995000 ;
      RECT  6.535000  0.995000  6.705000 2.715000 ;
      RECT  6.535000  2.715000  9.215000 2.885000 ;
      RECT  6.535000  2.885000  6.865000 3.455000 ;
      RECT  6.950000  1.915000  7.605000 2.085000 ;
      RECT  6.950000  2.085000  7.280000 2.535000 ;
      RECT  7.045000  0.435000  7.255000 1.175000 ;
      RECT  7.045000  1.175000  9.635000 1.345000 ;
      RECT  7.045000  1.345000  7.255000 1.735000 ;
      RECT  7.045000  3.065000  8.705000 3.235000 ;
      RECT  7.045000  3.235000  7.215000 3.635000 ;
      RECT  7.405000  3.415000  8.355000 3.705000 ;
      RECT  7.435000  1.525000 10.780000 1.695000 ;
      RECT  7.435000  1.695000  7.605000 1.915000 ;
      RECT  7.785000  1.875000 11.130000 2.045000 ;
      RECT  7.785000  2.045000  8.115000 2.535000 ;
      RECT  8.115000  0.365000  9.065000 0.995000 ;
      RECT  8.295000  2.225000  8.760000 2.535000 ;
      RECT  8.535000  3.235000  8.705000 3.635000 ;
      RECT  8.535000  3.635000  9.785000 3.805000 ;
      RECT  8.885000  2.885000  9.215000 3.455000 ;
      RECT  9.045000  2.225000 10.780000 2.395000 ;
      RECT  9.045000  2.395000  9.215000 2.715000 ;
      RECT  9.305000  0.885000  9.635000 1.175000 ;
      RECT  9.455000  2.695000  9.785000 3.135000 ;
      RECT  9.455000  3.135000 12.810000 3.305000 ;
      RECT  9.455000  3.305000  9.785000 3.635000 ;
      RECT  9.840000  0.365000 10.430000 1.345000 ;
      RECT  9.965000  3.485000 10.915000 3.735000 ;
      RECT 10.490000  2.395000 10.780000 2.555000 ;
      RECT 10.610000  0.265000 12.455000 0.435000 ;
      RECT 10.610000  0.435000 10.780000 1.525000 ;
      RECT 10.960000  0.615000 11.325000 1.285000 ;
      RECT 10.960000  1.285000 11.130000 1.875000 ;
      RECT 10.960000  2.045000 11.130000 2.675000 ;
      RECT 10.960000  2.675000 11.440000 2.955000 ;
      RECT 11.310000  1.465000 11.480000 2.285000 ;
      RECT 11.310000  2.285000 11.790000 2.455000 ;
      RECT 11.620000  2.455000 11.790000 3.135000 ;
      RECT 11.660000  0.615000 12.105000 1.365000 ;
      RECT 11.660000  1.365000 11.830000 1.935000 ;
      RECT 11.660000  1.935000 13.200000 2.105000 ;
      RECT 11.970000  2.105000 12.300000 2.955000 ;
      RECT 12.010000  1.545000 14.395000 1.715000 ;
      RECT 12.010000  1.715000 13.020000 1.755000 ;
      RECT 12.285000  0.435000 12.455000 1.545000 ;
      RECT 12.480000  2.285000 12.810000 3.135000 ;
      RECT 13.015000  3.370000 13.965000 3.705000 ;
      RECT 13.030000  2.105000 13.200000 3.020000 ;
      RECT 13.030000  3.020000 14.315000 3.190000 ;
      RECT 13.085000  0.365000 14.035000 1.365000 ;
      RECT 13.380000  1.895000 13.710000 2.670000 ;
      RECT 13.380000  2.670000 14.745000 2.840000 ;
      RECT 14.040000  1.895000 14.370000 2.490000 ;
      RECT 14.145000  3.190000 14.315000 3.355000 ;
      RECT 14.145000  3.355000 15.095000 3.525000 ;
      RECT 14.225000  0.535000 16.085000 0.705000 ;
      RECT 14.225000  0.705000 14.395000 1.545000 ;
      RECT 14.495000  2.840000 14.745000 3.175000 ;
      RECT 14.575000  1.175000 15.535000 1.345000 ;
      RECT 14.575000  1.345000 14.745000 2.670000 ;
      RECT 14.925000  1.605000 16.850000 1.775000 ;
      RECT 14.925000  1.775000 15.255000 2.275000 ;
      RECT 14.925000  2.275000 15.095000 3.355000 ;
      RECT 15.205000  0.885000 15.535000 1.175000 ;
      RECT 15.275000  2.675000 16.165000 3.705000 ;
      RECT 15.755000  0.705000 16.085000 1.255000 ;
      RECT 15.755000  1.255000 17.200000 1.425000 ;
      RECT 16.275000  0.365000 16.865000 0.995000 ;
      RECT 16.345000  1.955000 17.200000 2.125000 ;
      RECT 16.345000  2.125000 16.595000 3.505000 ;
      RECT 17.030000  1.425000 17.200000 1.955000 ;
      RECT 17.065000  2.305000 17.550000 3.005000 ;
      RECT 17.105000  0.825000 17.550000 1.075000 ;
      RECT 17.380000  1.075000 17.550000 1.485000 ;
      RECT 17.380000  1.485000 18.615000 1.815000 ;
      RECT 17.380000  1.815000 17.550000 2.305000 ;
      RECT 17.730000  0.365000 18.640000 1.305000 ;
      RECT 17.730000  2.175000 18.640000 3.755000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.985000  0.325000 4.155000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.985000  0.805000 4.155000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.985000  1.285000 4.155000 ;
      RECT  1.450000  3.505000  1.620000 3.675000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.985000  1.765000 4.155000 ;
      RECT  1.810000  3.505000  1.980000 3.675000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.985000  2.245000 4.155000 ;
      RECT  2.170000  3.505000  2.340000 3.675000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.985000  2.725000 4.155000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.985000  3.205000 4.155000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.985000  3.685000 4.155000 ;
      RECT  3.735000  3.505000  3.905000 3.675000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.985000  4.165000 4.155000 ;
      RECT  4.095000  3.505000  4.265000 3.675000 ;
      RECT  4.185000  0.395000  4.355000 0.565000 ;
      RECT  4.455000  3.505000  4.625000 3.675000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  2.320000  4.645000 2.490000 ;
      RECT  4.475000  3.985000  4.645000 4.155000 ;
      RECT  4.545000  0.395000  4.715000 0.565000 ;
      RECT  4.905000  0.395000  5.075000 0.565000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.985000  5.125000 4.155000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.985000  5.605000 4.155000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.985000  6.085000 4.155000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.985000  6.565000 4.155000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.985000  7.045000 4.155000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.985000  7.525000 4.155000 ;
      RECT  7.435000  3.505000  7.605000 3.675000 ;
      RECT  7.795000  3.505000  7.965000 3.675000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.985000  8.005000 4.155000 ;
      RECT  8.145000  0.395000  8.315000 0.565000 ;
      RECT  8.155000  3.505000  8.325000 3.675000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  2.320000  8.485000 2.490000 ;
      RECT  8.315000  3.985000  8.485000 4.155000 ;
      RECT  8.505000  0.395000  8.675000 0.565000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.985000  8.965000 4.155000 ;
      RECT  8.865000  0.395000  9.035000 0.565000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.985000  9.445000 4.155000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.985000  9.925000 4.155000 ;
      RECT  9.870000  0.395000 10.040000 0.565000 ;
      RECT  9.995000  3.515000 10.165000 3.685000 ;
      RECT 10.230000  0.395000 10.400000 0.565000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.985000 10.405000 4.155000 ;
      RECT 10.355000  3.515000 10.525000 3.685000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.515000 10.885000 3.685000 ;
      RECT 10.715000  3.985000 10.885000 4.155000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.985000 11.365000 4.155000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.985000 11.845000 4.155000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.985000 12.325000 4.155000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.985000 12.805000 4.155000 ;
      RECT 13.045000  3.505000 13.215000 3.675000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  0.395000 13.285000 0.565000 ;
      RECT 13.115000  3.985000 13.285000 4.155000 ;
      RECT 13.405000  3.505000 13.575000 3.675000 ;
      RECT 13.475000  0.395000 13.645000 0.565000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.985000 13.765000 4.155000 ;
      RECT 13.765000  3.505000 13.935000 3.675000 ;
      RECT 13.835000  0.395000 14.005000 0.565000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  2.320000 14.245000 2.490000 ;
      RECT 14.075000  3.985000 14.245000 4.155000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.985000 14.725000 4.155000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.985000 15.205000 4.155000 ;
      RECT 15.275000  3.505000 15.445000 3.675000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.985000 15.685000 4.155000 ;
      RECT 15.635000  3.505000 15.805000 3.675000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000  3.505000 16.165000 3.675000 ;
      RECT 15.995000  3.985000 16.165000 4.155000 ;
      RECT 16.305000  0.395000 16.475000 0.565000 ;
      RECT 16.475000 -0.085000 16.645000 0.085000 ;
      RECT 16.475000  3.985000 16.645000 4.155000 ;
      RECT 16.665000  0.395000 16.835000 0.565000 ;
      RECT 16.955000 -0.085000 17.125000 0.085000 ;
      RECT 16.955000  3.985000 17.125000 4.155000 ;
      RECT 17.435000 -0.085000 17.605000 0.085000 ;
      RECT 17.435000  3.985000 17.605000 4.155000 ;
      RECT 17.740000  0.395000 17.910000 0.565000 ;
      RECT 17.740000  3.505000 17.910000 3.675000 ;
      RECT 17.915000 -0.085000 18.085000 0.085000 ;
      RECT 17.915000  3.985000 18.085000 4.155000 ;
      RECT 18.100000  0.395000 18.270000 0.565000 ;
      RECT 18.100000  3.505000 18.270000 3.675000 ;
      RECT 18.395000 -0.085000 18.565000 0.085000 ;
      RECT 18.395000  3.985000 18.565000 4.155000 ;
      RECT 18.460000  0.395000 18.630000 0.565000 ;
      RECT 18.460000  3.505000 18.630000 3.675000 ;
      RECT 18.875000 -0.085000 19.045000 0.085000 ;
      RECT 18.875000  3.985000 19.045000 4.155000 ;
  END
END sky130_fd_sc_hvl__sdfrtp_1
MACRO sky130_fd_sc_hvl__xnor2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__xnor2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  2.250000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.580000 2.060000 1.750000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  2.250000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.575000 1.725000 0.905000 1.930000 ;
        RECT 0.575000 1.930000 3.255000 2.100000 ;
        RECT 1.565000 2.100000 3.255000 2.120000 ;
        RECT 2.925000 1.805000 3.255000 1.930000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  1.481250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.025000 1.905000 5.155000 2.075000 ;
        RECT 4.025000 2.075000 4.275000 3.755000 ;
        RECT 4.445000 1.545000 5.155000 1.905000 ;
        RECT 4.750000 0.535000 5.155000 1.545000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 5.280000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 5.280000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 5.280000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 5.280000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 5.610000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 5.280000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.280000 0.085000 ;
      RECT 0.000000  3.985000 5.280000 4.155000 ;
      RECT 0.090000  2.630000 0.985000 3.755000 ;
      RECT 0.110000  0.495000 0.440000 1.230000 ;
      RECT 0.110000  1.230000 2.410000 1.400000 ;
      RECT 0.110000  1.400000 0.360000 2.280000 ;
      RECT 0.110000  2.280000 1.335000 2.450000 ;
      RECT 0.610000  0.365000 2.410000 1.050000 ;
      RECT 1.165000  2.450000 1.335000 3.755000 ;
      RECT 1.515000  2.300000 3.845000 3.755000 ;
      RECT 2.240000  1.400000 2.410000 1.455000 ;
      RECT 2.240000  1.455000 3.980000 1.625000 ;
      RECT 2.590000  0.495000 2.920000 1.105000 ;
      RECT 2.590000  1.105000 4.300000 1.285000 ;
      RECT 3.100000  0.365000 3.630000 0.925000 ;
      RECT 3.650000  1.625000 3.980000 1.725000 ;
      RECT 3.970000  0.535000 4.300000 1.105000 ;
      RECT 4.465000  2.255000 5.055000 3.755000 ;
    LAYER mcon ;
      RECT 0.095000  3.505000 0.265000 3.675000 ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.455000  3.505000 0.625000 3.675000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.800000  0.395000 0.970000 0.565000 ;
      RECT 0.815000  3.505000 0.985000 3.675000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.160000  0.395000 1.330000 0.565000 ;
      RECT 1.515000  3.505000 1.685000 3.675000 ;
      RECT 1.520000  0.395000 1.690000 0.565000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.875000  3.505000 2.045000 3.675000 ;
      RECT 1.880000  0.395000 2.050000 0.565000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.235000  3.505000 2.405000 3.675000 ;
      RECT 2.240000  0.395000 2.410000 0.565000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 2.595000  3.505000 2.765000 3.675000 ;
      RECT 2.955000  3.505000 3.125000 3.675000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
      RECT 3.100000  0.395000 3.270000 0.565000 ;
      RECT 3.315000  3.505000 3.485000 3.675000 ;
      RECT 3.460000  0.395000 3.630000 0.565000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.985000 3.685000 4.155000 ;
      RECT 3.675000  3.505000 3.845000 3.675000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.985000 4.165000 4.155000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.985000 4.645000 4.155000 ;
      RECT 4.495000  3.505000 4.665000 3.675000 ;
      RECT 4.855000  3.505000 5.025000 3.675000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.985000 5.125000 4.155000 ;
  END
END sky130_fd_sc_hvl__xnor2_1
MACRO sky130_fd_sc_hvl__probec_p_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__probec_p_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.600000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  3.375000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.635000 1.580000 2.245000 1.815000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  2.520000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.410000 1.445000 3.590000 2.625000 ;
        RECT 5.010000 1.445000 6.190000 2.625000 ;
    END
    PORT
      LAYER met5 ;
        RECT 2.290000  1.235000 6.310000 2.835000 ;
        RECT 4.710000 -0.365000 6.310000 1.235000 ;
        RECT 4.710000  2.835000 6.310000 4.435000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 7.910000 -0.365000 10.410000 1.235000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 9.600000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 9.600000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 9.600000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 9.930000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 7.910000 2.835000 10.410000 4.435000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.600000 0.085000 ;
      RECT 0.000000  3.985000 9.600000 4.155000 ;
      RECT 0.245000  0.805000 0.455000 1.475000 ;
      RECT 0.245000  1.475000 0.435000 2.095000 ;
      RECT 0.245000  2.095000 2.595000 2.265000 ;
      RECT 0.245000  2.265000 0.435000 3.545000 ;
      RECT 0.615000  2.445000 1.865000 3.625000 ;
      RECT 0.615000  3.625000 9.505000 3.795000 ;
      RECT 0.675000  0.380000 9.505000 0.550000 ;
      RECT 0.675000  0.550000 1.925000 1.385000 ;
      RECT 2.045000  2.265000 2.595000 3.445000 ;
      RECT 2.105000  0.730000 2.315000 1.230000 ;
      RECT 2.105000  1.230000 2.595000 1.400000 ;
      RECT 2.425000  1.400000 2.595000 1.625000 ;
      RECT 2.425000  1.625000 3.380000 1.955000 ;
      RECT 2.425000  1.955000 2.595000 2.095000 ;
      RECT 2.605000  0.550000 3.495000 0.760000 ;
      RECT 2.765000  0.760000 3.495000 1.445000 ;
      RECT 2.765000  2.385000 3.435000 3.625000 ;
      RECT 3.605000  1.955000 8.965000 2.205000 ;
      RECT 3.605000  2.205000 3.935000 3.445000 ;
      RECT 3.665000  0.805000 3.875000 1.625000 ;
      RECT 3.665000  1.625000 8.965000 1.955000 ;
      RECT 4.045000  0.550000 5.055000 1.445000 ;
      RECT 4.105000  2.385000 4.995000 3.625000 ;
      RECT 5.165000  2.205000 5.495000 3.445000 ;
      RECT 5.225000  0.805000 5.435000 1.625000 ;
      RECT 5.605000  0.550000 6.615000 1.445000 ;
      RECT 5.665000  2.385000 6.555000 3.625000 ;
      RECT 6.725000  2.205000 7.055000 3.445000 ;
      RECT 6.785000  0.805000 6.995000 1.625000 ;
      RECT 7.165000  0.550000 8.175000 1.445000 ;
      RECT 7.225000  2.385000 8.115000 3.625000 ;
      RECT 8.285000  2.205000 8.965000 3.230000 ;
      RECT 8.285000  3.230000 8.735000 3.445000 ;
      RECT 8.345000  0.805000 8.965000 1.625000 ;
      RECT 8.905000  3.475000 9.505000 3.625000 ;
      RECT 8.975000  0.550000 9.505000 0.600000 ;
      RECT 9.135000  0.600000 9.505000 1.445000 ;
      RECT 9.135000  2.385000 9.505000 3.475000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.615000  3.475000 0.785000 3.645000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.975000  3.475000 1.145000 3.645000 ;
      RECT 1.035000  0.380000 1.205000 0.550000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.335000  3.475000 1.505000 3.645000 ;
      RECT 1.395000  0.380000 1.565000 0.550000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.695000  3.475000 1.865000 3.645000 ;
      RECT 1.755000  0.380000 1.925000 0.550000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 2.605000  0.380000 2.775000 0.550000 ;
      RECT 2.770000  3.475000 2.940000 3.645000 ;
      RECT 2.965000  0.380000 3.135000 0.550000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
      RECT 3.130000  3.475000 3.300000 3.645000 ;
      RECT 3.325000  0.380000 3.495000 0.550000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.985000 3.685000 4.155000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.985000 4.165000 4.155000 ;
      RECT 4.070000  0.380000 4.240000 0.550000 ;
      RECT 4.105000  3.475000 4.275000 3.645000 ;
      RECT 4.430000  0.380000 4.600000 0.550000 ;
      RECT 4.465000  3.475000 4.635000 3.645000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.985000 4.645000 4.155000 ;
      RECT 4.790000  0.380000 4.960000 0.550000 ;
      RECT 4.825000  3.475000 4.995000 3.645000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.985000 5.125000 4.155000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.985000 5.605000 4.155000 ;
      RECT 5.620000  1.950000 5.790000 2.120000 ;
      RECT 5.665000  3.475000 5.835000 3.645000 ;
      RECT 5.670000  0.380000 5.840000 0.550000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.985000 6.085000 4.155000 ;
      RECT 5.980000  1.950000 6.150000 2.120000 ;
      RECT 6.025000  3.475000 6.195000 3.645000 ;
      RECT 6.030000  0.380000 6.200000 0.550000 ;
      RECT 6.385000  3.475000 6.555000 3.645000 ;
      RECT 6.390000  0.380000 6.560000 0.550000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.985000 6.565000 4.155000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.985000 7.045000 4.155000 ;
      RECT 7.230000  3.475000 7.400000 3.645000 ;
      RECT 7.235000  0.380000 7.405000 0.550000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.985000 7.525000 4.155000 ;
      RECT 7.595000  0.380000 7.765000 0.550000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.985000 8.005000 4.155000 ;
      RECT 7.945000  3.475000 8.115000 3.645000 ;
      RECT 7.955000  0.380000 8.125000 0.550000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.985000 8.485000 4.155000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.985000 8.965000 4.155000 ;
      RECT 8.975000  0.380000 9.145000 0.550000 ;
      RECT 9.265000  3.475000 9.435000 3.645000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.985000 9.445000 4.155000 ;
      RECT 9.335000  0.380000 9.505000 0.550000 ;
    LAYER met1 ;
      RECT 0.000000 0.255000 9.600000 0.305000 ;
      RECT 0.000000 0.305000 9.920000 0.565000 ;
      RECT 0.000000 0.565000 9.600000 0.625000 ;
      RECT 0.000000 3.445000 9.600000 3.505000 ;
      RECT 0.000000 3.505000 9.920000 3.765000 ;
      RECT 0.000000 3.765000 9.600000 3.815000 ;
      RECT 5.560000 1.905000 6.210000 2.165000 ;
    LAYER met2 ;
      RECT 5.440000 1.895000 6.210000 2.175000 ;
      RECT 9.215000 0.285000 9.985000 0.565000 ;
      RECT 9.215000 3.505000 9.985000 3.785000 ;
    LAYER met3 ;
      RECT 2.835000 1.875000 3.615000 2.195000 ;
      RECT 5.435000 1.870000 6.215000 2.200000 ;
      RECT 9.210000 0.260000 9.990000 0.590000 ;
      RECT 9.210000 3.480000 9.990000 3.810000 ;
    LAYER met4 ;
      RECT 9.010000 -0.155000 10.190000 1.025000 ;
      RECT 9.010000  3.045000 10.190000 4.225000 ;
    LAYER via ;
      RECT 5.600000 1.905000 5.860000 2.165000 ;
      RECT 5.920000 1.905000 6.180000 2.165000 ;
      RECT 9.310000 0.305000 9.570000 0.565000 ;
      RECT 9.310000 3.505000 9.570000 3.765000 ;
      RECT 9.630000 0.305000 9.890000 0.565000 ;
      RECT 9.630000 3.505000 9.890000 3.765000 ;
    LAYER via2 ;
      RECT 5.485000 1.895000 5.765000 2.175000 ;
      RECT 5.885000 1.895000 6.165000 2.175000 ;
      RECT 9.260000 0.285000 9.540000 0.565000 ;
      RECT 9.260000 3.505000 9.540000 3.785000 ;
      RECT 9.660000 0.285000 9.940000 0.565000 ;
      RECT 9.660000 3.505000 9.940000 3.785000 ;
    LAYER via3 ;
      RECT 2.865000 1.875000 3.185000 2.195000 ;
      RECT 3.265000 1.875000 3.585000 2.195000 ;
      RECT 5.465000 1.875000 5.785000 2.195000 ;
      RECT 5.865000 1.875000 6.185000 2.195000 ;
      RECT 9.240000 0.265000 9.560000 0.585000 ;
      RECT 9.240000 3.485000 9.560000 3.805000 ;
      RECT 9.640000 0.265000 9.960000 0.585000 ;
      RECT 9.640000 3.485000 9.960000 3.805000 ;
  END
END sky130_fd_sc_hvl__probec_p_8
MACRO sky130_fd_sc_hvl__dfsbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__dfsbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  17.76000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN D
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.515000 2.875000 2.145000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.498750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 17.300000 0.495000 17.635000 1.325000 ;
        RECT 17.300000 2.355000 17.635000 3.435000 ;
        RECT 17.405000 1.325000 17.635000 2.355000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.641250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.015000 0.495000 15.375000 3.755000 ;
    END
  END Q_N
  PIN SET_B
    ANTENNAGATEAREA  0.840000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  6.985000 1.155000 10.330000 1.325000 ;
        RECT 10.160000 1.325000 10.330000 1.605000 ;
        RECT 10.160000 1.605000 10.885000 1.775000 ;
        RECT 10.715000 1.775000 10.885000 1.975000 ;
        RECT 10.715000 1.975000 12.830000 2.145000 ;
        RECT 12.150000 1.555000 12.830000 1.975000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.560000 1.550000 0.890000 2.520000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 17.760000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 17.760000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 17.760000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 17.760000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000  5.990000 2.385000 ;
        RECT -0.330000 2.385000 18.090000 4.485000 ;
        RECT 11.500000 1.885000 18.090000 2.385000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 17.760000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 17.760000 0.085000 ;
      RECT  0.000000  3.985000 17.760000 4.155000 ;
      RECT  0.110000  0.540000  0.360000 1.200000 ;
      RECT  0.110000  1.200000  1.590000 1.370000 ;
      RECT  0.110000  1.370000  0.380000 3.450000 ;
      RECT  0.540000  0.365000  1.490000 1.020000 ;
      RECT  0.650000  2.700000  1.240000 3.705000 ;
      RECT  1.260000  1.370000  1.590000 1.870000 ;
      RECT  1.420000  1.870000  1.590000 3.630000 ;
      RECT  1.420000  3.630000  2.290000 3.800000 ;
      RECT  1.670000  0.540000  2.000000 1.000000 ;
      RECT  1.770000  1.000000  2.000000 1.165000 ;
      RECT  1.770000  1.165000  2.820000 1.335000 ;
      RECT  1.770000  1.335000  1.940000 3.450000 ;
      RECT  2.120000  2.325000  3.025000 2.495000 ;
      RECT  2.120000  2.495000  2.290000 3.630000 ;
      RECT  2.220000  0.365000  2.470000 0.985000 ;
      RECT  2.470000  2.675000  2.675000 3.705000 ;
      RECT  2.650000  0.265000  4.460000 0.435000 ;
      RECT  2.650000  0.435000  2.820000 1.165000 ;
      RECT  2.855000  2.495000  3.025000 3.355000 ;
      RECT  2.855000  3.355000  5.500000 3.525000 ;
      RECT  3.000000  0.615000  3.375000 1.005000 ;
      RECT  3.205000  1.005000  3.375000 2.675000 ;
      RECT  3.205000  2.675000  3.545000 3.175000 ;
      RECT  3.555000  1.105000  3.725000 2.225000 ;
      RECT  3.555000  2.225000  4.800000 2.395000 ;
      RECT  3.725000  2.395000  3.895000 3.355000 ;
      RECT  3.780000  0.615000  4.110000 0.925000 ;
      RECT  3.905000  0.925000  4.075000 1.855000 ;
      RECT  3.905000  1.855000  8.060000 2.025000 ;
      RECT  4.075000  2.675000  4.405000 3.005000 ;
      RECT  4.075000  3.005000  5.150000 3.175000 ;
      RECT  4.255000  1.105000  4.585000 1.505000 ;
      RECT  4.255000  1.505000  9.470000 1.675000 ;
      RECT  4.290000  0.435000  4.460000 1.105000 ;
      RECT  4.585000  2.395000  4.800000 2.555000 ;
      RECT  4.650000  0.365000  5.600000 0.905000 ;
      RECT  4.945000  1.085000  6.150000 1.325000 ;
      RECT  4.980000  2.025000  5.150000 3.005000 ;
      RECT  5.330000  2.205000  7.025000 2.375000 ;
      RECT  5.330000  2.555000  6.595000 2.725000 ;
      RECT  5.330000  2.725000  5.500000 3.355000 ;
      RECT  5.680000  2.905000  6.245000 3.705000 ;
      RECT  5.820000  0.515000  6.150000 1.085000 ;
      RECT  6.425000  2.725000  6.595000 3.355000 ;
      RECT  6.425000  3.355000  7.675000 3.525000 ;
      RECT  6.775000  2.375000  7.025000 3.175000 ;
      RECT  6.785000  0.365000  7.735000 0.975000 ;
      RECT  7.505000  2.545000  9.120000 2.715000 ;
      RECT  7.505000  2.715000  7.675000 3.355000 ;
      RECT  7.730000  2.025000  8.060000 2.365000 ;
      RECT  7.855000  2.895000  8.805000 3.705000 ;
      RECT  8.185000  0.375000 11.110000 0.545000 ;
      RECT  8.185000  0.545000  8.515000 0.975000 ;
      RECT  8.755000  0.725000 10.680000 0.975000 ;
      RECT  8.870000  1.885000  9.120000 2.545000 ;
      RECT  9.300000  1.675000  9.470000 2.305000 ;
      RECT  9.300000  2.305000 10.185000 2.475000 ;
      RECT  9.345000  2.675000  9.675000 3.585000 ;
      RECT  9.345000  3.585000 10.535000 3.755000 ;
      RECT  9.650000  1.505000  9.980000 1.955000 ;
      RECT  9.650000  1.955000 10.535000 2.125000 ;
      RECT  9.855000  2.475000 10.185000 2.555000 ;
      RECT 10.365000  2.125000 10.535000 2.325000 ;
      RECT 10.365000  2.325000 13.180000 2.495000 ;
      RECT 10.365000  2.495000 10.535000 3.585000 ;
      RECT 10.510000  0.975000 10.680000 1.255000 ;
      RECT 10.510000  1.255000 11.460000 1.425000 ;
      RECT 10.715000  2.675000 11.665000 3.705000 ;
      RECT 10.860000  0.545000 11.110000 1.075000 ;
      RECT 11.290000  0.515000 11.660000 0.975000 ;
      RECT 11.290000  0.975000 11.460000 1.255000 ;
      RECT 11.640000  1.155000 11.970000 1.205000 ;
      RECT 11.640000  1.205000 14.395000 1.375000 ;
      RECT 11.640000  1.375000 11.970000 1.795000 ;
      RECT 12.035000  2.495000 13.180000 3.175000 ;
      RECT 12.200000  0.365000 13.150000 0.975000 ;
      RECT 13.010000  1.555000 14.045000 1.725000 ;
      RECT 13.010000  1.725000 13.180000 2.325000 ;
      RECT 13.360000  1.905000 14.395000 2.075000 ;
      RECT 13.360000  2.075000 13.690000 2.675000 ;
      RECT 13.390000  0.825000 13.720000 1.205000 ;
      RECT 13.870000  2.255000 14.820000 3.755000 ;
      RECT 13.900000  0.365000 14.835000 1.025000 ;
      RECT 14.225000  1.375000 14.395000 1.905000 ;
      RECT 15.625000  0.825000 15.975000 1.505000 ;
      RECT 15.625000  1.505000 17.175000 1.675000 ;
      RECT 15.625000  1.675000 15.955000 3.185000 ;
      RECT 16.135000  2.355000 17.085000 3.705000 ;
      RECT 16.155000  0.365000 17.105000 1.305000 ;
      RECT 16.845000  1.675000 17.175000 2.175000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.985000  0.325000 4.155000 ;
      RECT  0.570000  0.395000  0.740000 0.565000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.985000  0.805000 4.155000 ;
      RECT  0.680000  3.505000  0.850000 3.675000 ;
      RECT  0.930000  0.395000  1.100000 0.565000 ;
      RECT  1.040000  3.505000  1.210000 3.675000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.985000  1.285000 4.155000 ;
      RECT  1.290000  0.395000  1.460000 0.565000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.985000  1.765000 4.155000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.985000  2.245000 4.155000 ;
      RECT  2.250000  0.395000  2.420000 0.565000 ;
      RECT  2.490000  3.505000  2.660000 3.675000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.985000  2.725000 4.155000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.985000  3.205000 4.155000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.985000  3.685000 4.155000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.985000  4.165000 4.155000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.985000  4.645000 4.155000 ;
      RECT  4.680000  0.395000  4.850000 0.565000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.985000  5.125000 4.155000 ;
      RECT  5.040000  0.395000  5.210000 0.565000 ;
      RECT  5.400000  0.395000  5.570000 0.565000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.985000  5.605000 4.155000 ;
      RECT  5.695000  3.505000  5.865000 3.675000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.985000  6.085000 4.155000 ;
      RECT  6.055000  3.505000  6.225000 3.675000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.985000  6.565000 4.155000 ;
      RECT  6.815000  0.395000  6.985000 0.565000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.985000  7.045000 4.155000 ;
      RECT  7.175000  0.395000  7.345000 0.565000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.985000  7.525000 4.155000 ;
      RECT  7.535000  0.395000  7.705000 0.565000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.985000  8.005000 4.155000 ;
      RECT  7.885000  3.505000  8.055000 3.675000 ;
      RECT  8.245000  3.505000  8.415000 3.675000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.985000  8.485000 4.155000 ;
      RECT  8.605000  3.505000  8.775000 3.675000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.985000  8.965000 4.155000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.985000  9.445000 4.155000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.985000  9.925000 4.155000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.985000 10.405000 4.155000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.985000 10.885000 4.155000 ;
      RECT 10.745000  3.505000 10.915000 3.675000 ;
      RECT 11.105000  3.505000 11.275000 3.675000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.985000 11.365000 4.155000 ;
      RECT 11.465000  3.505000 11.635000 3.675000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.985000 11.845000 4.155000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.985000 12.325000 4.155000 ;
      RECT 12.230000  0.395000 12.400000 0.565000 ;
      RECT 12.590000  0.395000 12.760000 0.565000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.985000 12.805000 4.155000 ;
      RECT 12.950000  0.395000 13.120000 0.565000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.985000 13.285000 4.155000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.985000 13.765000 4.155000 ;
      RECT 13.900000  3.505000 14.070000 3.675000 ;
      RECT 13.920000  0.395000 14.090000 0.565000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.985000 14.245000 4.155000 ;
      RECT 14.260000  3.505000 14.430000 3.675000 ;
      RECT 14.280000  0.395000 14.450000 0.565000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.985000 14.725000 4.155000 ;
      RECT 14.620000  3.505000 14.790000 3.675000 ;
      RECT 14.640000  0.395000 14.810000 0.565000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.985000 15.205000 4.155000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.985000 15.685000 4.155000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000  3.985000 16.165000 4.155000 ;
      RECT 16.165000  3.505000 16.335000 3.675000 ;
      RECT 16.185000  0.395000 16.355000 0.565000 ;
      RECT 16.475000 -0.085000 16.645000 0.085000 ;
      RECT 16.475000  3.985000 16.645000 4.155000 ;
      RECT 16.525000  3.505000 16.695000 3.675000 ;
      RECT 16.545000  0.395000 16.715000 0.565000 ;
      RECT 16.885000  3.505000 17.055000 3.675000 ;
      RECT 16.905000  0.395000 17.075000 0.565000 ;
      RECT 16.955000 -0.085000 17.125000 0.085000 ;
      RECT 16.955000  3.985000 17.125000 4.155000 ;
      RECT 17.435000 -0.085000 17.605000 0.085000 ;
      RECT 17.435000  3.985000 17.605000 4.155000 ;
  END
END sky130_fd_sc_hvl__dfsbp_1
MACRO sky130_fd_sc_hvl__dlrtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__dlrtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.600000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN D
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.570000 1.930000 0.900000 2.600000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.641250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.735000 2.175000 9.475000 3.755000 ;
        RECT 9.140000 0.495000 9.475000 2.175000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.515000 0.810000 8.120000 1.780000 ;
        RECT 7.515000 1.780000 7.845000 1.855000 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.175000 1.795000 1.400000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 9.600000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 9.600000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 9.600000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 9.600000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 9.930000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 9.600000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.600000 0.085000 ;
      RECT 0.000000  3.985000 9.600000 4.155000 ;
      RECT 0.140000  0.495000 0.390000 1.580000 ;
      RECT 0.140000  1.580000 1.795000 1.675000 ;
      RECT 0.140000  1.675000 3.655000 1.750000 ;
      RECT 0.140000  1.750000 0.390000 3.610000 ;
      RECT 0.570000  0.365000 1.520000 0.995000 ;
      RECT 0.570000  2.780000 1.520000 3.705000 ;
      RECT 1.625000  1.750000 3.655000 1.845000 ;
      RECT 1.700000  0.495000 2.145000 0.995000 ;
      RECT 1.700000  2.025000 4.435000 2.195000 ;
      RECT 1.700000  2.195000 2.030000 3.610000 ;
      RECT 1.975000  0.995000 2.145000 1.325000 ;
      RECT 1.975000  1.325000 4.005000 1.495000 ;
      RECT 2.290000  2.375000 4.785000 2.545000 ;
      RECT 2.290000  2.545000 2.620000 3.245000 ;
      RECT 2.370000  0.495000 2.620000 0.975000 ;
      RECT 2.370000  0.975000 4.495000 1.145000 ;
      RECT 2.800000  0.365000 3.750000 0.795000 ;
      RECT 2.800000  2.725000 3.750000 3.705000 ;
      RECT 3.835000  1.495000 4.005000 1.605000 ;
      RECT 3.835000  1.605000 4.435000 2.025000 ;
      RECT 4.185000  1.145000 4.495000 1.225000 ;
      RECT 4.185000  1.225000 4.785000 1.395000 ;
      RECT 4.560000  2.725000 5.525000 2.895000 ;
      RECT 4.560000  2.895000 4.890000 3.245000 ;
      RECT 4.615000  1.395000 4.785000 1.965000 ;
      RECT 4.615000  1.965000 5.175000 2.295000 ;
      RECT 4.615000  2.295000 4.785000 2.375000 ;
      RECT 4.675000  0.495000 5.135000 0.995000 ;
      RECT 4.965000  0.995000 5.135000 1.175000 ;
      RECT 4.965000  1.175000 6.780000 1.345000 ;
      RECT 5.355000  1.345000 5.525000 2.725000 ;
      RECT 5.545000  0.365000 6.495000 0.995000 ;
      RECT 5.705000  2.255000 6.655000 3.705000 ;
      RECT 5.810000  1.525000 6.140000 1.905000 ;
      RECT 5.810000  1.905000 7.130000 2.035000 ;
      RECT 5.810000  2.035000 8.470000 2.075000 ;
      RECT 6.450000  1.345000 6.780000 1.725000 ;
      RECT 6.755000  0.495000 7.130000 0.995000 ;
      RECT 6.960000  0.995000 7.130000 1.905000 ;
      RECT 6.960000  2.075000 8.470000 2.205000 ;
      RECT 6.960000  2.205000 7.390000 3.005000 ;
      RECT 7.570000  2.385000 8.520000 3.755000 ;
      RECT 8.300000  0.365000 8.890000 1.325000 ;
      RECT 8.300000  1.665000 8.630000 1.995000 ;
      RECT 8.300000  1.995000 8.470000 2.035000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.600000  0.395000 0.770000 0.565000 ;
      RECT 0.600000  3.505000 0.770000 3.675000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.960000  0.395000 1.130000 0.565000 ;
      RECT 0.960000  3.505000 1.130000 3.675000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.320000  0.395000 1.490000 0.565000 ;
      RECT 1.320000  3.505000 1.490000 3.675000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 2.830000  0.395000 3.000000 0.565000 ;
      RECT 2.830000  3.505000 3.000000 3.675000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
      RECT 3.190000  0.395000 3.360000 0.565000 ;
      RECT 3.190000  3.505000 3.360000 3.675000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.985000 3.685000 4.155000 ;
      RECT 3.550000  0.395000 3.720000 0.565000 ;
      RECT 3.550000  3.505000 3.720000 3.675000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.985000 4.165000 4.155000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.985000 4.645000 4.155000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.985000 5.125000 4.155000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.985000 5.605000 4.155000 ;
      RECT 5.575000  0.395000 5.745000 0.565000 ;
      RECT 5.735000  3.505000 5.905000 3.675000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.985000 6.085000 4.155000 ;
      RECT 5.935000  0.395000 6.105000 0.565000 ;
      RECT 6.095000  3.505000 6.265000 3.675000 ;
      RECT 6.295000  0.395000 6.465000 0.565000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.985000 6.565000 4.155000 ;
      RECT 6.455000  3.505000 6.625000 3.675000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.985000 7.045000 4.155000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.985000 7.525000 4.155000 ;
      RECT 7.600000  3.505000 7.770000 3.675000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.985000 8.005000 4.155000 ;
      RECT 7.960000  3.505000 8.130000 3.675000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.985000 8.485000 4.155000 ;
      RECT 8.320000  3.505000 8.490000 3.675000 ;
      RECT 8.330000  0.395000 8.500000 0.565000 ;
      RECT 8.690000  0.395000 8.860000 0.565000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.985000 8.965000 4.155000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.985000 9.445000 4.155000 ;
  END
END sky130_fd_sc_hvl__dlrtp_1
MACRO sky130_fd_sc_hvl__o21ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__o21ai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A1
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.505000 0.855000 1.835000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 1.505000 1.795000 1.760000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.325000 1.805000 3.235000 2.120000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.633750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.940000 2.145000 2.110000 ;
        RECT 1.565000 2.110000 2.040000 3.755000 ;
        RECT 1.975000 1.455000 2.820000 1.625000 ;
        RECT 1.975000 1.625000 2.145000 1.940000 ;
        RECT 2.490000 0.495000 2.820000 1.455000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 3.360000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 3.360000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 3.360000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 3.360000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 3.690000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 3.360000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.985000 3.360000 4.155000 ;
      RECT 0.090000  2.175000 1.040000 3.755000 ;
      RECT 0.130000  0.495000 0.460000 1.105000 ;
      RECT 0.130000  1.105000 2.040000 1.275000 ;
      RECT 0.130000  1.275000 0.460000 1.325000 ;
      RECT 0.640000  0.365000 1.530000 0.925000 ;
      RECT 1.710000  0.495000 2.040000 1.105000 ;
      RECT 2.220000  2.300000 3.170000 3.755000 ;
    LAYER mcon ;
      RECT 0.120000  3.505000 0.290000 3.675000 ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.480000  3.505000 0.650000 3.675000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.640000  0.395000 0.810000 0.565000 ;
      RECT 0.840000  3.505000 1.010000 3.675000 ;
      RECT 1.000000  0.395000 1.170000 0.565000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.360000  0.395000 1.530000 0.565000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.250000  3.505000 2.420000 3.675000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 2.610000  3.505000 2.780000 3.675000 ;
      RECT 2.970000  3.505000 3.140000 3.675000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
  END
END sky130_fd_sc_hvl__o21ai_1
MACRO sky130_fd_sc_hvl__sdfrbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__sdfrbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  20.16000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN D
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.625000 2.330000 2.135000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.626250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 19.700000 0.685000 20.040000 3.755000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.596250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 17.435000 0.515000 17.835000 3.570000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  5.235000 1.295000  5.635000 2.150000 ;
        RECT 10.685000 1.625000 11.245000 2.135000 ;
      LAYER mcon ;
        RECT  5.435000 1.950000  5.605000 2.120000 ;
        RECT 10.715000 1.950000 10.885000 2.120000 ;
    END
    PORT
      LAYER li1 ;
        RECT 15.005000 1.425000 15.685000 2.120000 ;
      LAYER mcon ;
        RECT 15.035000 1.950000 15.205000 2.120000 ;
    END
    PORT
      LAYER met1 ;
        RECT  5.375000 1.920000  5.665000 1.965000 ;
        RECT  5.375000 1.965000 15.265000 2.105000 ;
        RECT  5.375000 2.105000  5.665000 2.150000 ;
        RECT 10.655000 1.920000 10.945000 1.965000 ;
        RECT 10.655000 2.105000 10.945000 2.150000 ;
        RECT 14.975000 1.920000 15.265000 1.965000 ;
        RECT 14.975000 2.105000 15.265000 2.150000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.710000 1.975000 4.705000 2.155000 ;
        RECT 3.710000 2.155000 4.040000 2.480000 ;
        RECT 4.375000 1.295000 4.705000 1.975000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.840000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.655000 1.295000 0.985000 1.965000 ;
        RECT 0.815000 0.265000 1.685000 0.435000 ;
        RECT 0.815000 0.435000 0.985000 1.295000 ;
        RECT 1.515000 0.435000 1.685000 1.275000 ;
        RECT 1.515000 1.275000 4.195000 1.445000 ;
        RECT 1.515000 2.665000 3.040000 2.835000 ;
        RECT 1.515000 2.835000 1.765000 2.995000 ;
        RECT 3.485000 1.445000 4.195000 1.795000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 5.870000 1.850000 6.200000 2.520000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 20.160000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 20.160000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 20.160000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 20.160000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 20.490000 4.485000 ;
        RECT 16.405000 1.720000 18.095000 1.885000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 20.160000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 20.160000 0.085000 ;
      RECT  0.000000  3.985000 20.160000 4.155000 ;
      RECT  0.090000  0.365000  0.635000 1.115000 ;
      RECT  0.090000  3.205000  0.985000 3.705000 ;
      RECT  1.165000  0.615000  1.335000 2.315000 ;
      RECT  1.165000  2.315000  3.440000 2.485000 ;
      RECT  1.165000  2.485000  1.335000 3.205000 ;
      RECT  1.165000  3.205000  1.415000 3.705000 ;
      RECT  1.675000  3.235000  2.115000 3.735000 ;
      RECT  1.865000  0.265000  5.095000 0.435000 ;
      RECT  1.865000  0.435000  2.115000 0.995000 ;
      RECT  1.945000  3.015000  6.325000 3.185000 ;
      RECT  1.945000  3.185000  2.115000 3.235000 ;
      RECT  2.545000  3.365000  3.495000 3.735000 ;
      RECT  2.730000  1.625000  3.060000 2.315000 ;
      RECT  3.270000  2.485000  3.440000 2.665000 ;
      RECT  3.270000  2.665000  4.680000 2.835000 ;
      RECT  3.275000  0.615000  3.605000 0.925000 ;
      RECT  3.275000  0.925000  5.055000 1.095000 ;
      RECT  4.350000  2.325000  4.680000 2.665000 ;
      RECT  4.655000  3.185000  4.905000 3.735000 ;
      RECT  4.765000  0.435000  5.095000 0.755000 ;
      RECT  4.885000  1.095000  5.055000 3.015000 ;
      RECT  5.085000  3.365000  5.975000 3.755000 ;
      RECT  5.275000  0.365000  6.225000 0.995000 ;
      RECT  6.155000  3.185000  6.325000 3.635000 ;
      RECT  6.155000  3.635000  7.025000 3.805000 ;
      RECT  6.505000  0.495000  6.675000 1.505000 ;
      RECT  6.505000  1.505000  7.695000 1.675000 ;
      RECT  6.505000  1.675000  6.675000 3.455000 ;
      RECT  6.855000  1.855000  7.725000 2.025000 ;
      RECT  6.855000  2.025000  7.025000 3.635000 ;
      RECT  6.870000  0.365000  7.720000 0.915000 ;
      RECT  7.205000  2.205000  7.375000 3.705000 ;
      RECT  7.365000  1.345000  7.695000 1.505000 ;
      RECT  7.555000  2.025000  7.725000 3.255000 ;
      RECT  7.555000  3.255000  8.955000 3.425000 ;
      RECT  7.900000  0.265000  9.975000 0.435000 ;
      RECT  7.900000  0.435000  8.150000 0.995000 ;
      RECT  7.905000  0.995000  8.150000 2.225000 ;
      RECT  7.905000  2.225000  8.605000 3.015000 ;
      RECT  8.275000  3.425000  8.605000 3.755000 ;
      RECT  8.355000  3.015000  8.605000 3.075000 ;
      RECT  8.410000  0.615000  8.955000 0.995000 ;
      RECT  8.785000  0.995000  8.955000 3.255000 ;
      RECT  9.135000  0.615000  9.520000 0.995000 ;
      RECT  9.135000  0.995000  9.305000 2.905000 ;
      RECT  9.135000  2.905000 11.775000 3.075000 ;
      RECT  9.135000  3.075000  9.385000 3.755000 ;
      RECT  9.510000  2.005000  9.840000 2.315000 ;
      RECT  9.510000  2.315000 11.595000 2.485000 ;
      RECT  9.510000  2.485000  9.840000 2.675000 ;
      RECT  9.700000  0.435000  9.975000 0.925000 ;
      RECT  9.700000  0.925000 12.145000 1.095000 ;
      RECT  9.700000  1.095000  9.975000 1.755000 ;
      RECT  9.925000  3.255000 10.875000 3.755000 ;
      RECT 10.225000  1.275000 12.645000 1.445000 ;
      RECT 10.225000  1.445000 10.505000 1.945000 ;
      RECT 10.770000  0.365000 11.805000 0.745000 ;
      RECT 11.325000  2.665000 11.945000 2.835000 ;
      RECT 11.325000  2.835000 11.775000 2.905000 ;
      RECT 11.325000  3.075000 11.775000 3.735000 ;
      RECT 11.425000  1.875000 12.295000 2.045000 ;
      RECT 11.425000  2.045000 11.595000 2.315000 ;
      RECT 11.775000  2.225000 11.945000 2.665000 ;
      RECT 11.955000  3.015000 12.545000 3.735000 ;
      RECT 11.975000  0.265000 14.270000 0.435000 ;
      RECT 11.975000  0.435000 12.145000 0.925000 ;
      RECT 12.125000  2.045000 12.295000 2.175000 ;
      RECT 12.125000  2.175000 13.220000 2.345000 ;
      RECT 12.315000  0.615000 12.645000 1.275000 ;
      RECT 12.475000  1.445000 12.645000 1.825000 ;
      RECT 12.475000  1.825000 13.570000 1.995000 ;
      RECT 12.735000  2.525000 13.570000 2.695000 ;
      RECT 12.735000  2.695000 12.985000 3.755000 ;
      RECT 12.825000  0.435000 12.995000 1.475000 ;
      RECT 12.825000  1.475000 13.155000 1.645000 ;
      RECT 13.175000  0.615000 13.425000 1.125000 ;
      RECT 13.175000  1.125000 13.920000 1.295000 ;
      RECT 13.400000  1.995000 13.570000 2.525000 ;
      RECT 13.435000  2.875000 14.620000 3.045000 ;
      RECT 13.435000  3.045000 13.765000 3.755000 ;
      RECT 13.750000  1.295000 13.920000 2.875000 ;
      RECT 14.100000  0.435000 14.270000 2.555000 ;
      RECT 14.450000  0.365000 15.400000 0.895000 ;
      RECT 14.450000  1.075000 16.195000 1.245000 ;
      RECT 14.450000  1.245000 14.620000 2.875000 ;
      RECT 14.800000  2.300000 16.150000 2.495000 ;
      RECT 14.800000  2.675000 15.720000 3.705000 ;
      RECT 15.865000  1.245000 16.195000 1.655000 ;
      RECT 15.900000  2.495000 16.150000 3.175000 ;
      RECT 15.980000  1.835000 16.545000 2.005000 ;
      RECT 15.980000  2.005000 16.150000 2.300000 ;
      RECT 16.175000  0.515000 16.545000 0.895000 ;
      RECT 16.330000  2.185000 17.255000 3.705000 ;
      RECT 16.375000  0.895000 16.545000 1.835000 ;
      RECT 16.725000  0.365000 17.255000 1.305000 ;
      RECT 18.025000  0.685000 18.385000 1.655000 ;
      RECT 18.025000  1.655000 19.520000 1.985000 ;
      RECT 18.025000  1.985000 18.355000 2.985000 ;
      RECT 18.535000  2.175000 19.485000 3.755000 ;
      RECT 18.565000  0.365000 19.515000 1.475000 ;
    LAYER mcon ;
      RECT  0.095000  0.395000  0.265000 0.565000 ;
      RECT  0.095000  3.505000  0.265000 3.675000 ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.985000  0.325000 4.155000 ;
      RECT  0.455000  0.395000  0.625000 0.565000 ;
      RECT  0.455000  3.505000  0.625000 3.675000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.985000  0.805000 4.155000 ;
      RECT  0.815000  3.505000  0.985000 3.675000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.985000  1.285000 4.155000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.985000  1.765000 4.155000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.985000  2.245000 4.155000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.985000  2.725000 4.155000 ;
      RECT  2.575000  3.505000  2.745000 3.675000 ;
      RECT  2.935000  3.505000  3.105000 3.675000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.985000  3.205000 4.155000 ;
      RECT  3.295000  3.505000  3.465000 3.675000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.985000  3.685000 4.155000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.985000  4.165000 4.155000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.985000  4.645000 4.155000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.985000  5.125000 4.155000 ;
      RECT  5.085000  3.505000  5.255000 3.675000 ;
      RECT  5.305000  0.395000  5.475000 0.565000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.985000  5.605000 4.155000 ;
      RECT  5.445000  3.505000  5.615000 3.675000 ;
      RECT  5.665000  0.395000  5.835000 0.565000 ;
      RECT  5.805000  3.505000  5.975000 3.675000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.985000  6.085000 4.155000 ;
      RECT  6.025000  0.395000  6.195000 0.565000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.985000  6.565000 4.155000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.985000  7.045000 4.155000 ;
      RECT  6.950000  0.395000  7.120000 0.565000 ;
      RECT  7.205000  3.505000  7.375000 3.675000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.985000  7.525000 4.155000 ;
      RECT  7.470000  0.395000  7.640000 0.565000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.985000  8.005000 4.155000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.985000  8.485000 4.155000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.985000  8.965000 4.155000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.985000  9.445000 4.155000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.985000  9.925000 4.155000 ;
      RECT  9.955000  3.505000 10.125000 3.675000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.985000 10.405000 4.155000 ;
      RECT 10.315000  3.505000 10.485000 3.675000 ;
      RECT 10.675000  3.505000 10.845000 3.675000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.985000 10.885000 4.155000 ;
      RECT 10.800000  0.395000 10.970000 0.565000 ;
      RECT 11.160000  0.395000 11.330000 0.565000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.985000 11.365000 4.155000 ;
      RECT 11.520000  0.395000 11.690000 0.565000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.985000 11.845000 4.155000 ;
      RECT 11.985000  3.505000 12.155000 3.675000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.985000 12.325000 4.155000 ;
      RECT 12.345000  3.505000 12.515000 3.675000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.985000 12.805000 4.155000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.985000 13.285000 4.155000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.985000 13.765000 4.155000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.985000 14.245000 4.155000 ;
      RECT 14.480000  0.395000 14.650000 0.565000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.985000 14.725000 4.155000 ;
      RECT 14.815000  3.505000 14.985000 3.675000 ;
      RECT 14.840000  0.395000 15.010000 0.565000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.985000 15.205000 4.155000 ;
      RECT 15.175000  3.505000 15.345000 3.675000 ;
      RECT 15.200000  0.395000 15.370000 0.565000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.985000 15.685000 4.155000 ;
      RECT 15.535000  3.505000 15.705000 3.675000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000  3.985000 16.165000 4.155000 ;
      RECT 16.345000  3.505000 16.515000 3.675000 ;
      RECT 16.475000 -0.085000 16.645000 0.085000 ;
      RECT 16.475000  3.985000 16.645000 4.155000 ;
      RECT 16.705000  3.505000 16.875000 3.675000 ;
      RECT 16.725000  0.395000 16.895000 0.565000 ;
      RECT 16.955000 -0.085000 17.125000 0.085000 ;
      RECT 16.955000  3.985000 17.125000 4.155000 ;
      RECT 17.065000  3.505000 17.235000 3.675000 ;
      RECT 17.085000  0.395000 17.255000 0.565000 ;
      RECT 17.435000 -0.085000 17.605000 0.085000 ;
      RECT 17.435000  3.985000 17.605000 4.155000 ;
      RECT 17.915000 -0.085000 18.085000 0.085000 ;
      RECT 17.915000  3.985000 18.085000 4.155000 ;
      RECT 18.395000 -0.085000 18.565000 0.085000 ;
      RECT 18.395000  3.985000 18.565000 4.155000 ;
      RECT 18.565000  3.505000 18.735000 3.675000 ;
      RECT 18.595000  0.395000 18.765000 0.565000 ;
      RECT 18.875000 -0.085000 19.045000 0.085000 ;
      RECT 18.875000  3.985000 19.045000 4.155000 ;
      RECT 18.925000  3.505000 19.095000 3.675000 ;
      RECT 18.955000  0.395000 19.125000 0.565000 ;
      RECT 19.285000  3.505000 19.455000 3.675000 ;
      RECT 19.315000  0.395000 19.485000 0.565000 ;
      RECT 19.355000 -0.085000 19.525000 0.085000 ;
      RECT 19.355000  3.985000 19.525000 4.155000 ;
      RECT 19.835000 -0.085000 20.005000 0.085000 ;
      RECT 19.835000  3.985000 20.005000 4.155000 ;
  END
END sky130_fd_sc_hvl__sdfrbp_1
MACRO sky130_fd_sc_hvl__nand3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__nand3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.455000 0.810000 2.725000 1.725000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.885000 0.810000 2.275000 1.725000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.505000 0.995000 1.835000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  1.065000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.200000 1.905000 3.235000 2.075000 ;
        RECT 1.200000 2.075000 1.370000 3.755000 ;
        RECT 2.905000 0.495000 3.235000 1.325000 ;
        RECT 2.980000 1.325000 3.235000 1.905000 ;
        RECT 2.980000 2.075000 3.235000 3.755000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 3.360000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 3.360000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 3.360000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 3.360000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 3.690000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 3.360000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.985000 3.360000 4.155000 ;
      RECT 0.090000  0.365000 1.705000 1.325000 ;
      RECT 0.090000  2.175000 1.020000 3.755000 ;
      RECT 1.550000  2.255000 2.800000 3.755000 ;
    LAYER mcon ;
      RECT 0.095000  0.395000 0.265000 0.565000 ;
      RECT 0.110000  3.505000 0.280000 3.675000 ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.455000  0.395000 0.625000 0.565000 ;
      RECT 0.470000  3.505000 0.640000 3.675000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.815000  0.395000 0.985000 0.565000 ;
      RECT 0.830000  3.505000 1.000000 3.675000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.175000  0.395000 1.345000 0.565000 ;
      RECT 1.535000  0.395000 1.705000 0.565000 ;
      RECT 1.550000  3.505000 1.720000 3.675000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.910000  3.505000 2.080000 3.675000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.270000  3.505000 2.440000 3.675000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 2.630000  3.505000 2.800000 3.675000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
  END
END sky130_fd_sc_hvl__nand3_1
MACRO sky130_fd_sc_hvl__o22ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__o22ai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A1
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.805000 3.715000 2.120000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.250000 1.805000 2.755000 2.120000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.535000 0.550000 1.865000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.535000 1.595000 1.750000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.742500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.735000 0.615000 1.270000 1.355000 ;
        RECT 0.735000 1.355000 0.905000 1.930000 ;
        RECT 0.735000 1.930000 1.795000 2.100000 ;
        RECT 1.525000 2.100000 1.795000 2.175000 ;
        RECT 1.525000 2.175000 2.045000 3.260000 ;
        RECT 1.875000 3.260000 2.045000 3.755000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 3.840000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 3.840000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 3.840000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 3.840000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 4.170000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 3.840000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.985000 3.840000 4.155000 ;
      RECT 0.090000  2.280000 1.345000 3.755000 ;
      RECT 0.160000  0.265000 1.970000 0.435000 ;
      RECT 0.160000  0.435000 0.490000 1.355000 ;
      RECT 1.800000  0.435000 1.970000 1.455000 ;
      RECT 1.800000  1.455000 3.670000 1.625000 ;
      RECT 2.150000  0.365000 3.250000 1.275000 ;
      RECT 2.305000  2.300000 3.615000 3.755000 ;
      RECT 3.420000  0.525000 3.670000 1.455000 ;
    LAYER mcon ;
      RECT 0.095000  3.505000 0.265000 3.675000 ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.455000  3.505000 0.625000 3.675000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.815000  3.505000 0.985000 3.675000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.175000  3.505000 1.345000 3.675000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.200000  0.395000 2.370000 0.565000 ;
      RECT 2.335000  3.505000 2.505000 3.675000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 2.560000  0.395000 2.730000 0.565000 ;
      RECT 2.695000  3.505000 2.865000 3.675000 ;
      RECT 2.920000  0.395000 3.090000 0.565000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
      RECT 3.055000  3.505000 3.225000 3.675000 ;
      RECT 3.415000  3.505000 3.585000 3.675000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.985000 3.685000 4.155000 ;
  END
END sky130_fd_sc_hvl__o22ai_1
MACRO sky130_fd_sc_hvl__mux2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__mux2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A0
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.295000 1.785000 2.905000 1.955000 ;
        RECT 2.295000 1.955000 2.625000 2.235000 ;
        RECT 2.735000 1.095000 3.685000 1.390000 ;
        RECT 2.735000 1.390000 2.905000 1.785000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.085000 1.570000 3.685000 1.955000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.840000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435000 1.705000 1.765000 3.095000 ;
        RECT 1.435000 3.095000 3.230000 3.265000 ;
        RECT 3.060000 2.135000 4.675000 2.305000 ;
        RECT 3.060000 2.305000 3.230000 3.095000 ;
        RECT 4.365000 1.550000 4.675000 2.135000 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  0.641250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.495000 0.415000 1.925000 ;
        RECT 0.125000 1.925000 0.495000 3.755000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 5.280000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 5.280000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 5.280000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 5.280000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 5.610000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 5.280000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.280000 0.085000 ;
      RECT 0.000000  3.985000 5.280000 4.155000 ;
      RECT 0.595000  0.365000 2.205000 1.175000 ;
      RECT 0.620000  1.355000 2.555000 1.525000 ;
      RECT 0.620000  1.525000 0.950000 1.745000 ;
      RECT 0.675000  2.175000 1.255000 3.755000 ;
      RECT 1.945000  1.525000 2.115000 2.415000 ;
      RECT 1.945000  2.415000 2.880000 2.585000 ;
      RECT 2.385000  0.495000 2.880000 0.915000 ;
      RECT 2.385000  0.915000 2.555000 1.355000 ;
      RECT 2.550000  2.585000 2.880000 2.915000 ;
      RECT 3.060000  0.365000 4.720000 0.915000 ;
      RECT 3.410000  2.495000 4.720000 3.705000 ;
      RECT 3.865000  1.105000 5.150000 1.275000 ;
      RECT 3.865000  1.275000 4.115000 1.775000 ;
      RECT 4.900000  0.495000 5.150000 1.105000 ;
      RECT 4.900000  1.275000 5.150000 2.915000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.595000  0.395000 0.765000 0.565000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.700000  3.505000 0.870000 3.675000 ;
      RECT 0.955000  0.395000 1.125000 0.565000 ;
      RECT 1.060000  3.505000 1.230000 3.675000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.315000  0.395000 1.485000 0.565000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.675000  0.395000 1.845000 0.565000 ;
      RECT 2.035000  0.395000 2.205000 0.565000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
      RECT 3.085000  0.395000 3.255000 0.565000 ;
      RECT 3.440000  3.505000 3.610000 3.675000 ;
      RECT 3.445000  0.395000 3.615000 0.565000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.985000 3.685000 4.155000 ;
      RECT 3.800000  3.505000 3.970000 3.675000 ;
      RECT 3.805000  0.395000 3.975000 0.565000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.985000 4.165000 4.155000 ;
      RECT 4.160000  3.505000 4.330000 3.675000 ;
      RECT 4.165000  0.395000 4.335000 0.565000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.985000 4.645000 4.155000 ;
      RECT 4.520000  3.505000 4.690000 3.675000 ;
      RECT 4.525000  0.395000 4.695000 0.565000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.985000 5.125000 4.155000 ;
  END
END sky130_fd_sc_hvl__mux2_1
MACRO sky130_fd_sc_hvl__conb_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__conb_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.400000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN HI
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.290000 0.430000 0.865000 1.070000 ;
        RECT 0.615000 1.070000 0.865000 1.935000 ;
        RECT 0.615000 1.935000 1.325000 2.185000 ;
        RECT 1.075000 2.185000 1.325000 3.530000 ;
    END
  END HI
  PIN LO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.035000 0.500000 1.365000 1.500000 ;
        RECT 1.035000 1.500000 1.795000 1.765000 ;
        RECT 1.530000 1.765000 1.795000 3.175000 ;
        RECT 1.530000 3.175000 2.110000 3.815000 ;
    END
  END LO
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 2.400000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 2.400000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 2.400000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 2.400000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 2.730000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 2.400000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.400000 0.085000 ;
      RECT 0.000000  3.985000 2.400000 4.155000 ;
      RECT 0.215000  3.175000 0.620000 3.445000 ;
      RECT 0.215000  3.445000 0.865000 3.785000 ;
      RECT 1.535000  0.285000 2.185000 0.625000 ;
      RECT 1.780000  0.625000 2.185000 1.070000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.275000  3.505000 0.445000 3.675000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.505000 0.805000 3.675000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  0.395000 1.765000 0.565000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.955000  0.395000 2.125000 0.565000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
  END
END sky130_fd_sc_hvl__conb_1
MACRO sky130_fd_sc_hvl__lsbuflv2hv_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__lsbuflv2hv_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.56000 BY  8.140000 ;
  SYMMETRY X Y ;
  SITE unithvdbl ;
  PIN A
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.495000 1.530000 2.805000 2.200000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.596250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.120000 4.405000 10.450000 6.055000 ;
        RECT 10.120000 6.725000 10.450000 7.625000 ;
        RECT 10.210000 6.055000 10.450000 6.725000 ;
    END
  END X
  PIN LVPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.070000 3.020000 10.490000 3.305000 ;
      LAYER nwell ;
        RECT 2.800000 2.015000 4.335000 4.325000 ;
    END
  END LVPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 7.515000 10.560000 7.885000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 8.025000 10.560000 8.255000 ;
      LAYER pwell ;
        RECT 0.000000 8.055000 10.560000 8.225000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 10.560000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000  0.800000 6.255000 ;
        RECT  6.335000 2.465000 10.890000 6.255000 ;
        RECT  9.800000 1.885000 10.890000 2.465000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 4.325000 10.560000 4.695000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.560000 0.085000 ;
      RECT 0.000000  3.985000  0.800000 4.155000 ;
      RECT 0.000000  8.055000 10.560000 8.225000 ;
      RECT 1.585000  6.085000  2.175000 7.715000 ;
      RECT 1.585000  7.715000  5.295000 7.885000 ;
      RECT 2.495000  5.665000  7.990000 5.995000 ;
      RECT 2.495000  5.995000  2.825000 7.545000 ;
      RECT 2.885000  2.765000  3.265000 3.055000 ;
      RECT 2.885000  3.055000  3.175000 5.495000 ;
      RECT 2.975000  0.735000  3.265000 1.745000 ;
      RECT 2.975000  1.745000  4.310000 1.995000 ;
      RECT 2.975000  1.995000  3.265000 2.765000 ;
      RECT 3.095000  0.335000  4.045000 0.565000 ;
      RECT 3.145000  6.165000  3.735000 7.715000 ;
      RECT 3.345000  3.225000  4.115000 4.200000 ;
      RECT 3.435000  0.565000  3.705000 1.575000 ;
      RECT 3.435000  2.165000  3.705000 3.075000 ;
      RECT 3.435000  3.075000  4.115000 3.225000 ;
      RECT 3.875000  0.735000  4.185000 1.245000 ;
      RECT 3.875000  1.245000  4.810000 1.575000 ;
      RECT 3.875000  2.165000  5.790000 2.475000 ;
      RECT 3.875000  2.475000  4.185000 2.905000 ;
      RECT 4.055000  5.995000  4.385000 7.545000 ;
      RECT 4.480000  1.575000  4.810000 2.145000 ;
      RECT 4.480000  2.145000  5.790000 2.165000 ;
      RECT 4.705000  6.165000  5.295000 7.715000 ;
      RECT 5.050000  0.255000  8.760000 0.425000 ;
      RECT 5.050000  0.425000  5.640000 1.975000 ;
      RECT 5.615000  5.995000  5.945000 7.625000 ;
      RECT 5.960000  0.595000  6.290000 2.145000 ;
      RECT 5.960000  2.145000  9.410000 2.475000 ;
      RECT 6.185000  3.135000  6.995000 3.465000 ;
      RECT 6.185000  3.465000  6.515000 5.665000 ;
      RECT 6.610000  0.425000  7.200000 1.975000 ;
      RECT 6.665000  2.795000  6.995000 3.135000 ;
      RECT 6.685000  4.470000  7.495000 4.800000 ;
      RECT 7.165000  2.475000  7.495000 3.395000 ;
      RECT 7.165000  3.395000  7.835000 3.805000 ;
      RECT 7.165000  3.805000  7.495000 4.470000 ;
      RECT 7.520000  0.595000  7.850000 2.145000 ;
      RECT 7.660000  5.205000  7.990000 5.665000 ;
      RECT 7.660000  5.995000  7.990000 6.555000 ;
      RECT 7.755000  3.985000 10.560000 4.155000 ;
      RECT 7.755000  4.405000  8.345000 4.800000 ;
      RECT 8.005000  2.795000  8.595000 3.705000 ;
      RECT 8.170000  0.425000  8.760000 1.975000 ;
      RECT 8.515000  4.405000  8.845000 6.225000 ;
      RECT 8.515000  6.225000 10.040000 6.555000 ;
      RECT 8.515000  6.555000  8.845000 7.625000 ;
      RECT 9.080000  0.515000  9.410000 2.145000 ;
      RECT 9.210000  4.405000  9.800000 5.945000 ;
      RECT 9.210000  6.835000  9.800000 7.745000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.985000  0.325000 4.155000 ;
      RECT  0.155000  8.055000  0.325000 8.225000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  8.055000  0.805000 8.225000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  8.055000  1.285000 8.225000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  8.055000  1.765000 8.225000 ;
      RECT  1.615000  7.545000  1.785000 7.715000 ;
      RECT  1.975000  7.545000  2.145000 7.715000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  8.055000  2.245000 8.225000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  8.055000  2.725000 8.225000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  8.055000  3.205000 8.225000 ;
      RECT  3.125000  0.365000  3.295000 0.535000 ;
      RECT  3.175000  7.545000  3.345000 7.715000 ;
      RECT  3.485000  0.425000  3.655000 0.595000 ;
      RECT  3.485000  3.050000  3.655000 3.220000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  8.055000  3.685000 8.225000 ;
      RECT  3.535000  7.545000  3.705000 7.715000 ;
      RECT  3.845000  0.365000  4.015000 0.535000 ;
      RECT  3.845000  3.105000  4.015000 3.275000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  8.055000  4.165000 8.225000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  8.055000  4.645000 8.225000 ;
      RECT  4.735000  7.545000  4.905000 7.715000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  8.055000  5.125000 8.225000 ;
      RECT  5.080000  0.425000  5.250000 0.595000 ;
      RECT  5.095000  7.545000  5.265000 7.715000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  8.055000  5.605000 8.225000 ;
      RECT  5.440000  0.425000  5.610000 0.595000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  8.055000  6.085000 8.225000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  8.055000  6.565000 8.225000 ;
      RECT  6.640000  0.425000  6.810000 0.595000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  8.055000  7.045000 8.225000 ;
      RECT  7.000000  0.425000  7.170000 0.595000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  8.055000  7.525000 8.225000 ;
      RECT  7.785000  4.495000  7.955000 4.665000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.985000  8.005000 4.155000 ;
      RECT  7.835000  8.055000  8.005000 8.225000 ;
      RECT  8.035000  3.475000  8.205000 3.645000 ;
      RECT  8.145000  4.495000  8.315000 4.665000 ;
      RECT  8.200000  0.425000  8.370000 0.595000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.985000  8.485000 4.155000 ;
      RECT  8.315000  8.055000  8.485000 8.225000 ;
      RECT  8.395000  3.475000  8.565000 3.645000 ;
      RECT  8.560000  0.425000  8.730000 0.595000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.985000  8.965000 4.155000 ;
      RECT  8.795000  8.055000  8.965000 8.225000 ;
      RECT  9.240000  4.495000  9.410000 4.665000 ;
      RECT  9.240000  7.545000  9.410000 7.715000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.985000  9.445000 4.155000 ;
      RECT  9.275000  8.055000  9.445000 8.225000 ;
      RECT  9.600000  4.495000  9.770000 4.665000 ;
      RECT  9.600000  7.545000  9.770000 7.715000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.985000  9.925000 4.155000 ;
      RECT  9.755000  8.055000  9.925000 8.225000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.985000 10.405000 4.155000 ;
      RECT 10.235000  8.055000 10.405000 8.225000 ;
    LAYER met1 ;
      RECT 0.000000 -0.115000 10.560000 0.115000 ;
      RECT 0.000000  0.255000 10.560000 0.625000 ;
      RECT 0.000000  3.445000 10.560000 3.815000 ;
    LAYER pwell ;
      RECT 0.000000 -0.085000 10.560000 0.085000 ;
  END
END sky130_fd_sc_hvl__lsbuflv2hv_1
MACRO sky130_fd_sc_hvl__lsbuflv2hv_isosrchvaon_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__lsbuflv2hv_isosrchvaon_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.92000 BY  8.140000 ;
  SYMMETRY X Y ;
  SITE unithvdbl ;
  PIN A
    ANTENNAGATEAREA  0.279000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.205000 1.685000 9.895000 2.015000 ;
    END
  END A
  PIN SLEEP_B
    ANTENNAGATEAREA  7.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.730000 1.830000 5.400000 2.160000 ;
    END
  END SLEEP_B
  PIN X
    ANTENNADIFFAREA  0.397500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.755000 1.315000 1.175000 1.605000 ;
        RECT 0.755000 1.605000 0.975000 2.405000 ;
        RECT 0.755000 2.405000 1.175000 2.695000 ;
        RECT 0.955000 0.895000 1.175000 1.315000 ;
        RECT 0.955000 2.695000 1.175000 3.075000 ;
    END
  END X
  PIN LVPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.070000 3.020000 13.850000 3.305000 ;
      LAYER nwell ;
        RECT 8.890000 2.045000 10.710000 6.095000 ;
    END
  END LVPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 7.515000 13.920000 7.885000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 8.025000 13.920000 8.255000 ;
      LAYER pwell ;
        RECT 0.000000 8.055000 13.920000 8.225000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 13.920000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 0.510000 2.095000 ;
        RECT -0.330000 2.095000 6.020000 6.005000 ;
        RECT -0.330000 6.005000 0.510000 6.255000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 4.325000 13.920000 4.695000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.920000 0.085000 ;
      RECT  0.000000  3.985000  0.685000 4.155000 ;
      RECT  0.000000  8.055000 13.920000 8.225000 ;
      RECT  0.360000  4.155000  0.530000 5.280000 ;
      RECT  0.895000  4.575000  2.780000 4.795000 ;
      RECT  0.895000  4.795000  1.115000 6.055000 ;
      RECT  0.895000  6.055000  1.955000 6.275000 ;
      RECT  0.955000  6.445000  1.175000 7.625000 ;
      RECT  0.955000  7.625000  4.900000 7.845000 ;
      RECT  1.365000  5.555000  2.035000 5.665000 ;
      RECT  1.365000  5.665000  5.675000 5.885000 ;
      RECT  1.400000  0.395000  1.990000 0.625000 ;
      RECT  1.735000  6.275000  1.955000 7.455000 ;
      RECT  1.760000  0.625000  1.990000 1.565000 ;
      RECT  1.760000  2.405000  1.930000 3.445000 ;
      RECT  1.760000  3.445000  2.350000 3.735000 ;
      RECT  2.110000  4.295000  2.780000 4.575000 ;
      RECT  2.260000  0.645000  2.480000 2.860000 ;
      RECT  2.260000  2.860000  2.780000 3.085000 ;
      RECT  2.515000  6.445000  2.735000 7.625000 ;
      RECT  2.560000  3.085000  2.780000 4.295000 ;
      RECT  2.650000  1.830000  3.320000 1.940000 ;
      RECT  2.650000  1.940000  4.425000 2.160000 ;
      RECT  3.060000  3.445000  3.645000 3.735000 ;
      RECT  3.175000  0.395000  3.765000 0.625000 ;
      RECT  3.175000  4.410000  3.645000 4.630000 ;
      RECT  3.175000  4.630000  3.395000 5.405000 ;
      RECT  3.295000  5.885000  3.515000 7.455000 ;
      RECT  3.360000  0.625000  3.590000 1.655000 ;
      RECT  3.425000  2.405000  3.645000 3.445000 ;
      RECT  3.425000  3.735000  3.645000 4.410000 ;
      RECT  4.075000  6.445000  4.295000 7.625000 ;
      RECT  4.205000  0.645000  4.425000 1.940000 ;
      RECT  4.205000  2.160000  4.425000 3.755000 ;
      RECT  4.680000  6.295000  8.445000 6.515000 ;
      RECT  4.680000  6.515000  4.900000 7.625000 ;
      RECT  5.455000  4.945000  5.675000 5.665000 ;
      RECT  6.465000  1.305000  6.685000 6.295000 ;
      RECT  7.155000  0.395000  7.745000 0.625000 ;
      RECT  7.340000  0.625000  7.570000 6.055000 ;
      RECT  7.750000  7.075000  9.535000 7.405000 ;
      RECT  8.225000  1.305000  8.445000 6.295000 ;
      RECT  9.100000  3.905000 10.035000 4.235000 ;
      RECT  9.205000  4.775000  9.535000 7.075000 ;
      RECT  9.305000  0.395000  9.895000 0.625000 ;
      RECT  9.305000  3.020000  9.895000 3.365000 ;
      RECT  9.565000  0.625000  9.895000 1.515000 ;
      RECT  9.565000  2.335000  9.895000 3.020000 ;
      RECT  9.565000  3.365000  9.895000 3.905000 ;
      RECT  9.705000  4.235000 10.035000 5.805000 ;
      RECT  9.705000  6.125000 10.535000 6.455000 ;
      RECT  9.705000  6.625000 10.035000 7.520000 ;
      RECT  9.705000  7.520000 10.295000 7.750000 ;
      RECT 10.065000  0.735000 10.395000 3.035000 ;
      RECT 10.065000  3.035000 10.535000 3.365000 ;
      RECT 10.205000  3.365000 10.535000 6.125000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.985000  0.325000 4.155000 ;
      RECT  0.155000  8.055000  0.325000 8.225000 ;
      RECT  0.515000  3.985000  0.685000 4.155000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  8.055000  0.805000 8.225000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  8.055000  1.285000 8.225000 ;
      RECT  1.430000  0.425000  1.600000 0.595000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  8.055000  1.765000 8.225000 ;
      RECT  1.790000  0.425000  1.960000 0.595000 ;
      RECT  1.790000  3.505000  1.960000 3.675000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  8.055000  2.245000 8.225000 ;
      RECT  2.150000  3.505000  2.320000 3.675000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  8.055000  2.725000 8.225000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  8.055000  3.205000 8.225000 ;
      RECT  3.090000  3.505000  3.260000 3.675000 ;
      RECT  3.205000  0.425000  3.375000 0.595000 ;
      RECT  3.450000  3.505000  3.620000 3.675000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  8.055000  3.685000 8.225000 ;
      RECT  3.565000  0.425000  3.735000 0.595000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  8.055000  4.165000 8.225000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  8.055000  4.645000 8.225000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  8.055000  5.125000 8.225000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  8.055000  5.605000 8.225000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  8.055000  6.085000 8.225000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  8.055000  6.565000 8.225000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  8.055000  7.045000 8.225000 ;
      RECT  7.185000  0.425000  7.355000 0.595000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  8.055000  7.525000 8.225000 ;
      RECT  7.545000  0.425000  7.715000 0.595000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  8.055000  8.005000 8.225000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  8.055000  8.485000 8.225000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  8.055000  8.965000 8.225000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  8.055000  9.445000 8.225000 ;
      RECT  9.335000  0.425000  9.505000 0.595000 ;
      RECT  9.335000  3.080000  9.505000 3.250000 ;
      RECT  9.695000  0.425000  9.865000 0.595000 ;
      RECT  9.695000  3.080000  9.865000 3.250000 ;
      RECT  9.735000  7.550000  9.905000 7.720000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  8.055000  9.925000 8.225000 ;
      RECT 10.095000  7.550000 10.265000 7.720000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  8.055000 10.405000 8.225000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  8.055000 10.885000 8.225000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  8.055000 11.365000 8.225000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  8.055000 11.845000 8.225000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  8.055000 12.325000 8.225000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  8.055000 12.805000 8.225000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  8.055000 13.285000 8.225000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  8.055000 13.765000 8.225000 ;
    LAYER met1 ;
      RECT 0.000000 -0.115000 13.920000 0.115000 ;
      RECT 0.000000  0.255000 13.920000 0.625000 ;
      RECT 0.000000  3.445000 13.920000 3.815000 ;
    LAYER pwell ;
      RECT 0.000000 -0.085000 13.920000 0.085000 ;
  END
END sky130_fd_sc_hvl__lsbuflv2hv_isosrchvaon_1
MACRO sky130_fd_sc_hvl__lsbufhv2hv_hl_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__lsbufhv2hv_hl_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  8.140000 ;
  SYMMETRY X Y ;
  SITE unithvdbl ;
  PIN A
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.355000 1.775000 4.685000 2.900000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.626250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.995000 0.495000 3.395000 4.065000 ;
    END
  END X
  PIN LOWHVPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.070000 3.020000 8.570000 3.305000 ;
      LAYER nwell ;
        RECT 2.800000 1.885000 5.425000 5.135000 ;
    END
  END LOWHVPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 7.515000 8.640000 7.885000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 8.025000 8.640000 8.255000 ;
      LAYER pwell ;
        RECT 0.000000 8.055000 8.640000 8.225000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 8.640000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 0.800000 6.255000 ;
        RECT  7.425000 1.885000 8.970000 6.255000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 4.325000 8.640000 4.695000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.640000 0.085000 ;
      RECT 0.000000  3.985000 0.800000 4.155000 ;
      RECT 0.000000  8.055000 8.640000 8.225000 ;
      RECT 3.130000  4.265000 5.095000 4.835000 ;
      RECT 3.565000  0.365000 4.515000 1.265000 ;
      RECT 3.565000  1.435000 5.115000 1.605000 ;
      RECT 3.565000  1.605000 3.895000 2.065000 ;
      RECT 3.565000  2.485000 4.185000 4.265000 ;
      RECT 4.865000  0.495000 5.115000 1.435000 ;
      RECT 4.865000  1.605000 5.115000 3.315000 ;
      RECT 7.425000  3.985000 8.640000 4.155000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.155000  8.055000 0.325000 8.225000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  8.055000 0.805000 8.225000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  8.055000 1.285000 8.225000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  8.055000 1.765000 8.225000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  8.055000 2.245000 8.225000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  8.055000 2.725000 8.225000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  8.055000 3.205000 8.225000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  8.055000 3.685000 8.225000 ;
      RECT 3.595000  0.395000 3.765000 0.565000 ;
      RECT 3.630000  3.075000 3.800000 3.245000 ;
      RECT 3.955000  0.395000 4.125000 0.565000 ;
      RECT 3.990000  3.075000 4.160000 3.245000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  8.055000 4.165000 8.225000 ;
      RECT 4.315000  0.395000 4.485000 0.565000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  8.055000 4.645000 8.225000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  8.055000 5.125000 8.225000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  8.055000 5.605000 8.225000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  8.055000 6.085000 8.225000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  8.055000 6.565000 8.225000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  8.055000 7.045000 8.225000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  8.055000 7.525000 8.225000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.985000 8.005000 4.155000 ;
      RECT 7.835000  8.055000 8.005000 8.225000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.985000 8.485000 4.155000 ;
      RECT 8.315000  8.055000 8.485000 8.225000 ;
    LAYER met1 ;
      RECT 0.000000 -0.115000 8.640000 0.115000 ;
      RECT 0.000000  0.255000 8.640000 0.625000 ;
      RECT 0.000000  3.445000 8.640000 3.815000 ;
    LAYER pwell ;
      RECT 0.000000 -0.085000 8.640000 0.085000 ;
  END
END sky130_fd_sc_hvl__lsbufhv2hv_hl_1
MACRO sky130_fd_sc_hvl__lsbufhv2hv_lh_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__lsbufhv2hv_lh_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.56000 BY  8.140000 ;
  SYMMETRY X Y ;
  SITE unithvdbl ;
  PIN A
    ANTENNAGATEAREA  0.750000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.495000 1.530000 2.805000 2.200000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.596250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.120000 4.405000 10.450000 7.625000 ;
    END
  END X
  PIN LOWHVPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.070000 3.020000 10.490000 3.305000 ;
      LAYER nwell ;
        RECT 2.800000 2.015000 5.270000 4.315000 ;
    END
  END LOWHVPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 7.515000 10.560000 7.885000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 8.025000 10.560000 8.255000 ;
      LAYER pwell ;
        RECT 0.000000 8.055000 10.560000 8.225000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 10.560000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000  0.800000 6.255000 ;
        RECT  7.270000 2.465000 10.890000 6.255000 ;
        RECT  9.800000 1.885000 10.890000 2.465000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 4.325000 10.560000 4.695000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.560000 0.085000 ;
      RECT 0.000000  3.985000  0.800000 4.155000 ;
      RECT 0.000000  8.055000 10.560000 8.225000 ;
      RECT 3.090000  0.685000  3.420000 1.745000 ;
      RECT 3.090000  1.745000  4.845000 1.995000 ;
      RECT 3.090000  1.995000  3.420000 5.165000 ;
      RECT 3.090000  5.165000  5.660000 5.495000 ;
      RECT 3.300000  6.085000  3.890000 7.715000 ;
      RECT 3.300000  7.715000  7.010000 7.885000 ;
      RECT 3.590000  3.355000  4.780000 4.025000 ;
      RECT 3.740000  0.255000  9.540000 0.425000 ;
      RECT 3.740000  0.425000  4.330000 1.475000 ;
      RECT 3.740000  2.325000  4.330000 3.355000 ;
      RECT 4.210000  5.665000  7.930000 5.995000 ;
      RECT 4.210000  5.995000  4.540000 7.545000 ;
      RECT 4.650000  0.685000  4.980000 1.145000 ;
      RECT 4.650000  1.145000  5.660000 1.475000 ;
      RECT 4.650000  2.165000  6.570000 2.475000 ;
      RECT 4.650000  2.475000  4.980000 3.115000 ;
      RECT 4.860000  6.165000  5.450000 7.715000 ;
      RECT 5.330000  1.475000  5.660000 2.145000 ;
      RECT 5.330000  2.145000  6.570000 2.165000 ;
      RECT 5.770000  5.995000  6.100000 7.545000 ;
      RECT 5.830000  0.425000  6.420000 1.975000 ;
      RECT 6.420000  6.165000  7.010000 7.715000 ;
      RECT 6.740000  0.595000  7.070000 2.145000 ;
      RECT 6.740000  2.145000  8.630000 2.475000 ;
      RECT 7.375000  3.605000  8.045000 3.935000 ;
      RECT 7.390000  0.425000  7.980000 1.975000 ;
      RECT 7.600000  2.795000  8.545000 3.125000 ;
      RECT 7.600000  3.125000  7.930000 3.435000 ;
      RECT 7.600000  3.935000  7.930000 5.665000 ;
      RECT 8.215000  2.475000  8.545000 2.795000 ;
      RECT 8.215000  3.125000  8.545000 5.205000 ;
      RECT 8.215000  5.205000  8.965000 5.535000 ;
      RECT 8.300000  0.595000  8.630000 2.145000 ;
      RECT 8.635000  5.535000  8.965000 6.555000 ;
      RECT 8.715000  3.985000 10.560000 4.155000 ;
      RECT 8.790000  4.405000  9.800000 4.800000 ;
      RECT 8.940000  2.795000  9.530000 3.705000 ;
      RECT 8.950000  0.425000  9.540000 1.975000 ;
      RECT 9.210000  4.800000  9.800000 5.945000 ;
      RECT 9.210000  6.835000  9.800000 7.745000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.985000  0.325000 4.155000 ;
      RECT  0.155000  8.055000  0.325000 8.225000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  8.055000  0.805000 8.225000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  8.055000  1.285000 8.225000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  8.055000  1.765000 8.225000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  8.055000  2.245000 8.225000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  8.055000  2.725000 8.225000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  8.055000  3.205000 8.225000 ;
      RECT  3.330000  7.545000  3.500000 7.715000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  8.055000  3.685000 8.225000 ;
      RECT  3.690000  7.545000  3.860000 7.715000 ;
      RECT  3.770000  0.425000  3.940000 0.595000 ;
      RECT  3.770000  3.050000  3.940000 3.220000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  8.055000  4.165000 8.225000 ;
      RECT  4.130000  0.425000  4.300000 0.595000 ;
      RECT  4.130000  3.050000  4.300000 3.220000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  8.055000  4.645000 8.225000 ;
      RECT  4.890000  7.545000  5.060000 7.715000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  8.055000  5.125000 8.225000 ;
      RECT  5.250000  7.545000  5.420000 7.715000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  8.055000  5.605000 8.225000 ;
      RECT  5.860000  0.425000  6.030000 0.595000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  8.055000  6.085000 8.225000 ;
      RECT  6.220000  0.425000  6.390000 0.595000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  8.055000  6.565000 8.225000 ;
      RECT  6.450000  7.545000  6.620000 7.715000 ;
      RECT  6.810000  7.545000  6.980000 7.715000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  8.055000  7.045000 8.225000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  8.055000  7.525000 8.225000 ;
      RECT  7.420000  0.425000  7.590000 0.595000 ;
      RECT  7.780000  0.425000  7.950000 0.595000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  8.055000  8.005000 8.225000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  8.055000  8.485000 8.225000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.985000  8.965000 4.155000 ;
      RECT  8.795000  8.055000  8.965000 8.225000 ;
      RECT  8.880000  4.495000  9.050000 4.665000 ;
      RECT  8.970000  3.475000  9.140000 3.645000 ;
      RECT  8.980000  0.425000  9.150000 0.595000 ;
      RECT  9.240000  4.495000  9.410000 4.665000 ;
      RECT  9.240000  7.545000  9.410000 7.715000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.985000  9.445000 4.155000 ;
      RECT  9.275000  8.055000  9.445000 8.225000 ;
      RECT  9.330000  3.475000  9.500000 3.645000 ;
      RECT  9.340000  0.425000  9.510000 0.595000 ;
      RECT  9.600000  4.495000  9.770000 4.665000 ;
      RECT  9.600000  7.545000  9.770000 7.715000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.985000  9.925000 4.155000 ;
      RECT  9.755000  8.055000  9.925000 8.225000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.985000 10.405000 4.155000 ;
      RECT 10.235000  8.055000 10.405000 8.225000 ;
    LAYER met1 ;
      RECT 0.000000 -0.115000 10.560000 0.115000 ;
      RECT 0.000000  0.255000 10.560000 0.625000 ;
      RECT 0.000000  3.445000 10.560000 3.815000 ;
    LAYER pwell ;
      RECT 0.000000 -0.085000 10.560000 0.085000 ;
  END
END sky130_fd_sc_hvl__lsbufhv2hv_lh_1
MACRO sky130_fd_sc_hvl__lsbuflv2hv_symmetric_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__lsbuflv2hv_symmetric_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  8.140000 ;
  SYMMETRY X Y ;
  SITE unithvdbl ;
  PIN A
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.495000 1.530000 2.805000 2.200000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.596250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.600000 4.405000 10.930000 6.055000 ;
        RECT 10.600000 6.725000 10.930000 7.625000 ;
        RECT 10.690000 6.055000 10.930000 6.725000 ;
    END
  END X
  PIN LVPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.070000 3.020000 10.970000 3.305000 ;
      LAYER nwell ;
        RECT 2.800000 2.015000 4.335000 4.325000 ;
    END
  END LVPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 7.515000 11.040000 7.885000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 8.025000 11.040000 8.255000 ;
      LAYER pwell ;
        RECT 0.000000 8.055000 11.040000 8.225000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 11.040000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000  0.800000 6.255000 ;
        RECT  6.335000 2.465000 11.370000 6.255000 ;
        RECT  9.800000 1.885000 11.370000 2.465000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 4.325000 11.040000 4.695000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  3.985000  0.800000 4.155000 ;
      RECT  0.000000  8.055000 11.040000 8.225000 ;
      RECT  2.885000  2.765000  3.265000 3.055000 ;
      RECT  2.885000  3.055000  3.175000 5.495000 ;
      RECT  2.975000  0.735000  3.265000 1.745000 ;
      RECT  2.975000  1.745000  4.310000 1.995000 ;
      RECT  2.975000  1.995000  3.265000 2.765000 ;
      RECT  3.095000  0.335000  4.045000 0.565000 ;
      RECT  3.145000  6.165000  3.735000 7.715000 ;
      RECT  3.145000  7.715000  5.295000 7.885000 ;
      RECT  3.345000  3.225000  4.115000 4.200000 ;
      RECT  3.435000  0.565000  3.705000 1.575000 ;
      RECT  3.435000  2.165000  3.705000 3.075000 ;
      RECT  3.435000  3.075000  4.115000 3.225000 ;
      RECT  3.875000  0.735000  4.185000 1.245000 ;
      RECT  3.875000  1.245000  4.810000 1.575000 ;
      RECT  3.875000  2.165000  5.790000 2.475000 ;
      RECT  3.875000  2.475000  4.185000 2.905000 ;
      RECT  4.055000  5.665000  7.025000 5.995000 ;
      RECT  4.055000  5.995000  4.385000 7.545000 ;
      RECT  4.480000  1.575000  4.810000 2.145000 ;
      RECT  4.480000  2.145000  5.790000 2.165000 ;
      RECT  4.705000  6.165000  5.295000 7.715000 ;
      RECT  5.050000  0.255000  7.200000 0.425000 ;
      RECT  5.050000  0.425000  5.640000 1.975000 ;
      RECT  5.960000  0.595000  6.290000 2.145000 ;
      RECT  5.960000  2.145000  7.850000 2.325000 ;
      RECT  6.565000  2.795000  6.895000 4.405000 ;
      RECT  6.565000  4.405000  7.025000 4.735000 ;
      RECT  6.610000  0.425000  7.200000 1.975000 ;
      RECT  6.695000  4.735000  7.025000 5.665000 ;
      RECT  6.695000  5.995000  7.025000 6.285000 ;
      RECT  6.695000  6.285000  8.815000 6.615000 ;
      RECT  7.095000  2.495000  9.835000 2.705000 ;
      RECT  7.095000  2.705000  7.765000 4.215000 ;
      RECT  7.390000  4.405000  7.980000 5.945000 ;
      RECT  7.520000  0.255000  9.410000 0.425000 ;
      RECT  7.520000  0.425000  7.850000 2.145000 ;
      RECT  7.955000  2.875000  8.545000 3.705000 ;
      RECT  8.170000  0.595000  8.760000 2.495000 ;
      RECT  8.235000  3.985000 11.040000 4.155000 ;
      RECT  8.300000  4.405000  8.630000 6.285000 ;
      RECT  8.535000  6.615000  8.815000 6.955000 ;
      RECT  8.915000  2.705000  9.835000 3.465000 ;
      RECT  8.995000  4.405000  9.325000 6.225000 ;
      RECT  8.995000  6.225000 10.520000 6.555000 ;
      RECT  8.995000  6.555000  9.325000 7.625000 ;
      RECT  9.080000  0.425000  9.410000 2.055000 ;
      RECT  9.690000  4.405000 10.280000 5.945000 ;
      RECT  9.690000  6.835000 10.280000 7.745000 ;
      RECT 10.125000  2.795000 10.715000 3.705000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.985000  0.325000 4.155000 ;
      RECT  0.155000  8.055000  0.325000 8.225000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  8.055000  0.805000 8.225000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  8.055000  1.285000 8.225000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  8.055000  1.765000 8.225000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  8.055000  2.245000 8.225000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  8.055000  2.725000 8.225000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  8.055000  3.205000 8.225000 ;
      RECT  3.125000  0.365000  3.295000 0.535000 ;
      RECT  3.175000  7.545000  3.345000 7.715000 ;
      RECT  3.485000  0.425000  3.655000 0.595000 ;
      RECT  3.485000  3.050000  3.655000 3.220000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  8.055000  3.685000 8.225000 ;
      RECT  3.535000  7.545000  3.705000 7.715000 ;
      RECT  3.845000  0.365000  4.015000 0.535000 ;
      RECT  3.845000  3.105000  4.015000 3.275000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  8.055000  4.165000 8.225000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  8.055000  4.645000 8.225000 ;
      RECT  4.735000  7.545000  4.905000 7.715000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  8.055000  5.125000 8.225000 ;
      RECT  5.080000  0.425000  5.250000 0.595000 ;
      RECT  5.095000  7.545000  5.265000 7.715000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  8.055000  5.605000 8.225000 ;
      RECT  5.440000  0.425000  5.610000 0.595000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  8.055000  6.085000 8.225000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  8.055000  6.565000 8.225000 ;
      RECT  6.640000  0.425000  6.810000 0.595000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  8.055000  7.045000 8.225000 ;
      RECT  7.000000  0.425000  7.170000 0.595000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  8.055000  7.525000 8.225000 ;
      RECT  7.420000  4.495000  7.590000 4.665000 ;
      RECT  7.780000  4.495000  7.950000 4.665000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  8.055000  8.005000 8.225000 ;
      RECT  7.985000  3.475000  8.155000 3.645000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.985000  8.485000 4.155000 ;
      RECT  8.315000  8.055000  8.485000 8.225000 ;
      RECT  8.345000  3.475000  8.515000 3.645000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.985000  8.965000 4.155000 ;
      RECT  8.795000  8.055000  8.965000 8.225000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.985000  9.445000 4.155000 ;
      RECT  9.275000  8.055000  9.445000 8.225000 ;
      RECT  9.720000  4.495000  9.890000 4.665000 ;
      RECT  9.720000  7.545000  9.890000 7.715000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.985000  9.925000 4.155000 ;
      RECT  9.755000  8.055000  9.925000 8.225000 ;
      RECT 10.080000  4.495000 10.250000 4.665000 ;
      RECT 10.080000  7.545000 10.250000 7.715000 ;
      RECT 10.155000  3.475000 10.325000 3.645000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.985000 10.405000 4.155000 ;
      RECT 10.235000  8.055000 10.405000 8.225000 ;
      RECT 10.515000  3.475000 10.685000 3.645000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.985000 10.885000 4.155000 ;
      RECT 10.715000  8.055000 10.885000 8.225000 ;
    LAYER met1 ;
      RECT 0.000000 -0.115000 11.040000 0.115000 ;
      RECT 0.000000  0.255000 11.040000 0.625000 ;
      RECT 0.000000  3.445000 11.040000 3.815000 ;
    LAYER pwell ;
      RECT 0.000000 -0.085000 11.040000 0.085000 ;
  END
END sky130_fd_sc_hvl__lsbuflv2hv_symmetric_1
MACRO sky130_fd_sc_hvl__dfrtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__dfrtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  15.36000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN D
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.415000 0.810000 3.745000 2.105000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.611250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.900000 0.665000 15.235000 3.735000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  2.695000 1.620000  3.235000 2.490000 ;
        RECT  3.065000 0.460000  6.010000 0.630000 ;
        RECT  3.065000 0.630000  3.235000 1.620000 ;
        RECT  5.840000 0.630000  6.010000 1.125000 ;
        RECT  5.840000 1.125000  8.460000 1.295000 ;
        RECT  6.605000 1.825000  8.460000 1.995000 ;
        RECT  8.290000 0.265000 10.950000 0.435000 ;
        RECT  8.290000 0.435000  8.460000 1.125000 ;
        RECT  8.290000 1.295000  8.460000 1.825000 ;
        RECT 10.780000 0.435000 10.950000 1.095000 ;
        RECT 10.780000 1.095000 11.785000 1.265000 ;
        RECT 11.455000 1.265000 11.785000 1.655000 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.560000 1.175000 0.890000 2.150000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 15.360000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 15.360000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 15.360000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 15.360000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 15.690000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 15.360000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 15.360000 0.085000 ;
      RECT  0.000000  3.985000 15.360000 4.155000 ;
      RECT  0.110000  0.495000  0.380000 2.355000 ;
      RECT  0.110000  2.355000  1.570000 2.525000 ;
      RECT  0.110000  2.525000  0.440000 3.455000 ;
      RECT  0.560000  0.365000  1.510000 0.995000 ;
      RECT  0.630000  2.725000  1.220000 3.705000 ;
      RECT  1.240000  1.855000  1.570000 2.355000 ;
      RECT  1.400000  2.525000  1.570000 3.635000 ;
      RECT  1.400000  3.635000  2.840000 3.805000 ;
      RECT  1.690000  0.495000  2.020000 0.995000 ;
      RECT  1.750000  0.995000  2.020000 1.920000 ;
      RECT  1.750000  1.920000  2.275000 2.150000 ;
      RECT  1.750000  2.150000  2.000000 3.455000 ;
      RECT  2.200000  0.365000  2.790000 1.245000 ;
      RECT  2.240000  2.670000  4.050000 2.840000 ;
      RECT  2.240000  2.840000  2.490000 3.455000 ;
      RECT  2.670000  3.020000  3.700000 3.190000 ;
      RECT  2.670000  3.190000  2.840000 3.635000 ;
      RECT  3.020000  3.370000  3.350000 3.705000 ;
      RECT  3.530000  3.190000  3.700000 3.635000 ;
      RECT  3.530000  3.635000  5.270000 3.805000 ;
      RECT  3.880000  2.320000  4.100000 2.490000 ;
      RECT  3.880000  2.490000  4.050000 2.670000 ;
      RECT  3.880000  2.840000  4.050000 3.455000 ;
      RECT  3.930000  0.825000  4.200000 1.325000 ;
      RECT  3.930000  1.325000  4.100000 2.320000 ;
      RECT  4.230000  2.670000  4.450000 3.000000 ;
      RECT  4.280000  1.920000  5.305000 2.150000 ;
      RECT  4.280000  2.150000  4.450000 2.670000 ;
      RECT  4.580000  3.200000  4.910000 3.455000 ;
      RECT  4.630000  2.330000  5.660000 2.500000 ;
      RECT  4.630000  2.500000  4.800000 3.200000 ;
      RECT  4.650000  0.825000  4.980000 1.075000 ;
      RECT  4.650000  1.075000  5.660000 1.245000 ;
      RECT  4.975000  1.425000  5.305000 1.920000 ;
      RECT  4.980000  2.680000  5.310000 2.875000 ;
      RECT  4.980000  2.875000  6.750000 3.000000 ;
      RECT  5.100000  3.000000  6.750000 3.045000 ;
      RECT  5.100000  3.045000  5.270000 3.635000 ;
      RECT  5.450000  3.225000  6.400000 3.705000 ;
      RECT  5.490000  1.245000  5.660000 1.475000 ;
      RECT  5.490000  1.475000  8.110000 1.645000 ;
      RECT  5.490000  1.645000  5.660000 2.330000 ;
      RECT  5.490000  2.500000  5.660000 2.525000 ;
      RECT  5.490000  2.525000  7.260000 2.695000 ;
      RECT  5.840000  1.825000  6.170000 2.175000 ;
      RECT  5.840000  2.175000  8.900000 2.345000 ;
      RECT  6.580000  3.045000  6.750000 3.635000 ;
      RECT  6.580000  3.635000  7.610000 3.805000 ;
      RECT  6.930000  2.695000  7.260000 3.455000 ;
      RECT  7.160000  0.365000  8.110000 0.945000 ;
      RECT  7.440000  3.105000  9.250000 3.275000 ;
      RECT  7.440000  3.275000  7.610000 3.635000 ;
      RECT  7.790000  3.455000  8.740000 3.755000 ;
      RECT  8.570000  2.345000  8.900000 2.925000 ;
      RECT  8.640000  0.615000  8.970000 1.325000 ;
      RECT  8.640000  1.325000  8.900000 2.175000 ;
      RECT  9.080000  1.585000 10.250000 1.755000 ;
      RECT  9.080000  1.755000  9.250000 3.105000 ;
      RECT  9.430000  0.615000 10.600000 0.785000 ;
      RECT  9.430000  0.785000  9.760000 1.325000 ;
      RECT  9.430000  2.675000 10.305000 2.845000 ;
      RECT  9.430000  2.845000  9.680000 3.755000 ;
      RECT  9.625000  1.935000  9.955000 2.435000 ;
      RECT  9.965000  1.085000 10.250000 1.585000 ;
      RECT 10.135000  2.185000 12.495000 2.355000 ;
      RECT 10.135000  2.355000 10.305000 2.675000 ;
      RECT 10.430000  0.785000 10.600000 2.185000 ;
      RECT 10.485000  2.675000 11.435000 3.705000 ;
      RECT 10.805000  1.445000 11.135000 1.835000 ;
      RECT 10.805000  1.835000 12.845000 2.005000 ;
      RECT 11.130000  0.365000 12.080000 0.915000 ;
      RECT 11.840000  2.535000 12.845000 2.705000 ;
      RECT 11.840000  2.705000 12.090000 3.175000 ;
      RECT 12.270000  2.885000 13.165000 3.705000 ;
      RECT 12.620000  0.495000 12.950000 0.995000 ;
      RECT 12.620000  0.995000 12.845000 1.835000 ;
      RECT 12.675000  2.005000 12.845000 2.535000 ;
      RECT 13.225000  0.995000 13.555000 1.495000 ;
      RECT 13.345000  1.495000 13.555000 1.675000 ;
      RECT 13.345000  1.675000 14.720000 2.005000 ;
      RECT 13.345000  2.005000 13.595000 3.005000 ;
      RECT 13.735000  0.365000 14.685000 1.495000 ;
      RECT 13.775000  2.195000 14.720000 3.735000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.985000  0.325000 4.155000 ;
      RECT  0.590000  0.395000  0.760000 0.565000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.985000  0.805000 4.155000 ;
      RECT  0.660000  3.505000  0.830000 3.675000 ;
      RECT  0.950000  0.395000  1.120000 0.565000 ;
      RECT  1.020000  3.505000  1.190000 3.675000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.985000  1.285000 4.155000 ;
      RECT  1.310000  0.395000  1.480000 0.565000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.985000  1.765000 4.155000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  1.950000  2.245000 2.120000 ;
      RECT  2.075000  3.985000  2.245000 4.155000 ;
      RECT  2.230000  0.395000  2.400000 0.565000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.985000  2.725000 4.155000 ;
      RECT  2.590000  0.395000  2.760000 0.565000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.985000  3.205000 4.155000 ;
      RECT  3.050000  3.505000  3.220000 3.675000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.985000  3.685000 4.155000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.985000  4.165000 4.155000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  1.950000  4.645000 2.120000 ;
      RECT  4.475000  3.985000  4.645000 4.155000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.985000  5.125000 4.155000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.985000  5.605000 4.155000 ;
      RECT  5.480000  3.505000  5.650000 3.675000 ;
      RECT  5.840000  3.505000  6.010000 3.675000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.985000  6.085000 4.155000 ;
      RECT  6.200000  3.505000  6.370000 3.675000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.985000  6.565000 4.155000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.985000  7.045000 4.155000 ;
      RECT  7.190000  0.395000  7.360000 0.565000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.985000  7.525000 4.155000 ;
      RECT  7.550000  0.395000  7.720000 0.565000 ;
      RECT  7.820000  3.505000  7.990000 3.675000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.985000  8.005000 4.155000 ;
      RECT  7.910000  0.395000  8.080000 0.565000 ;
      RECT  8.180000  3.505000  8.350000 3.675000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.985000  8.485000 4.155000 ;
      RECT  8.540000  3.505000  8.710000 3.675000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.985000  8.965000 4.155000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.985000  9.445000 4.155000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  1.950000  9.925000 2.120000 ;
      RECT  9.755000  3.985000  9.925000 4.155000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.985000 10.405000 4.155000 ;
      RECT 10.515000  3.505000 10.685000 3.675000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.985000 10.885000 4.155000 ;
      RECT 10.875000  3.505000 11.045000 3.675000 ;
      RECT 11.160000  0.395000 11.330000 0.565000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.985000 11.365000 4.155000 ;
      RECT 11.235000  3.505000 11.405000 3.675000 ;
      RECT 11.520000  0.395000 11.690000 0.565000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.985000 11.845000 4.155000 ;
      RECT 11.880000  0.395000 12.050000 0.565000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.985000 12.325000 4.155000 ;
      RECT 12.270000  3.505000 12.440000 3.675000 ;
      RECT 12.630000  3.505000 12.800000 3.675000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.985000 12.805000 4.155000 ;
      RECT 12.990000  3.505000 13.160000 3.675000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.985000 13.285000 4.155000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.985000 13.765000 4.155000 ;
      RECT 13.765000  0.395000 13.935000 0.565000 ;
      RECT 13.800000  3.505000 13.970000 3.675000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.985000 14.245000 4.155000 ;
      RECT 14.125000  0.395000 14.295000 0.565000 ;
      RECT 14.160000  3.505000 14.330000 3.675000 ;
      RECT 14.485000  0.395000 14.655000 0.565000 ;
      RECT 14.520000  3.505000 14.690000 3.675000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.985000 14.725000 4.155000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.985000 15.205000 4.155000 ;
    LAYER met1 ;
      RECT 2.015000 1.920000 2.305000 1.965000 ;
      RECT 2.015000 1.965000 9.985000 2.105000 ;
      RECT 2.015000 2.105000 2.305000 2.150000 ;
      RECT 4.415000 1.920000 4.705000 1.965000 ;
      RECT 4.415000 2.105000 4.705000 2.150000 ;
      RECT 9.695000 1.920000 9.985000 1.965000 ;
      RECT 9.695000 2.105000 9.985000 2.150000 ;
  END
END sky130_fd_sc_hvl__dfrtp_1
MACRO sky130_fd_sc_hvl__mux4_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__mux4_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.48000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A0
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.770000 1.550000 7.100000 2.520000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.400000 2.300000 4.730000 3.260000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.525000 1.515000 2.150000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 2.300000 3.845000 2.915000 ;
    END
  END A3
  PIN S0
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.565000 2.330000 2.155000 2.500000 ;
        RECT 0.565000 2.500000 0.895000 2.915000 ;
        RECT 1.905000 2.305000 2.155000 2.330000 ;
        RECT 1.905000 2.500000 2.155000 3.635000 ;
        RECT 1.905000 3.635000 3.060000 3.805000 ;
        RECT 2.685000 1.445000 5.420000 1.770000 ;
        RECT 2.685000 1.770000 2.855000 2.800000 ;
        RECT 2.685000 2.800000 3.060000 2.970000 ;
        RECT 2.890000 2.970000 3.060000 3.635000 ;
        RECT 4.925000 0.810000 5.420000 1.445000 ;
    END
  END S0
  PIN S1
    ANTENNAGATEAREA  0.840000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.810000 1.920000 8.220000 2.885000 ;
        RECT 7.810000 2.885000 9.290000 2.915000 ;
        RECT 8.050000 2.915000 9.290000 3.055000 ;
        RECT 9.120000 1.315000 9.370000 1.985000 ;
        RECT 9.120000 1.985000 9.290000 2.885000 ;
    END
  END S1
  PIN X
    ANTENNADIFFAREA  0.596250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.120000 0.605000 12.370000 3.735000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 12.480000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 12.480000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 12.480000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 12.480000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 12.810000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 12.480000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.480000 0.085000 ;
      RECT  0.000000  3.985000 12.480000 4.155000 ;
      RECT  0.110000  0.515000  0.440000 1.175000 ;
      RECT  0.110000  1.175000  2.155000 1.345000 ;
      RECT  0.110000  1.345000  0.280000 3.115000 ;
      RECT  0.110000  3.115000  0.440000 3.575000 ;
      RECT  0.620000  0.365000  1.570000 0.995000 ;
      RECT  0.620000  3.095000  1.570000 3.705000 ;
      RECT  1.905000  1.345000  2.155000 2.035000 ;
      RECT  2.335000  0.495000  2.710000 1.095000 ;
      RECT  2.335000  1.095000  4.550000 1.265000 ;
      RECT  2.335000  1.265000  2.505000 3.175000 ;
      RECT  2.335000  3.175000  2.710000 3.455000 ;
      RECT  3.035000  1.950000  6.240000 2.120000 ;
      RECT  3.035000  2.120000  3.285000 2.620000 ;
      RECT  3.250000  0.365000  4.200000 0.915000 ;
      RECT  3.270000  3.095000  4.220000 3.705000 ;
      RECT  4.380000  0.265000  6.940000 0.435000 ;
      RECT  4.380000  0.435000  4.550000 1.095000 ;
      RECT  5.005000  2.120000  5.335000 2.915000 ;
      RECT  5.460000  3.095000  5.790000 3.595000 ;
      RECT  5.600000  0.615000  6.590000 0.915000 ;
      RECT  5.620000  2.745000  7.630000 2.915000 ;
      RECT  5.620000  2.915000  5.790000 3.095000 ;
      RECT  5.910000  1.095000  6.240000 1.950000 ;
      RECT  6.330000  3.095000  7.280000 3.705000 ;
      RECT  6.420000  0.915000  6.590000 2.745000 ;
      RECT  6.770000  0.435000  6.940000 1.175000 ;
      RECT  6.770000  1.175000  8.000000 1.345000 ;
      RECT  7.120000  0.365000  7.650000 0.995000 ;
      RECT  7.460000  1.570000  8.350000 1.740000 ;
      RECT  7.460000  1.740000  7.630000 2.745000 ;
      RECT  7.460000  2.915000  7.630000 3.115000 ;
      RECT  7.460000  3.115000  7.870000 3.535000 ;
      RECT  7.830000  0.265000  8.700000 0.435000 ;
      RECT  7.830000  0.435000  8.000000 1.175000 ;
      RECT  8.180000  0.615000  8.350000 1.570000 ;
      RECT  8.320000  3.235000  8.650000 3.635000 ;
      RECT  8.320000  3.635000 10.870000 3.805000 ;
      RECT  8.530000  0.435000  8.700000 0.965000 ;
      RECT  8.530000  0.965000  9.990000 1.035000 ;
      RECT  8.530000  1.035000  9.720000 1.135000 ;
      RECT  8.880000  0.265000 10.870000 0.435000 ;
      RECT  8.880000  0.435000  9.210000 0.785000 ;
      RECT  9.470000  3.115000  9.800000 3.455000 ;
      RECT  9.550000  0.615000  9.990000 0.965000 ;
      RECT  9.550000  1.135000  9.720000 3.115000 ;
      RECT  9.900000  2.115000 10.520000 2.655000 ;
      RECT  9.900000  2.655000 10.150000 2.915000 ;
      RECT 10.270000  0.915000 10.520000 2.115000 ;
      RECT 10.700000  0.435000 10.870000 1.595000 ;
      RECT 10.700000  1.595000 11.915000 1.925000 ;
      RECT 10.700000  1.925000 10.870000 3.635000 ;
      RECT 11.050000  0.365000 11.940000 1.415000 ;
      RECT 11.050000  2.175000 11.940000 3.755000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.985000  0.325000 4.155000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.985000  0.805000 4.155000 ;
      RECT  0.650000  0.395000  0.820000 0.565000 ;
      RECT  0.650000  3.505000  0.820000 3.675000 ;
      RECT  1.010000  0.395000  1.180000 0.565000 ;
      RECT  1.010000  3.505000  1.180000 3.675000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.985000  1.285000 4.155000 ;
      RECT  1.370000  0.395000  1.540000 0.565000 ;
      RECT  1.370000  3.505000  1.540000 3.675000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.985000  1.765000 4.155000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.985000  2.245000 4.155000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.985000  2.725000 4.155000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.985000  3.205000 4.155000 ;
      RECT  3.280000  0.395000  3.450000 0.565000 ;
      RECT  3.300000  3.505000  3.470000 3.675000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.985000  3.685000 4.155000 ;
      RECT  3.640000  0.395000  3.810000 0.565000 ;
      RECT  3.660000  3.505000  3.830000 3.675000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.985000  4.165000 4.155000 ;
      RECT  4.000000  0.395000  4.170000 0.565000 ;
      RECT  4.020000  3.505000  4.190000 3.675000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.985000  4.645000 4.155000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.985000  5.125000 4.155000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.985000  5.605000 4.155000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.985000  6.085000 4.155000 ;
      RECT  6.360000  3.505000  6.530000 3.675000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.985000  6.565000 4.155000 ;
      RECT  6.720000  3.505000  6.890000 3.675000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.985000  7.045000 4.155000 ;
      RECT  7.080000  3.505000  7.250000 3.675000 ;
      RECT  7.120000  0.395000  7.290000 0.565000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.985000  7.525000 4.155000 ;
      RECT  7.480000  0.395000  7.650000 0.565000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.985000  8.005000 4.155000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.985000  8.485000 4.155000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.985000  8.965000 4.155000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.985000  9.445000 4.155000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.985000  9.925000 4.155000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.985000 10.405000 4.155000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.985000 10.885000 4.155000 ;
      RECT 11.050000  0.395000 11.220000 0.565000 ;
      RECT 11.050000  3.505000 11.220000 3.675000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.985000 11.365000 4.155000 ;
      RECT 11.410000  0.395000 11.580000 0.565000 ;
      RECT 11.410000  3.505000 11.580000 3.675000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.985000 11.845000 4.155000 ;
      RECT 11.770000  0.395000 11.940000 0.565000 ;
      RECT 11.770000  3.505000 11.940000 3.675000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.985000 12.325000 4.155000 ;
  END
END sky130_fd_sc_hvl__mux4_1
MACRO sky130_fd_sc_hvl__a22o_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__a22o_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A1
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.505000 4.645000 1.750000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.825000 1.505000 5.155000 1.750000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.035000 0.810000 3.205000 1.750000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.990000 1.775000 2.320000 3.260000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.626250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.495000 0.380000 3.755000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 5.280000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 5.280000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 5.280000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 5.280000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 5.610000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 5.280000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.280000 0.085000 ;
      RECT 0.000000  3.985000 5.280000 4.155000 ;
      RECT 0.550000  0.365000 2.260000 1.245000 ;
      RECT 0.560000  2.175000 1.460000 3.755000 ;
      RECT 0.585000  1.425000 2.855000 1.595000 ;
      RECT 0.585000  1.595000 0.915000 1.755000 ;
      RECT 1.640000  2.175000 1.810000 3.635000 ;
      RECT 1.640000  3.635000 3.530000 3.805000 ;
      RECT 2.500000  1.595000 2.830000 3.455000 ;
      RECT 2.685000  0.460000 3.635000 0.630000 ;
      RECT 2.685000  0.630000 2.855000 1.425000 ;
      RECT 3.280000  1.930000 5.170000 2.100000 ;
      RECT 3.280000  2.100000 3.530000 3.635000 ;
      RECT 3.385000  0.630000 3.635000 1.325000 ;
      RECT 3.710000  2.280000 4.660000 3.755000 ;
      RECT 3.815000  0.365000 5.125000 1.325000 ;
      RECT 4.840000  2.100000 5.170000 3.735000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.565000  3.505000 0.735000 3.675000 ;
      RECT 0.600000  0.395000 0.770000 0.565000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.925000  3.505000 1.095000 3.675000 ;
      RECT 0.960000  0.395000 1.130000 0.565000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.285000  3.505000 1.455000 3.675000 ;
      RECT 1.320000  0.395000 1.490000 0.565000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.680000  0.395000 1.850000 0.565000 ;
      RECT 2.040000  0.395000 2.210000 0.565000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.985000 3.685000 4.155000 ;
      RECT 3.740000  3.505000 3.910000 3.675000 ;
      RECT 3.845000  0.395000 4.015000 0.565000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.985000 4.165000 4.155000 ;
      RECT 4.100000  3.505000 4.270000 3.675000 ;
      RECT 4.205000  0.395000 4.375000 0.565000 ;
      RECT 4.460000  3.505000 4.630000 3.675000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.985000 4.645000 4.155000 ;
      RECT 4.565000  0.395000 4.735000 0.565000 ;
      RECT 4.925000  0.395000 5.095000 0.565000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.985000 5.125000 4.155000 ;
  END
END sky130_fd_sc_hvl__a22o_1
MACRO sky130_fd_sc_hvl__or2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__or2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.530000 1.175000 1.860000 1.725000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.175000 0.935000 1.725000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.641250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.980000 0.495000 3.235000 3.755000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 3.360000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 3.360000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 3.360000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 3.360000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 3.690000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 3.360000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.985000 3.360000 4.155000 ;
      RECT 0.090000  0.365000 1.000000 0.995000 ;
      RECT 0.400000  1.905000 2.775000 2.075000 ;
      RECT 0.400000  2.075000 0.650000 2.675000 ;
      RECT 0.830000  2.255000 2.800000 3.755000 ;
      RECT 1.180000  0.495000 1.510000 0.995000 ;
      RECT 1.180000  0.995000 1.350000 1.905000 ;
      RECT 2.040000  0.365000 2.630000 1.325000 ;
      RECT 2.445000  1.725000 2.775000 1.905000 ;
    LAYER mcon ;
      RECT 0.100000  0.395000 0.270000 0.565000 ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.460000  0.395000 0.630000 0.565000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.820000  0.395000 0.990000 0.565000 ;
      RECT 0.830000  3.505000 1.000000 3.675000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.190000  3.505000 1.360000 3.675000 ;
      RECT 1.550000  3.505000 1.720000 3.675000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.910000  3.505000 2.080000 3.675000 ;
      RECT 2.070000  0.395000 2.240000 0.565000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.270000  3.505000 2.440000 3.675000 ;
      RECT 2.430000  0.395000 2.600000 0.565000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 2.630000  3.505000 2.800000 3.675000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
  END
END sky130_fd_sc_hvl__or2_1
MACRO sky130_fd_sc_hvl__o21a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__o21a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A1
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.505000 4.195000 1.835000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.555000 1.550000 2.785000 3.260000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.805000 2.000000 2.120000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.626250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.525000 0.380000 1.975000 ;
        RECT 0.125000 1.975000 0.595000 3.755000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 4.320000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 4.320000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 4.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 4.320000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 4.650000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 4.320000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.985000 4.320000 4.155000 ;
      RECT 0.550000  0.365000 1.315000 1.275000 ;
      RECT 0.550000  1.455000 2.375000 1.625000 ;
      RECT 0.550000  1.625000 0.835000 1.795000 ;
      RECT 0.775000  2.300000 2.025000 3.755000 ;
      RECT 1.495000  0.495000 1.825000 1.455000 ;
      RECT 2.205000  1.625000 2.375000 3.755000 ;
      RECT 2.275000  0.495000 2.605000 1.105000 ;
      RECT 2.275000  1.105000 4.185000 1.275000 ;
      RECT 2.785000  0.365000 3.675000 0.925000 ;
      RECT 2.965000  2.175000 4.230000 3.755000 ;
      RECT 3.855000  0.495000 4.185000 1.105000 ;
      RECT 3.855000  1.275000 4.185000 1.325000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.600000  0.395000 0.770000 0.565000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.775000  3.505000 0.945000 3.675000 ;
      RECT 1.105000  0.395000 1.275000 0.565000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.135000  3.505000 1.305000 3.675000 ;
      RECT 1.495000  3.505000 1.665000 3.675000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.855000  3.505000 2.025000 3.675000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 2.785000  0.395000 2.955000 0.565000 ;
      RECT 2.970000  3.505000 3.140000 3.675000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
      RECT 3.145000  0.395000 3.315000 0.565000 ;
      RECT 3.330000  3.505000 3.500000 3.675000 ;
      RECT 3.505000  0.395000 3.675000 0.565000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.985000 3.685000 4.155000 ;
      RECT 3.690000  3.505000 3.860000 3.675000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.985000 4.165000 4.155000 ;
      RECT 4.050000  3.505000 4.220000 3.675000 ;
  END
END sky130_fd_sc_hvl__o21a_1
MACRO sky130_fd_sc_hvl__sdfxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__sdfxtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.88000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN D
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 2.205000 2.755000 2.520000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.596250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.660000 0.615000 14.020000 1.505000 ;
        RECT 13.660000 2.195000 14.020000 3.735000 ;
        RECT 13.850000 1.505000 14.755000 1.780000 ;
        RECT 13.850000 1.780000 14.020000 2.195000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.600000 2.215000 4.195000 2.765000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.840000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.445000 1.795000 1.855000 ;
        RECT 0.605000 1.855000 3.050000 2.025000 ;
        RECT 2.720000 1.095000 3.050000 1.855000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.345000 1.175000 4.675000 1.685000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 14.880000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 14.880000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 14.880000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 14.880000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 15.210000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 14.880000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 14.880000 0.085000 ;
      RECT  0.000000  3.985000 14.880000 4.155000 ;
      RECT  0.125000  0.515000  0.455000 1.095000 ;
      RECT  0.125000  1.095000  2.305000 1.265000 ;
      RECT  0.125000  1.265000  0.380000 3.425000 ;
      RECT  0.905000  0.365000  1.855000 0.915000 ;
      RECT  0.910000  2.925000  1.860000 3.705000 ;
      RECT  1.975000  1.265000  2.305000 1.675000 ;
      RECT  2.395000  0.495000  2.725000 0.745000 ;
      RECT  2.395000  0.745000  3.400000 0.915000 ;
      RECT  2.400000  2.925000  3.400000 3.095000 ;
      RECT  2.400000  3.095000  2.730000 3.425000 ;
      RECT  3.230000  0.915000  3.400000 1.865000 ;
      RECT  3.230000  1.865000  6.780000 2.035000 ;
      RECT  3.230000  2.035000  3.400000 2.925000 ;
      RECT  3.580000  0.365000  4.485000 0.995000 ;
      RECT  3.635000  2.945000  4.585000 3.735000 ;
      RECT  4.665000  0.515000  5.025000 0.975000 ;
      RECT  4.765000  2.595000  5.605000 2.765000 ;
      RECT  4.765000  2.765000  5.095000 3.735000 ;
      RECT  4.855000  0.975000  5.025000 1.155000 ;
      RECT  4.855000  1.155000  5.870000 1.325000 ;
      RECT  5.215000  0.365000  5.805000 0.975000 ;
      RECT  5.275000  2.215000  5.605000 2.595000 ;
      RECT  5.315000  2.945000  5.905000 3.735000 ;
      RECT  5.540000  1.325000  5.870000 1.685000 ;
      RECT  5.995000  0.265000  8.210000 0.435000 ;
      RECT  5.995000  0.435000  6.325000 0.975000 ;
      RECT  6.095000  2.945000  6.425000 3.335000 ;
      RECT  6.095000  3.335000  7.325000 3.505000 ;
      RECT  6.095000  3.505000  6.425000 3.735000 ;
      RECT  6.565000  0.615000  6.895000 0.995000 ;
      RECT  6.565000  0.995000  6.780000 1.865000 ;
      RECT  6.610000  2.035000  6.780000 2.695000 ;
      RECT  6.610000  2.695000  6.975000 3.155000 ;
      RECT  6.960000  2.225000  7.325000 2.515000 ;
      RECT  7.075000  0.435000  7.245000 2.225000 ;
      RECT  7.155000  2.515000  7.325000 3.335000 ;
      RECT  7.425000  0.615000  7.755000 0.995000 ;
      RECT  7.505000  0.995000  7.755000 1.605000 ;
      RECT  7.505000  1.605000  9.685000 1.775000 ;
      RECT  7.505000  1.775000  7.675000 2.675000 ;
      RECT  7.505000  2.675000  7.755000 3.175000 ;
      RECT  7.880000  1.955000  8.210000 2.495000 ;
      RECT  7.935000  0.435000  8.210000 1.255000 ;
      RECT  7.935000  1.255000 10.295000 1.425000 ;
      RECT  8.040000  2.495000  8.210000 3.155000 ;
      RECT  8.040000  3.155000 10.490000 3.325000 ;
      RECT  8.620000  1.955000 10.645000 2.125000 ;
      RECT  8.620000  2.125000  8.950000 2.555000 ;
      RECT  8.680000  0.365000  9.630000 1.075000 ;
      RECT  9.030000  3.505000  9.980000 3.755000 ;
      RECT  9.810000  0.495000 10.140000 0.905000 ;
      RECT  9.810000  0.905000 10.645000 1.075000 ;
      RECT  9.810000  2.125000  9.980000 2.675000 ;
      RECT  9.810000  2.675000 10.140000 2.975000 ;
      RECT 10.045000  1.425000 10.295000 1.775000 ;
      RECT 10.160000  2.305000 10.490000 2.495000 ;
      RECT 10.320000  2.495000 10.490000 3.155000 ;
      RECT 10.320000  3.325000 11.450000 3.495000 ;
      RECT 10.475000  1.075000 10.645000 1.955000 ;
      RECT 10.670000  2.675000 11.075000 3.145000 ;
      RECT 10.825000  0.495000 11.800000 0.665000 ;
      RECT 10.825000  0.665000 11.075000 2.675000 ;
      RECT 11.255000  1.085000 11.450000 3.325000 ;
      RECT 11.630000  0.665000 11.800000 2.345000 ;
      RECT 11.630000  2.345000 12.930000 2.515000 ;
      RECT 11.980000  0.365000 12.930000 1.305000 ;
      RECT 11.980000  1.485000 13.440000 1.655000 ;
      RECT 11.980000  1.655000 12.310000 2.155000 ;
      RECT 11.980000  2.695000 12.930000 3.735000 ;
      RECT 12.600000  1.845000 12.930000 2.345000 ;
      RECT 13.110000  0.515000 13.440000 1.485000 ;
      RECT 13.110000  1.655000 13.440000 1.685000 ;
      RECT 13.110000  1.685000 13.670000 2.015000 ;
      RECT 13.110000  2.015000 13.440000 3.735000 ;
      RECT 14.200000  0.365000 14.790000 1.325000 ;
      RECT 14.200000  2.195000 14.790000 3.735000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.985000  0.325000 4.155000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.985000  0.805000 4.155000 ;
      RECT  0.935000  0.395000  1.105000 0.565000 ;
      RECT  0.940000  3.505000  1.110000 3.675000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.985000  1.285000 4.155000 ;
      RECT  1.295000  0.395000  1.465000 0.565000 ;
      RECT  1.300000  3.505000  1.470000 3.675000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.985000  1.765000 4.155000 ;
      RECT  1.655000  0.395000  1.825000 0.565000 ;
      RECT  1.660000  3.505000  1.830000 3.675000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.985000  2.245000 4.155000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.985000  2.725000 4.155000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.985000  3.205000 4.155000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.985000  3.685000 4.155000 ;
      RECT  3.590000  0.395000  3.760000 0.565000 ;
      RECT  3.665000  3.505000  3.835000 3.675000 ;
      RECT  3.950000  0.395000  4.120000 0.565000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.985000  4.165000 4.155000 ;
      RECT  4.025000  3.505000  4.195000 3.675000 ;
      RECT  4.310000  0.395000  4.480000 0.565000 ;
      RECT  4.385000  3.505000  4.555000 3.675000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.985000  4.645000 4.155000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.985000  5.125000 4.155000 ;
      RECT  5.245000  0.395000  5.415000 0.565000 ;
      RECT  5.345000  3.505000  5.515000 3.675000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.985000  5.605000 4.155000 ;
      RECT  5.605000  0.395000  5.775000 0.565000 ;
      RECT  5.705000  3.505000  5.875000 3.675000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.985000  6.085000 4.155000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.985000  6.565000 4.155000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.985000  7.045000 4.155000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.985000  7.525000 4.155000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.985000  8.005000 4.155000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.985000  8.485000 4.155000 ;
      RECT  8.710000  0.395000  8.880000 0.565000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.985000  8.965000 4.155000 ;
      RECT  9.060000  3.535000  9.230000 3.705000 ;
      RECT  9.070000  0.395000  9.240000 0.565000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.985000  9.445000 4.155000 ;
      RECT  9.420000  3.535000  9.590000 3.705000 ;
      RECT  9.430000  0.395000  9.600000 0.565000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.985000  9.925000 4.155000 ;
      RECT  9.780000  3.535000  9.950000 3.705000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.985000 10.405000 4.155000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.985000 10.885000 4.155000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.985000 11.365000 4.155000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.985000 11.845000 4.155000 ;
      RECT 12.010000  0.395000 12.180000 0.565000 ;
      RECT 12.010000  3.505000 12.180000 3.675000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.985000 12.325000 4.155000 ;
      RECT 12.370000  0.395000 12.540000 0.565000 ;
      RECT 12.370000  3.505000 12.540000 3.675000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.985000 12.805000 4.155000 ;
      RECT 12.730000  0.395000 12.900000 0.565000 ;
      RECT 12.730000  3.505000 12.900000 3.675000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.985000 13.285000 4.155000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.985000 13.765000 4.155000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.985000 14.245000 4.155000 ;
      RECT 14.230000  0.395000 14.400000 0.565000 ;
      RECT 14.230000  3.505000 14.400000 3.675000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.985000 14.725000 4.155000 ;
      RECT 14.590000  0.395000 14.760000 0.565000 ;
      RECT 14.590000  3.505000 14.760000 3.675000 ;
  END
END sky130_fd_sc_hvl__sdfxtp_1
MACRO sky130_fd_sc_hvl__nor3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__nor3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.525000 0.425000 2.120000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.775000 1.795000 2.120000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.975000 1.775000 2.305000 3.260000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  0.836250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.930000 0.495000 1.180000 1.425000 ;
        RECT 0.930000 1.425000 2.755000 1.595000 ;
        RECT 2.490000 0.495000 2.755000 1.425000 ;
        RECT 2.490000 1.595000 2.755000 3.755000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 3.360000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 3.360000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 3.360000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 3.360000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 3.690000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 3.360000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.985000 3.360000 4.155000 ;
      RECT 0.090000  0.365000 0.680000 1.325000 ;
      RECT 0.090000  2.300000 1.760000 3.755000 ;
      RECT 1.360000  0.365000 2.310000 1.245000 ;
    LAYER mcon ;
      RECT 0.120000  0.395000 0.290000 0.565000 ;
      RECT 0.120000  3.505000 0.290000 3.675000 ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.480000  0.395000 0.650000 0.565000 ;
      RECT 0.480000  3.505000 0.650000 3.675000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.840000  3.505000 1.010000 3.675000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.200000  3.505000 1.370000 3.675000 ;
      RECT 1.390000  0.395000 1.560000 0.565000 ;
      RECT 1.560000  3.505000 1.730000 3.675000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.750000  0.395000 1.920000 0.565000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.110000  0.395000 2.280000 0.565000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
  END
END sky130_fd_sc_hvl__nor3_1
MACRO sky130_fd_sc_hvl__dfxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__dfxtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.00000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN D
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.595000 1.555000 2.470000 1.750000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.596250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.560000 2.185000 11.890000 3.735000 ;
        RECT 11.640000 0.685000 11.890000 2.185000 ;
    END
  END Q
  PIN CLK
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.540000 1.905000 0.870000 2.575000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 12.000000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 12.000000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 12.000000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 12.000000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 12.330000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 12.000000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.000000 0.085000 ;
      RECT  0.000000  3.985000 12.000000 4.155000 ;
      RECT  0.110000  0.595000  0.380000 1.555000 ;
      RECT  0.110000  1.555000  1.415000 1.725000 ;
      RECT  0.110000  1.725000  0.360000 3.565000 ;
      RECT  0.540000  2.755000  1.490000 3.705000 ;
      RECT  0.560000  0.365000  1.510000 1.095000 ;
      RECT  1.165000  1.725000  1.415000 1.930000 ;
      RECT  1.165000  1.930000  2.820000 2.225000 ;
      RECT  1.670000  2.445000  2.820000 2.615000 ;
      RECT  1.670000  2.615000  2.000000 3.565000 ;
      RECT  1.690000  0.595000  2.020000 1.205000 ;
      RECT  1.690000  1.205000  3.115000 1.375000 ;
      RECT  2.200000  0.365000  2.765000 1.025000 ;
      RECT  2.220000  2.795000  2.470000 3.705000 ;
      RECT  2.650000  1.760000  3.685000 1.930000 ;
      RECT  2.650000  2.615000  2.820000 3.305000 ;
      RECT  2.650000  3.305000  3.680000 3.475000 ;
      RECT  2.945000  0.265000  5.055000 0.435000 ;
      RECT  2.945000  0.435000  3.115000 1.205000 ;
      RECT  3.000000  2.110000  4.035000 2.280000 ;
      RECT  3.000000  2.280000  3.330000 3.125000 ;
      RECT  3.295000  0.615000  4.035000 1.025000 ;
      RECT  3.430000  1.205000  3.685000 1.760000 ;
      RECT  3.510000  2.460000  3.840000 3.135000 ;
      RECT  3.510000  3.135000  7.655000 3.305000 ;
      RECT  3.865000  1.025000  4.035000 2.110000 ;
      RECT  4.055000  2.675000  4.385000 2.955000 ;
      RECT  4.215000  0.615000  4.545000 1.525000 ;
      RECT  4.215000  1.525000  6.345000 1.695000 ;
      RECT  4.215000  1.695000  4.385000 2.675000 ;
      RECT  4.565000  1.885000  4.890000 2.385000 ;
      RECT  4.565000  2.385000  6.955000 2.555000 ;
      RECT  4.725000  0.435000  5.055000 1.175000 ;
      RECT  4.725000  1.175000  6.555000 1.345000 ;
      RECT  5.070000  3.485000  6.020000 3.735000 ;
      RECT  5.255000  0.365000  6.205000 0.995000 ;
      RECT  5.435000  1.875000  7.305000 2.045000 ;
      RECT  5.435000  2.045000  5.765000 2.205000 ;
      RECT  6.385000  0.265000  7.450000 0.435000 ;
      RECT  6.385000  0.435000  6.555000 1.175000 ;
      RECT  6.470000  2.755000  7.305000 2.955000 ;
      RECT  6.705000  2.225000  6.955000 2.385000 ;
      RECT  6.735000  0.615000  7.065000 1.875000 ;
      RECT  7.135000  2.045000  7.305000 2.755000 ;
      RECT  7.280000  0.435000  7.450000 1.125000 ;
      RECT  7.280000  1.125000  7.655000 1.445000 ;
      RECT  7.485000  1.445000  7.655000 2.225000 ;
      RECT  7.485000  2.225000  8.250000 2.515000 ;
      RECT  7.485000  2.515000  7.655000 3.135000 ;
      RECT  7.630000  0.525000  8.005000 0.855000 ;
      RECT  7.630000  0.855000  8.600000 0.945000 ;
      RECT  7.835000  0.945000  8.600000 1.025000 ;
      RECT  7.835000  2.695000  8.600000 2.865000 ;
      RECT  7.835000  2.865000  8.085000 3.735000 ;
      RECT  8.430000  1.025000  8.600000 2.275000 ;
      RECT  8.430000  2.275000 10.035000 2.445000 ;
      RECT  8.430000  2.445000  8.600000 2.695000 ;
      RECT  8.780000  0.365000  9.730000 1.245000 ;
      RECT  8.815000  2.695000  9.765000 3.735000 ;
      RECT  9.000000  1.425000 10.510000 1.595000 ;
      RECT  9.000000  1.595000  9.330000 2.015000 ;
      RECT  9.705000  1.775000 10.035000 2.275000 ;
      RECT 10.180000  0.525000 10.510000 1.425000 ;
      RECT 10.215000  1.595000 10.510000 1.675000 ;
      RECT 10.215000  1.675000 11.460000 2.005000 ;
      RECT 10.215000  2.005000 10.545000 3.735000 ;
      RECT 10.690000  0.365000 11.280000 1.495000 ;
      RECT 10.725000  2.195000 11.315000 3.735000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.985000  0.325000 4.155000 ;
      RECT  0.570000  3.505000  0.740000 3.675000 ;
      RECT  0.590000  0.395000  0.760000 0.565000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.985000  0.805000 4.155000 ;
      RECT  0.930000  3.505000  1.100000 3.675000 ;
      RECT  0.950000  0.395000  1.120000 0.565000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.985000  1.285000 4.155000 ;
      RECT  1.290000  3.505000  1.460000 3.675000 ;
      RECT  1.310000  0.395000  1.480000 0.565000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.985000  1.765000 4.155000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.985000  2.245000 4.155000 ;
      RECT  2.215000  0.395000  2.385000 0.565000 ;
      RECT  2.250000  3.505000  2.420000 3.675000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.985000  2.725000 4.155000 ;
      RECT  2.575000  0.395000  2.745000 0.565000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.985000  3.205000 4.155000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.985000  3.685000 4.155000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.985000  4.165000 4.155000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.985000  4.645000 4.155000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.985000  5.125000 4.155000 ;
      RECT  5.100000  3.515000  5.270000 3.685000 ;
      RECT  5.285000  0.395000  5.455000 0.565000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.985000  5.605000 4.155000 ;
      RECT  5.460000  3.515000  5.630000 3.685000 ;
      RECT  5.645000  0.395000  5.815000 0.565000 ;
      RECT  5.820000  3.515000  5.990000 3.685000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.985000  6.085000 4.155000 ;
      RECT  6.005000  0.395000  6.175000 0.565000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.985000  6.565000 4.155000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.985000  7.045000 4.155000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.985000  7.525000 4.155000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.985000  8.005000 4.155000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.985000  8.485000 4.155000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.985000  8.965000 4.155000 ;
      RECT  8.810000  0.395000  8.980000 0.565000 ;
      RECT  8.845000  3.505000  9.015000 3.675000 ;
      RECT  9.170000  0.395000  9.340000 0.565000 ;
      RECT  9.205000  3.505000  9.375000 3.675000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.985000  9.445000 4.155000 ;
      RECT  9.530000  0.395000  9.700000 0.565000 ;
      RECT  9.565000  3.505000  9.735000 3.675000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.985000  9.925000 4.155000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.985000 10.405000 4.155000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.985000 10.885000 4.155000 ;
      RECT 10.720000  0.395000 10.890000 0.565000 ;
      RECT 10.755000  3.505000 10.925000 3.675000 ;
      RECT 11.080000  0.395000 11.250000 0.565000 ;
      RECT 11.115000  3.505000 11.285000 3.675000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.985000 11.365000 4.155000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.985000 11.845000 4.155000 ;
  END
END sky130_fd_sc_hvl__dfxtp_1
MACRO sky130_fd_sc_hvl__einvp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__einvp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.275000 1.625000 2.865000 1.955000 ;
        RECT 2.445000 1.160000 2.810000 1.625000 ;
        RECT 2.445000 1.955000 2.810000 2.540000 ;
    END
  END A
  PIN TE
    ANTENNAGATEAREA  0.960000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.505000 1.305000 1.750000 ;
    END
  END TE
  PIN Z
    ANTENNADIFFAREA  0.641250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.980000 0.575000 3.235000 1.455000 ;
        RECT 2.980000 2.125000 3.235000 3.755000 ;
        RECT 3.035000 1.455000 3.235000 2.125000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 3.360000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 3.360000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 3.360000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 3.360000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 3.690000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 3.360000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.985000 3.360000 4.155000 ;
      RECT 0.175000  0.905000 0.380000 1.335000 ;
      RECT 0.175000  1.335000 0.345000 1.930000 ;
      RECT 0.175000  1.930000 2.065000 2.100000 ;
      RECT 0.175000  2.100000 0.650000 3.005000 ;
      RECT 0.470000  0.365000 2.800000 0.735000 ;
      RECT 0.550000  0.735000 2.800000 0.990000 ;
      RECT 0.550000  0.990000 2.275000 1.335000 ;
      RECT 0.830000  2.280000 2.275000 2.710000 ;
      RECT 0.830000  2.710000 2.800000 3.755000 ;
      RECT 1.475000  1.725000 2.065000 1.930000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.470000  0.395000 0.640000 0.565000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.830000  0.395000 1.000000 0.565000 ;
      RECT 0.830000  3.505000 1.000000 3.675000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.190000  0.395000 1.360000 0.565000 ;
      RECT 1.190000  3.505000 1.360000 3.675000 ;
      RECT 1.550000  0.395000 1.720000 0.565000 ;
      RECT 1.550000  3.505000 1.720000 3.675000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.910000  0.395000 2.080000 0.565000 ;
      RECT 1.910000  3.505000 2.080000 3.675000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.270000  0.395000 2.440000 0.565000 ;
      RECT 2.270000  3.505000 2.440000 3.675000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 2.630000  0.395000 2.800000 0.565000 ;
      RECT 2.630000  3.505000 2.800000 3.675000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
  END
END sky130_fd_sc_hvl__einvp_1
MACRO sky130_fd_sc_hvl__and2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__and2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.175000 0.535000 1.845000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 0.810000 1.455000 1.725000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.626250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.980000 0.495000 3.255000 3.755000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 3.360000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 3.360000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 3.360000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 3.360000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 3.690000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 3.360000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.985000 3.360000 4.155000 ;
      RECT 0.090000  2.255000 1.020000 3.705000 ;
      RECT 0.130000  0.495000 0.380000 0.825000 ;
      RECT 0.130000  0.825000 0.885000 0.995000 ;
      RECT 0.715000  0.995000 0.885000 1.905000 ;
      RECT 0.715000  1.905000 2.775000 2.075000 ;
      RECT 1.200000  2.075000 1.370000 2.675000 ;
      RECT 1.550000  2.255000 2.800000 3.755000 ;
      RECT 1.635000  0.365000 2.625000 1.325000 ;
      RECT 2.445000  1.725000 2.775000 1.905000 ;
    LAYER mcon ;
      RECT 0.110000  3.505000 0.280000 3.675000 ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.470000  3.505000 0.640000 3.675000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.830000  3.505000 1.000000 3.675000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.550000  3.505000 1.720000 3.675000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.685000  0.395000 1.855000 0.565000 ;
      RECT 1.910000  3.505000 2.080000 3.675000 ;
      RECT 2.045000  0.395000 2.215000 0.565000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.270000  3.505000 2.440000 3.675000 ;
      RECT 2.405000  0.395000 2.575000 0.565000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 2.630000  3.505000 2.800000 3.675000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
  END
END sky130_fd_sc_hvl__and2_1
MACRO sky130_fd_sc_hvl__and3_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__and3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.810000 0.935000 1.645000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 2.175000 1.565000 2.490000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.115000 0.810000 2.255000 1.645000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.626250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.365000 2.175000 3.715000 3.755000 ;
        RECT 3.410000 0.495000 3.715000 2.175000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 3.840000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 3.840000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 3.840000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 3.840000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 4.170000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 3.840000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.985000 3.840000 4.155000 ;
      RECT 0.130000  0.825000 0.425000 1.825000 ;
      RECT 0.130000  1.825000 3.240000 1.995000 ;
      RECT 0.130000  1.995000 0.380000 3.045000 ;
      RECT 0.560000  2.670000 1.510000 3.705000 ;
      RECT 1.770000  1.995000 2.020000 3.045000 ;
      RECT 2.200000  2.175000 3.150000 3.755000 ;
      RECT 2.435000  0.365000 3.240000 1.325000 ;
      RECT 2.910000  1.665000 3.240000 1.825000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.590000  3.505000 0.760000 3.675000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.950000  3.505000 1.120000 3.675000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.310000  3.505000 1.480000 3.675000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.230000  3.505000 2.400000 3.675000 ;
      RECT 2.485000  0.395000 2.655000 0.565000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 2.590000  3.505000 2.760000 3.675000 ;
      RECT 2.950000  3.505000 3.120000 3.675000 ;
      RECT 3.015000  0.395000 3.185000 0.565000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.985000 3.685000 4.155000 ;
  END
END sky130_fd_sc_hvl__and3_1
MACRO sky130_fd_sc_hvl__o22a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__o22a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A1
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.420000 1.775000 2.150000 2.055000 ;
        RECT 1.980000 1.400000 2.775000 1.570000 ;
        RECT 1.980000 1.570000 2.150000 1.775000 ;
        RECT 2.605000 1.230000 4.880000 1.400000 ;
        RECT 3.035000 1.210000 3.710000 1.230000 ;
        RECT 4.550000 1.400000 4.880000 2.015000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.580000 4.195000 1.910000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.330000 1.750000 2.755000 2.120000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.955000 1.580000 3.250000 2.120000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.641250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.495000 0.380000 3.755000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 5.280000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 5.280000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 5.280000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 5.280000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 5.610000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 5.280000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.280000 0.085000 ;
      RECT 0.000000  3.985000 5.280000 4.155000 ;
      RECT 0.560000  0.365000 1.450000 1.245000 ;
      RECT 0.560000  2.650000 3.250000 3.755000 ;
      RECT 0.585000  1.425000 1.800000 1.595000 ;
      RECT 0.585000  1.595000 0.915000 2.300000 ;
      RECT 0.585000  2.300000 3.680000 2.470000 ;
      RECT 1.630000  1.050000 2.425000 1.220000 ;
      RECT 1.630000  1.220000 1.800000 1.425000 ;
      RECT 1.745000  0.265000 3.680000 0.435000 ;
      RECT 1.745000  0.435000 2.075000 0.870000 ;
      RECT 2.255000  0.880000 2.855000 1.050000 ;
      RECT 2.525000  0.615000 2.855000 0.880000 ;
      RECT 3.350000  0.435000 3.680000 1.030000 ;
      RECT 3.430000  2.175000 3.680000 2.300000 ;
      RECT 3.430000  2.470000 3.680000 3.755000 ;
      RECT 3.860000  2.195000 5.170000 3.735000 ;
      RECT 3.890000  0.365000 5.190000 1.050000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.560000  0.395000 0.730000 0.565000 ;
      RECT 0.560000  3.505000 0.730000 3.675000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.920000  0.395000 1.090000 0.565000 ;
      RECT 0.920000  3.505000 1.090000 3.675000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.280000  0.395000 1.450000 0.565000 ;
      RECT 1.280000  3.505000 1.450000 3.675000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.640000  3.505000 1.810000 3.675000 ;
      RECT 2.000000  3.505000 2.170000 3.675000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.360000  3.505000 2.530000 3.675000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 2.720000  3.505000 2.890000 3.675000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
      RECT 3.080000  3.505000 3.250000 3.675000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.985000 3.685000 4.155000 ;
      RECT 3.890000  3.505000 4.060000 3.675000 ;
      RECT 3.915000  0.395000 4.085000 0.565000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.985000 4.165000 4.155000 ;
      RECT 4.250000  3.505000 4.420000 3.675000 ;
      RECT 4.275000  0.395000 4.445000 0.565000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.985000 4.645000 4.155000 ;
      RECT 4.610000  3.505000 4.780000 3.675000 ;
      RECT 4.635000  0.395000 4.805000 0.565000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.985000 5.125000 4.155000 ;
      RECT 4.970000  3.505000 5.140000 3.675000 ;
      RECT 4.995000  0.395000 5.165000 0.565000 ;
  END
END sky130_fd_sc_hvl__o22a_1
MACRO sky130_fd_sc_hvl__einvn_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__einvn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.275000 1.725000 2.780000 2.540000 ;
        RECT 2.505000 1.160000 2.780000 1.725000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  1.335000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.825000 1.795000 2.025000 ;
        RECT 0.635000 2.025000 1.795000 2.120000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.641250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.950000 0.495000 3.235000 3.755000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 3.360000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 3.360000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 3.360000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 3.360000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 3.690000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 3.360000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.985000 3.360000 4.155000 ;
      RECT 0.090000  0.910000 0.440000 1.425000 ;
      RECT 0.090000  1.425000 2.065000 1.645000 ;
      RECT 0.090000  1.645000 0.345000 2.195000 ;
      RECT 0.090000  2.195000 0.455000 2.300000 ;
      RECT 0.090000  2.300000 0.535000 3.025000 ;
      RECT 0.440000  0.365000 2.770000 0.740000 ;
      RECT 0.610000  0.740000 2.770000 0.900000 ;
      RECT 0.610000  0.900000 2.335000 1.245000 ;
      RECT 0.740000  2.300000 2.105000 2.710000 ;
      RECT 0.740000  2.710000 2.770000 3.755000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.440000  0.395000 0.610000 0.565000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.770000  3.505000 0.940000 3.675000 ;
      RECT 0.800000  0.395000 0.970000 0.565000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.130000  3.505000 1.300000 3.675000 ;
      RECT 1.160000  0.395000 1.330000 0.565000 ;
      RECT 1.490000  3.505000 1.660000 3.675000 ;
      RECT 1.520000  0.395000 1.690000 0.565000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.850000  3.505000 2.020000 3.675000 ;
      RECT 1.880000  0.395000 2.050000 0.565000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.210000  3.505000 2.380000 3.675000 ;
      RECT 2.240000  0.395000 2.410000 0.565000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 2.570000  3.505000 2.740000 3.675000 ;
      RECT 2.600000  0.395000 2.770000 0.565000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
  END
END sky130_fd_sc_hvl__einvn_1
MACRO sky130_fd_sc_hvl__diode_2
  CLASS CORE ANTENNACELL ;
  FOREIGN sky130_fd_sc_hvl__diode_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  0.960000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN DIODE
    ANTENNADIFFAREA  0.607200 ;
    ANTENNAGATEAREA  0.607200 ;
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.515000 0.855000 3.280000 ;
    END
  END DIODE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 0.960000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 0.960000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 0.960000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 0.960000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 1.290000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 0.960000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 0.960000 0.085000 ;
      RECT 0.000000  3.985000 0.960000 4.155000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
  END
END sky130_fd_sc_hvl__diode_2
MACRO sky130_fd_sc_hvl__lsbuflv2hv_clkiso_hlkg_3
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__lsbuflv2hv_clkiso_hlkg_3 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  24.96000 BY  8.140000 ;
  SYMMETRY X Y ;
  SITE unithvdbl ;
  PIN A
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 21.070000 5.975000 21.400000 6.455000 ;
    END
  END A
  PIN SLEEP_B
    ANTENNAGATEAREA  0.750000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.315000 5.545000 14.985000 5.875000 ;
    END
  END SLEEP_B
  PIN X
    ANTENNADIFFAREA  2.180000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.060000 0.645000 1.280000 1.920000 ;
        RECT 1.060000 1.920000 2.840000 2.140000 ;
        RECT 1.060000 2.140000 1.280000 5.115000 ;
        RECT 2.620000 0.645000 2.840000 1.920000 ;
        RECT 2.620000 2.140000 2.840000 5.115000 ;
    END
  END X
  PIN LVPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.070000 3.020000 24.890000 3.305000 ;
      LAYER nwell ;
        RECT 17.395000 2.045000 21.695000 6.095000 ;
    END
  END LVPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 7.515000 24.960000 7.885000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 8.025000 24.960000 8.255000 ;
      LAYER pwell ;
        RECT 0.000000 8.055000 24.960000 8.225000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 24.960000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000  0.510000 2.095000 ;
        RECT -0.330000 2.095000 15.395000 5.755000 ;
        RECT -0.330000 5.755000  0.510000 6.255000 ;
        RECT  9.415000 1.705000 15.395000 2.095000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 4.325000 24.960000 4.695000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 24.960000 0.085000 ;
      RECT  0.000000  3.985000  0.685000 4.155000 ;
      RECT  0.000000  8.055000 24.960000 8.225000 ;
      RECT  0.360000  4.155000  0.530000 5.180000 ;
      RECT  1.060000  6.195000  1.280000 6.850000 ;
      RECT  1.060000  6.850000  1.810000 7.180000 ;
      RECT  1.060000  7.180000  1.280000 7.570000 ;
      RECT  1.060000  7.570000 14.885000 7.800000 ;
      RECT  1.655000  4.395000  2.245000 4.625000 ;
      RECT  1.835000  0.255000  2.425000 0.485000 ;
      RECT  1.835000  0.485000  2.065000 1.655000 ;
      RECT  1.835000  2.405000  2.065000 4.395000 ;
      RECT  1.835000  4.625000  2.065000 5.115000 ;
      RECT  1.840000  5.755000  6.520000 5.975000 ;
      RECT  1.840000  5.975000  2.060000 6.525000 ;
      RECT  2.360000  6.195000  2.585000 7.205000 ;
      RECT  2.360000  7.205000  2.580000 7.570000 ;
      RECT  3.010000  1.865000  4.170000 1.920000 ;
      RECT  3.010000  1.920000  5.730000 2.140000 ;
      RECT  3.010000  2.140000  4.170000 2.195000 ;
      RECT  3.035000  0.255000  3.625000 0.485000 ;
      RECT  3.215000  4.395000  3.805000 4.625000 ;
      RECT  3.395000  0.485000  3.625000 1.655000 ;
      RECT  3.395000  2.405000  3.625000 4.395000 ;
      RECT  3.395000  4.625000  3.625000 5.115000 ;
      RECT  3.570000  5.975000  3.790000 7.205000 ;
      RECT  3.950000  0.645000  4.170000 1.865000 ;
      RECT  3.950000  2.195000  4.170000 3.755000 ;
      RECT  4.545000  0.255000  5.135000 0.485000 ;
      RECT  4.725000  0.485000  4.955000 1.655000 ;
      RECT  4.725000  2.405000  4.955000 3.515000 ;
      RECT  4.725000  3.515000  5.310000 3.755000 ;
      RECT  4.750000  6.195000  4.970000 7.570000 ;
      RECT  5.510000  0.645000  5.730000 1.920000 ;
      RECT  5.510000  2.140000  5.730000 3.755000 ;
      RECT  5.930000  5.975000  6.150000 7.205000 ;
      RECT  6.300000  2.185000  6.995000 2.515000 ;
      RECT  6.300000  2.515000  6.520000 5.755000 ;
      RECT  7.075000  2.835000  7.435000 3.065000 ;
      RECT  7.075000  3.065000  7.305000 4.345000 ;
      RECT  7.110000  6.195000  7.330000 7.570000 ;
      RECT  7.205000  2.425000  7.805000 2.655000 ;
      RECT  7.205000  2.655000  7.435000 2.835000 ;
      RECT  7.345000  4.905000  8.080000 5.235000 ;
      RECT  7.575000  1.585000 12.770000 1.805000 ;
      RECT  7.575000  1.805000  7.805000 2.425000 ;
      RECT  7.860000  2.835000  8.080000 4.905000 ;
      RECT  7.860000  5.235000  8.080000 5.755000 ;
      RECT  7.860000  5.755000 12.775000 5.975000 ;
      RECT  8.290000  5.975000  8.510000 7.205000 ;
      RECT  9.135000  3.985000  9.925000 4.155000 ;
      RECT  9.470000  6.195000  9.690000 7.570000 ;
      RECT 10.025000  3.515000 10.615000 3.745000 ;
      RECT 10.210000  2.015000 10.430000 3.515000 ;
      RECT 10.210000  3.745000 10.430000 5.035000 ;
      RECT 10.210000  5.035000 13.550000 5.255000 ;
      RECT 10.650000  5.975000 10.870000 7.205000 ;
      RECT 10.990000  1.805000 11.210000 4.725000 ;
      RECT 11.585000  3.515000 12.175000 3.745000 ;
      RECT 11.770000  2.015000 11.990000 3.515000 ;
      RECT 11.770000  3.745000 11.990000 5.035000 ;
      RECT 11.830000  6.195000 12.050000 7.570000 ;
      RECT 12.550000  1.805000 12.770000 4.725000 ;
      RECT 12.555000  5.975000 12.775000 6.525000 ;
      RECT 13.090000  5.425000 14.105000 5.755000 ;
      RECT 13.145000  3.515000 13.735000 3.745000 ;
      RECT 13.330000  2.015000 13.550000 3.515000 ;
      RECT 13.330000  3.745000 13.550000 5.035000 ;
      RECT 13.335000  6.195000 13.555000 7.570000 ;
      RECT 13.885000  4.265000 14.105000 5.425000 ;
      RECT 13.885000  5.755000 14.105000 6.865000 ;
      RECT 13.965000  1.345000 18.530000 1.395000 ;
      RECT 13.965000  1.395000 19.940000 1.565000 ;
      RECT 13.965000  1.565000 14.295000 2.285000 ;
      RECT 14.295000  4.395000 14.885000 4.625000 ;
      RECT 14.655000  4.265000 14.885000 4.395000 ;
      RECT 14.655000  4.625000 14.885000 5.055000 ;
      RECT 14.665000  6.195000 14.885000 7.570000 ;
      RECT 17.160000  1.735000 19.465000 2.165000 ;
      RECT 17.160000  2.165000 17.380000 5.635000 ;
      RECT 17.160000  5.635000 19.465000 5.805000 ;
      RECT 17.160000  5.805000 18.020000 5.855000 ;
      RECT 17.780000  0.395000 19.950000 0.625000 ;
      RECT 17.780000  0.625000 18.110000 1.175000 ;
      RECT 17.780000  6.915000 18.110000 7.515000 ;
      RECT 17.780000  7.515000 21.375000 7.745000 ;
      RECT 17.785000  4.435000 21.400000 4.605000 ;
      RECT 17.785000  4.605000 18.035000 5.465000 ;
      RECT 17.790000  5.855000 18.020000 6.575000 ;
      RECT 17.790000  6.575000 19.450000 6.745000 ;
      RECT 17.795000  3.905000 20.420000 4.235000 ;
      RECT 17.815000  2.335000 18.065000 3.535000 ;
      RECT 17.815000  3.535000 20.420000 3.705000 ;
      RECT 18.235000  4.775000 18.565000 5.635000 ;
      RECT 18.265000  2.335000 19.940000 2.505000 ;
      RECT 18.265000  2.505000 18.595000 3.365000 ;
      RECT 18.265000  5.975000 19.940000 6.185000 ;
      RECT 18.265000  6.185000 20.900000 6.405000 ;
      RECT 18.280000  0.795000 18.530000 1.345000 ;
      RECT 18.290000  6.745000 18.460000 7.345000 ;
      RECT 18.690000  6.915000 19.020000 7.515000 ;
      RECT 18.710000  0.625000 19.040000 1.225000 ;
      RECT 18.765000  4.605000 18.935000 5.465000 ;
      RECT 18.795000  2.675000 18.965000 3.535000 ;
      RECT 19.135000  4.775000 19.465000 5.635000 ;
      RECT 19.165000  2.505000 19.495000 3.365000 ;
      RECT 19.200000  6.745000 19.450000 7.345000 ;
      RECT 19.270000  0.795000 19.440000 1.395000 ;
      RECT 19.620000  0.625000 19.950000 1.225000 ;
      RECT 19.620000  6.625000 19.950000 7.515000 ;
      RECT 19.665000  3.705000 20.420000 3.905000 ;
      RECT 19.665000  4.235000 20.420000 4.435000 ;
      RECT 19.665000  4.605000 20.420000 5.805000 ;
      RECT 19.695000  2.675000 19.945000 3.020000 ;
      RECT 19.695000  3.020000 20.420000 3.535000 ;
      RECT 19.710000  1.565000 19.940000 2.335000 ;
      RECT 20.170000  5.805000 20.420000 5.935000 ;
      RECT 20.185000  6.625000 20.435000 7.515000 ;
      RECT 20.615000  4.775000 20.900000 6.185000 ;
      RECT 20.615000  6.405000 20.900000 6.625000 ;
      RECT 20.615000  6.625000 20.945000 7.345000 ;
      RECT 21.070000  4.605000 21.400000 5.805000 ;
      RECT 21.125000  6.625000 21.375000 7.515000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.985000  0.325000 4.155000 ;
      RECT  0.155000  8.055000  0.325000 8.225000 ;
      RECT  0.515000  3.985000  0.685000 4.155000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  8.055000  0.805000 8.225000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  7.600000  1.285000 7.770000 ;
      RECT  1.115000  8.055000  1.285000 8.225000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  7.600000  1.765000 7.770000 ;
      RECT  1.595000  8.055000  1.765000 8.225000 ;
      RECT  1.685000  4.425000  1.855000 4.595000 ;
      RECT  1.865000  0.285000  2.035000 0.455000 ;
      RECT  2.045000  4.425000  2.215000 4.595000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  7.600000  2.245000 7.770000 ;
      RECT  2.075000  8.055000  2.245000 8.225000 ;
      RECT  2.225000  0.285000  2.395000 0.455000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  7.600000  2.725000 7.770000 ;
      RECT  2.555000  8.055000  2.725000 8.225000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  7.600000  3.205000 7.770000 ;
      RECT  3.035000  8.055000  3.205000 8.225000 ;
      RECT  3.065000  0.285000  3.235000 0.455000 ;
      RECT  3.245000  4.425000  3.415000 4.595000 ;
      RECT  3.425000  0.285000  3.595000 0.455000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  7.600000  3.685000 7.770000 ;
      RECT  3.515000  8.055000  3.685000 8.225000 ;
      RECT  3.605000  4.425000  3.775000 4.595000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  7.600000  4.165000 7.770000 ;
      RECT  3.995000  8.055000  4.165000 8.225000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  7.600000  4.645000 7.770000 ;
      RECT  4.475000  8.055000  4.645000 8.225000 ;
      RECT  4.575000  0.285000  4.745000 0.455000 ;
      RECT  4.750000  3.545000  4.920000 3.715000 ;
      RECT  4.935000  0.285000  5.105000 0.455000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  7.600000  5.125000 7.770000 ;
      RECT  4.955000  8.055000  5.125000 8.225000 ;
      RECT  5.110000  3.545000  5.280000 3.715000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  7.600000  5.605000 7.770000 ;
      RECT  5.435000  8.055000  5.605000 8.225000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  7.600000  6.085000 7.770000 ;
      RECT  5.915000  8.055000  6.085000 8.225000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  7.600000  6.565000 7.770000 ;
      RECT  6.395000  8.055000  6.565000 8.225000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  7.600000  7.045000 7.770000 ;
      RECT  6.875000  8.055000  7.045000 8.225000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  7.600000  7.525000 7.770000 ;
      RECT  7.355000  8.055000  7.525000 8.225000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  7.600000  8.005000 7.770000 ;
      RECT  7.835000  8.055000  8.005000 8.225000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  7.600000  8.485000 7.770000 ;
      RECT  8.315000  8.055000  8.485000 8.225000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  7.600000  8.965000 7.770000 ;
      RECT  8.795000  8.055000  8.965000 8.225000 ;
      RECT  9.265000  3.985000  9.435000 4.155000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  7.600000  9.445000 7.770000 ;
      RECT  9.275000  8.055000  9.445000 8.225000 ;
      RECT  9.625000  3.985000  9.795000 4.155000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  7.600000  9.925000 7.770000 ;
      RECT  9.755000  8.055000  9.925000 8.225000 ;
      RECT 10.055000  3.545000 10.225000 3.715000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  7.600000 10.405000 7.770000 ;
      RECT 10.235000  8.055000 10.405000 8.225000 ;
      RECT 10.415000  3.545000 10.585000 3.715000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  7.600000 10.885000 7.770000 ;
      RECT 10.715000  8.055000 10.885000 8.225000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  7.600000 11.365000 7.770000 ;
      RECT 11.195000  8.055000 11.365000 8.225000 ;
      RECT 11.615000  3.545000 11.785000 3.715000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  7.600000 11.845000 7.770000 ;
      RECT 11.675000  8.055000 11.845000 8.225000 ;
      RECT 11.975000  3.545000 12.145000 3.715000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  7.600000 12.325000 7.770000 ;
      RECT 12.155000  8.055000 12.325000 8.225000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  7.600000 12.805000 7.770000 ;
      RECT 12.635000  8.055000 12.805000 8.225000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  7.600000 13.285000 7.770000 ;
      RECT 13.115000  8.055000 13.285000 8.225000 ;
      RECT 13.175000  3.545000 13.345000 3.715000 ;
      RECT 13.535000  3.545000 13.705000 3.715000 ;
      RECT 13.590000  7.600000 13.760000 7.770000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  8.055000 13.765000 8.225000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  7.600000 14.245000 7.770000 ;
      RECT 14.075000  8.055000 14.245000 8.225000 ;
      RECT 14.325000  4.425000 14.495000 4.595000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  7.600000 14.725000 7.770000 ;
      RECT 14.555000  8.055000 14.725000 8.225000 ;
      RECT 14.685000  4.425000 14.855000 4.595000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  8.055000 15.205000 8.225000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  8.055000 15.685000 8.225000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000  8.055000 16.165000 8.225000 ;
      RECT 16.475000 -0.085000 16.645000 0.085000 ;
      RECT 16.475000  8.055000 16.645000 8.225000 ;
      RECT 16.955000 -0.085000 17.125000 0.085000 ;
      RECT 16.955000  8.055000 17.125000 8.225000 ;
      RECT 17.435000 -0.085000 17.605000 0.085000 ;
      RECT 17.435000  8.055000 17.605000 8.225000 ;
      RECT 17.820000  0.425000 17.990000 0.595000 ;
      RECT 17.820000  7.545000 17.990000 7.715000 ;
      RECT 17.915000 -0.085000 18.085000 0.085000 ;
      RECT 17.915000  8.055000 18.085000 8.225000 ;
      RECT 18.300000  0.425000 18.470000 0.595000 ;
      RECT 18.300000  7.545000 18.470000 7.715000 ;
      RECT 18.395000 -0.085000 18.565000 0.085000 ;
      RECT 18.395000  8.055000 18.565000 8.225000 ;
      RECT 18.780000  0.425000 18.950000 0.595000 ;
      RECT 18.780000  7.545000 18.950000 7.715000 ;
      RECT 18.875000 -0.085000 19.045000 0.085000 ;
      RECT 18.875000  8.055000 19.045000 8.225000 ;
      RECT 19.260000  0.425000 19.430000 0.595000 ;
      RECT 19.260000  7.545000 19.430000 7.715000 ;
      RECT 19.355000 -0.085000 19.525000 0.085000 ;
      RECT 19.355000  8.055000 19.525000 8.225000 ;
      RECT 19.740000  0.425000 19.910000 0.595000 ;
      RECT 19.740000  7.545000 19.910000 7.715000 ;
      RECT 19.800000  3.070000 19.970000 3.240000 ;
      RECT 19.835000 -0.085000 20.005000 0.085000 ;
      RECT 19.835000  8.055000 20.005000 8.225000 ;
      RECT 20.160000  3.070000 20.330000 3.240000 ;
      RECT 20.220000  7.545000 20.390000 7.715000 ;
      RECT 20.315000 -0.085000 20.485000 0.085000 ;
      RECT 20.315000  8.055000 20.485000 8.225000 ;
      RECT 20.700000  7.545000 20.870000 7.715000 ;
      RECT 20.795000 -0.085000 20.965000 0.085000 ;
      RECT 20.795000  8.055000 20.965000 8.225000 ;
      RECT 21.180000  7.545000 21.350000 7.715000 ;
      RECT 21.275000 -0.085000 21.445000 0.085000 ;
      RECT 21.275000  8.055000 21.445000 8.225000 ;
      RECT 21.755000 -0.085000 21.925000 0.085000 ;
      RECT 21.755000  8.055000 21.925000 8.225000 ;
      RECT 22.235000 -0.085000 22.405000 0.085000 ;
      RECT 22.235000  8.055000 22.405000 8.225000 ;
      RECT 22.715000 -0.085000 22.885000 0.085000 ;
      RECT 22.715000  8.055000 22.885000 8.225000 ;
      RECT 23.195000 -0.085000 23.365000 0.085000 ;
      RECT 23.195000  8.055000 23.365000 8.225000 ;
      RECT 23.675000 -0.085000 23.845000 0.085000 ;
      RECT 23.675000  8.055000 23.845000 8.225000 ;
      RECT 24.155000 -0.085000 24.325000 0.085000 ;
      RECT 24.155000  8.055000 24.325000 8.225000 ;
      RECT 24.635000 -0.085000 24.805000 0.085000 ;
      RECT 24.635000  8.055000 24.805000 8.225000 ;
    LAYER met1 ;
      RECT 0.000000 -0.115000 24.960000 0.115000 ;
      RECT 0.000000  0.255000 24.960000 0.625000 ;
      RECT 0.000000  3.445000 24.960000 3.815000 ;
    LAYER pwell ;
      RECT 0.000000 -0.085000 24.960000 0.085000 ;
  END
END sky130_fd_sc_hvl__lsbuflv2hv_clkiso_hlkg_3
MACRO sky130_fd_sc_hvl__nand2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__nand2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.400000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN A
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.975000 1.525000 2.275000 1.855000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.125000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.550000 1.015000 1.935000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.633750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.220000 1.525000 1.795000 1.695000 ;
        RECT 1.220000 1.695000 1.470000 3.755000 ;
        RECT 1.580000 1.175000 2.180000 1.345000 ;
        RECT 1.580000 1.345000 1.795000 1.525000 ;
        RECT 1.850000 0.515000 2.180000 1.175000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 2.400000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 2.400000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 2.400000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 2.400000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 2.730000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 2.400000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.400000 0.085000 ;
      RECT 0.000000  3.985000 2.400000 4.155000 ;
      RECT 0.090000  0.365000 1.400000 1.345000 ;
      RECT 0.090000  2.175000 1.040000 3.755000 ;
      RECT 1.660000  2.175000 2.250000 3.755000 ;
    LAYER mcon ;
      RECT 0.120000  0.395000 0.290000 0.565000 ;
      RECT 0.120000  3.505000 0.290000 3.675000 ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.480000  0.395000 0.650000 0.565000 ;
      RECT 0.480000  3.505000 0.650000 3.675000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.840000  0.395000 1.010000 0.565000 ;
      RECT 0.840000  3.505000 1.010000 3.675000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.200000  0.395000 1.370000 0.565000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.690000  3.505000 1.860000 3.675000 ;
      RECT 2.050000  3.505000 2.220000 3.675000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
  END
END sky130_fd_sc_hvl__nand2_1
MACRO sky130_fd_sc_hvl__decap_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__decap_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.920000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 1.920000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 1.920000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 1.920000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 1.920000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 2.250000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 1.920000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.920000 0.085000 ;
      RECT 0.000000  3.985000 1.920000 4.155000 ;
      RECT 0.170000  0.365000 1.780000 0.845000 ;
      RECT 0.250000  2.685000 1.700000 3.755000 ;
      RECT 0.475000  0.845000 1.780000 1.250000 ;
      RECT 0.475000  1.250000 0.805000 2.030000 ;
      RECT 1.015000  1.700000 1.345000 2.685000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.215000  0.395000 0.385000 0.565000 ;
      RECT 0.495000  3.560000 0.665000 3.730000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.655000  0.395000 0.825000 0.565000 ;
      RECT 0.860000  3.560000 1.030000 3.730000 ;
      RECT 1.095000  0.395000 1.265000 0.565000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.300000  3.560000 1.470000 3.730000 ;
      RECT 1.510000  0.395000 1.680000 0.565000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
  END
END sky130_fd_sc_hvl__decap_4
MACRO sky130_fd_sc_hvl__decap_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__decap_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 3.840000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 3.840000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 3.840000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 3.840000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 4.170000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 3.840000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.985000 3.840000 4.155000 ;
      RECT 0.500000  2.680000 3.240000 3.750000 ;
      RECT 0.575000  0.360000 3.305000 1.360000 ;
      RECT 0.735000  1.360000 1.065000 2.025000 ;
      RECT 1.470000  1.695000 1.800000 2.680000 ;
      RECT 2.015000  1.360000 2.345000 2.025000 ;
      RECT 2.750000  1.695000 3.080000 2.680000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.705000  3.555000 0.875000 3.725000 ;
      RECT 0.745000  0.390000 0.915000 0.560000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.145000  3.555000 1.315000 3.725000 ;
      RECT 1.185000  0.390000 1.355000 0.560000 ;
      RECT 1.560000  3.555000 1.730000 3.725000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.600000  0.390000 1.770000 0.560000 ;
      RECT 1.985000  3.555000 2.155000 3.725000 ;
      RECT 2.025000  0.390000 2.195000 0.560000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.425000  3.555000 2.595000 3.725000 ;
      RECT 2.465000  0.390000 2.635000 0.560000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 2.840000  3.555000 3.010000 3.725000 ;
      RECT 2.880000  0.390000 3.050000 0.560000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.985000 3.685000 4.155000 ;
  END
END sky130_fd_sc_hvl__decap_8
MACRO sky130_fd_sc_hvl__sdlxtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__sdlxtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.52000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN D
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.040000 2.185000 2.370000 3.260000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.626250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.060000 0.515000 11.400000 3.755000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.515000 1.525000 3.860000 2.495000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  1.005000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.585000 1.835000 2.770000 2.005000 ;
        RECT 0.585000 2.005000 1.795000 2.775000 ;
        RECT 2.600000 1.445000 2.985000 1.695000 ;
        RECT 2.600000 1.695000 2.770000 1.835000 ;
    END
  END SCE
  PIN GATE
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.370000 1.145000 4.665000 2.495000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 11.520000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 11.520000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 11.520000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 11.520000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 11.850000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 11.520000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.520000 0.085000 ;
      RECT  0.000000  3.985000 11.520000 4.155000 ;
      RECT  0.130000  0.495000  0.480000 1.175000 ;
      RECT  0.130000  1.175000  3.335000 1.265000 ;
      RECT  0.130000  1.265000  2.295000 1.345000 ;
      RECT  0.130000  1.345000  0.380000 3.395000 ;
      RECT  0.560000  2.995000  1.510000 3.705000 ;
      RECT  0.660000  0.365000  1.610000 0.995000 ;
      RECT  1.965000  1.095000  3.335000 1.175000 ;
      RECT  1.965000  1.345000  2.295000 1.655000 ;
      RECT  2.420000  0.495000  2.750000 0.745000 ;
      RECT  2.420000  0.745000  3.685000 0.915000 ;
      RECT  2.575000  2.675000  4.665000 2.845000 ;
      RECT  2.575000  2.845000  2.825000 3.725000 ;
      RECT  2.950000  1.905000  3.335000 2.495000 ;
      RECT  3.165000  1.265000  3.335000 1.905000 ;
      RECT  3.365000  3.025000  4.315000 3.725000 ;
      RECT  3.515000  0.915000  3.685000 1.175000 ;
      RECT  3.515000  1.175000  4.200000 1.345000 ;
      RECT  3.865000  0.365000  4.455000 0.975000 ;
      RECT  4.030000  1.345000  4.200000 2.675000 ;
      RECT  4.495000  2.845000  4.665000 3.635000 ;
      RECT  4.495000  3.635000  5.365000 3.805000 ;
      RECT  4.695000  0.515000  5.025000 0.975000 ;
      RECT  4.845000  0.975000  5.015000 1.175000 ;
      RECT  4.845000  1.175000  5.920000 1.345000 ;
      RECT  4.845000  1.345000  5.015000 3.455000 ;
      RECT  5.195000  2.235000  6.065000 2.405000 ;
      RECT  5.195000  2.405000  5.365000 3.635000 ;
      RECT  5.205000  0.365000  5.795000 0.995000 ;
      RECT  5.545000  2.585000  5.715000 3.705000 ;
      RECT  5.590000  1.345000  5.920000 1.845000 ;
      RECT  5.895000  2.405000  6.065000 3.595000 ;
      RECT  5.895000  3.595000  7.250000 3.765000 ;
      RECT  6.045000  0.265000  7.275000 0.435000 ;
      RECT  6.045000  0.435000  6.415000 0.975000 ;
      RECT  6.245000  0.975000  6.415000 2.585000 ;
      RECT  6.245000  2.585000  6.575000 3.415000 ;
      RECT  6.595000  0.615000  6.925000 0.975000 ;
      RECT  6.755000  0.975000  6.925000 2.925000 ;
      RECT  6.755000  2.925000  7.250000 3.595000 ;
      RECT  7.105000  0.435000  7.275000 1.585000 ;
      RECT  7.105000  1.585000  8.010000 1.755000 ;
      RECT  7.455000  0.495000  7.705000 1.075000 ;
      RECT  7.455000  1.075000  8.360000 1.245000 ;
      RECT  7.700000  2.925000  8.030000 3.755000 ;
      RECT  7.840000  1.755000  8.010000 2.215000 ;
      RECT  7.840000  2.215000  8.570000 2.475000 ;
      RECT  7.860000  2.655000  8.920000 2.825000 ;
      RECT  7.860000  2.825000  8.030000 2.925000 ;
      RECT  8.190000  1.245000  8.360000 1.835000 ;
      RECT  8.190000  1.835000 10.200000 2.005000 ;
      RECT  8.245000  0.365000  9.195000 0.895000 ;
      RECT  8.540000  1.075000  8.870000 1.405000 ;
      RECT  8.540000  1.405000 10.550000 1.575000 ;
      RECT  8.540000  1.575000  8.870000 1.655000 ;
      RECT  8.685000  3.005000  9.635000 3.705000 ;
      RECT  8.750000  2.005000  8.920000 2.655000 ;
      RECT  9.385000  2.185000 10.550000 2.355000 ;
      RECT  9.385000  2.355000  9.715000 2.675000 ;
      RECT  9.415000  0.845000  9.745000 1.405000 ;
      RECT  9.870000  1.755000 10.200000 1.835000 ;
      RECT  9.895000  2.535000 10.845000 3.755000 ;
      RECT  9.925000  0.365000 10.875000 1.225000 ;
      RECT 10.380000  1.575000 10.550000 2.185000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.985000  0.325000 4.155000 ;
      RECT  0.590000  3.505000  0.760000 3.675000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.985000  0.805000 4.155000 ;
      RECT  0.690000  0.395000  0.860000 0.565000 ;
      RECT  0.950000  3.505000  1.120000 3.675000 ;
      RECT  1.050000  0.395000  1.220000 0.565000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.985000  1.285000 4.155000 ;
      RECT  1.310000  3.505000  1.480000 3.675000 ;
      RECT  1.410000  0.395000  1.580000 0.565000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.985000  1.765000 4.155000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.985000  2.245000 4.155000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.985000  2.725000 4.155000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.985000  3.205000 4.155000 ;
      RECT  3.395000  3.505000  3.565000 3.675000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.985000  3.685000 4.155000 ;
      RECT  3.755000  3.505000  3.925000 3.675000 ;
      RECT  3.895000  0.395000  4.065000 0.565000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.985000  4.165000 4.155000 ;
      RECT  4.115000  3.505000  4.285000 3.675000 ;
      RECT  4.255000  0.395000  4.425000 0.565000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.985000  4.645000 4.155000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.985000  5.125000 4.155000 ;
      RECT  5.235000  0.395000  5.405000 0.565000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.985000  5.605000 4.155000 ;
      RECT  5.545000  3.505000  5.715000 3.675000 ;
      RECT  5.595000  0.395000  5.765000 0.565000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.985000  6.085000 4.155000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.985000  6.565000 4.155000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.985000  7.045000 4.155000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.985000  7.525000 4.155000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.985000  8.005000 4.155000 ;
      RECT  8.275000  0.395000  8.445000 0.565000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.985000  8.485000 4.155000 ;
      RECT  8.635000  0.395000  8.805000 0.565000 ;
      RECT  8.715000  3.505000  8.885000 3.675000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.985000  8.965000 4.155000 ;
      RECT  8.995000  0.395000  9.165000 0.565000 ;
      RECT  9.075000  3.505000  9.245000 3.675000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.985000  9.445000 4.155000 ;
      RECT  9.435000  3.505000  9.605000 3.675000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.985000  9.925000 4.155000 ;
      RECT  9.925000  3.505000 10.095000 3.675000 ;
      RECT  9.955000  0.395000 10.125000 0.565000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.985000 10.405000 4.155000 ;
      RECT 10.285000  3.505000 10.455000 3.675000 ;
      RECT 10.315000  0.395000 10.485000 0.565000 ;
      RECT 10.645000  3.505000 10.815000 3.675000 ;
      RECT 10.675000  0.395000 10.845000 0.565000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.985000 10.885000 4.155000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.985000 11.365000 4.155000 ;
  END
END sky130_fd_sc_hvl__sdlxtp_1
MACRO sky130_fd_sc_hvl__sdlclkp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__sdlclkp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN GATE
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.475000 1.535000 1.805000 2.125000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.596250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.590000 0.515000 10.955000 1.215000 ;
        RECT 10.590000 1.895000 10.955000 3.735000 ;
        RECT 10.685000 1.215000 10.955000 1.895000 ;
    END
  END GCLK
  PIN SCE
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595000 1.535000 0.925000 2.125000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  1.170000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.320000 1.465000 4.650000 1.975000 ;
        RECT 9.195000 3.125000 9.560000 3.445000 ;
        RECT 9.310000 1.725000 9.640000 2.025000 ;
        RECT 9.310000 2.025000 9.560000 3.125000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 11.040000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 11.040000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 11.040000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 11.040000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 11.370000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 11.040000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 11.040000 0.085000 ;
      RECT 0.000000  3.985000 11.040000 4.155000 ;
      RECT 0.290000  0.840000  0.620000 1.195000 ;
      RECT 0.290000  1.195000  2.145000 1.365000 ;
      RECT 0.290000  2.295000  0.620000 3.445000 ;
      RECT 0.290000  3.445000  1.985000 3.615000 ;
      RECT 0.290000  3.615000  4.290000 3.815000 ;
      RECT 0.730000  0.365000  1.740000 0.625000 ;
      RECT 1.070000  0.625000  1.400000 1.025000 ;
      RECT 1.850000  0.840000  2.145000 1.195000 ;
      RECT 1.850000  2.295000  2.145000 3.055000 ;
      RECT 1.975000  1.365000  2.145000 2.295000 ;
      RECT 2.115000  0.365000  3.770000 0.535000 ;
      RECT 2.115000  0.535000  2.825000 0.670000 ;
      RECT 2.155000  3.225000  3.455000 3.445000 ;
      RECT 2.555000  1.555000  3.065000 1.885000 ;
      RECT 2.630000  0.840000  2.960000 1.555000 ;
      RECT 2.630000  1.885000  2.960000 3.055000 ;
      RECT 3.180000  0.705000  3.430000 1.080000 ;
      RECT 3.235000  1.080000  3.430000 2.145000 ;
      RECT 3.235000  2.145000  4.650000 2.315000 ;
      RECT 3.235000  2.315000  3.455000 3.225000 ;
      RECT 3.600000  0.535000  3.770000 1.125000 ;
      RECT 3.600000  1.125000  5.030000 1.295000 ;
      RECT 3.600000  1.295000  3.930000 1.965000 ;
      RECT 3.625000  3.445000  4.290000 3.615000 ;
      RECT 3.940000  0.255000  4.885000 0.535000 ;
      RECT 3.940000  0.535000  4.610000 0.625000 ;
      RECT 3.940000  0.625000  4.290000 0.955000 ;
      RECT 3.960000  2.485000  4.290000 3.445000 ;
      RECT 4.480000  2.315000  4.650000 3.385000 ;
      RECT 4.480000  3.385000  6.475000 3.555000 ;
      RECT 4.780000  0.705000  5.030000 1.125000 ;
      RECT 4.820000  1.295000  5.030000 3.005000 ;
      RECT 4.820000  3.005000  6.135000 3.215000 ;
      RECT 5.055000  0.255000  5.620000 0.535000 ;
      RECT 5.335000  0.535000  5.620000 1.195000 ;
      RECT 5.335000  1.195000  7.450000 1.365000 ;
      RECT 5.335000  1.365000  5.505000 2.330000 ;
      RECT 5.335000  2.330000  5.620000 2.660000 ;
      RECT 5.675000  1.615000  6.265000 1.945000 ;
      RECT 5.790000  0.255000  7.110000 0.625000 ;
      RECT 6.095000  1.945000  6.265000 2.425000 ;
      RECT 6.095000  2.425000  6.475000 2.595000 ;
      RECT 6.305000  2.595000  6.475000 3.385000 ;
      RECT 6.475000  1.535000  6.805000 1.875000 ;
      RECT 6.475000  1.875000  7.890000 2.085000 ;
      RECT 6.645000  3.445000  9.025000 3.615000 ;
      RECT 6.645000  3.615000 10.420000 3.815000 ;
      RECT 6.780000  0.625000  7.110000 1.025000 ;
      RECT 6.780000  2.330000  7.110000 3.445000 ;
      RECT 7.085000  1.365000  7.450000 1.655000 ;
      RECT 7.280000  0.355000  7.870000 0.670000 ;
      RECT 7.280000  0.670000  7.450000 1.195000 ;
      RECT 7.620000  0.840000  7.890000 1.615000 ;
      RECT 7.620000  1.615000  8.745000 1.825000 ;
      RECT 7.620000  1.825000  7.890000 1.875000 ;
      RECT 7.620000  2.085000  7.890000 2.660000 ;
      RECT 8.040000  0.255000 10.420000 0.625000 ;
      RECT 8.110000  0.885000  9.140000 1.215000 ;
      RECT 8.110000  2.225000  8.440000 3.445000 ;
      RECT 8.415000  1.385000  8.745000 1.615000 ;
      RECT 8.415000  1.825000  8.745000 2.055000 ;
      RECT 8.915000  1.215000  9.140000 1.385000 ;
      RECT 8.915000  1.385000 10.515000 1.555000 ;
      RECT 8.915000  1.555000  9.140000 2.955000 ;
      RECT 9.730000  0.625000 10.060000 1.215000 ;
      RECT 9.730000  2.195000 10.060000 3.445000 ;
      RECT 9.730000  3.445000 10.420000 3.615000 ;
      RECT 9.905000  1.555000 10.515000 1.725000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.985000  0.325000 4.155000 ;
      RECT  0.380000  3.475000  0.550000 3.645000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.985000  0.805000 4.155000 ;
      RECT  0.740000  3.475000  0.910000 3.645000 ;
      RECT  0.790000  0.425000  0.960000 0.595000 ;
      RECT  1.100000  3.475000  1.270000 3.645000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.985000  1.285000 4.155000 ;
      RECT  1.150000  0.425000  1.320000 0.595000 ;
      RECT  1.460000  3.475000  1.630000 3.645000 ;
      RECT  1.510000  0.425000  1.680000 0.595000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.985000  1.765000 4.155000 ;
      RECT  1.820000  3.615000  1.990000 3.785000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.985000  2.245000 4.155000 ;
      RECT  2.180000  3.615000  2.350000 3.785000 ;
      RECT  2.540000  3.615000  2.710000 3.785000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.985000  2.725000 4.155000 ;
      RECT  2.955000  3.615000  3.125000 3.785000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.985000  3.205000 4.155000 ;
      RECT  3.315000  3.615000  3.485000 3.785000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.985000  3.685000 4.155000 ;
      RECT  3.675000  3.475000  3.845000 3.645000 ;
      RECT  3.955000  0.425000  4.125000 0.595000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.985000  4.165000 4.155000 ;
      RECT  4.035000  3.475000  4.205000 3.645000 ;
      RECT  4.315000  0.425000  4.485000 0.595000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.985000  4.645000 4.155000 ;
      RECT  4.675000  0.355000  4.845000 0.525000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.985000  5.125000 4.155000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.985000  5.605000 4.155000 ;
      RECT  5.830000  0.355000  6.000000 0.525000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.985000  6.085000 4.155000 ;
      RECT  6.190000  0.355000  6.360000 0.525000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.985000  6.565000 4.155000 ;
      RECT  6.550000  0.425000  6.720000 0.595000 ;
      RECT  6.675000  3.475000  6.845000 3.645000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.985000  7.045000 4.155000 ;
      RECT  6.910000  0.425000  7.080000 0.595000 ;
      RECT  7.035000  3.475000  7.205000 3.645000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.985000  7.525000 4.155000 ;
      RECT  7.395000  3.545000  7.565000 3.715000 ;
      RECT  7.755000  3.545000  7.925000 3.715000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.985000  8.005000 4.155000 ;
      RECT  8.060000  0.355000  8.230000 0.525000 ;
      RECT  8.115000  3.475000  8.285000 3.645000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.985000  8.485000 4.155000 ;
      RECT  8.420000  0.355000  8.590000 0.525000 ;
      RECT  8.475000  3.475000  8.645000 3.645000 ;
      RECT  8.780000  0.355000  8.950000 0.525000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.985000  8.965000 4.155000 ;
      RECT  9.140000  0.355000  9.310000 0.525000 ;
      RECT  9.155000  3.615000  9.325000 3.785000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.985000  9.445000 4.155000 ;
      RECT  9.500000  0.425000  9.670000 0.595000 ;
      RECT  9.515000  3.615000  9.685000 3.785000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.985000  9.925000 4.155000 ;
      RECT  9.860000  0.425000 10.030000 0.595000 ;
      RECT  9.875000  3.475000 10.045000 3.645000 ;
      RECT 10.220000  0.425000 10.390000 0.595000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.475000 10.405000 3.645000 ;
      RECT 10.235000  3.985000 10.405000 4.155000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.985000 10.885000 4.155000 ;
  END
END sky130_fd_sc_hvl__sdlclkp_1
MACRO sky130_fd_sc_hvl__dfstp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__dfstp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.88000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN D
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.505000 1.525000 2.835000 2.095000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.478750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.420000 0.645000 14.770000 3.615000 ;
    END
  END Q
  PIN SET_B
    ANTENNAGATEAREA  0.840000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  7.165000 1.555000  8.100000 1.795000 ;
        RECT  7.930000 0.840000 11.160000 1.010000 ;
        RECT  7.930000 1.010000  8.100000 1.555000 ;
        RECT  8.285000 0.555000 11.160000 0.840000 ;
        RECT 10.885000 1.010000 11.160000 1.040000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.545000 2.075000 0.875000 2.745000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 14.880000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 14.880000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 14.880000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 14.880000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000  5.145000 2.245000 ;
        RECT -0.330000 2.245000 15.210000 4.485000 ;
        RECT  7.170000 1.885000 15.210000 2.245000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 14.880000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 14.880000 0.085000 ;
      RECT  0.000000  3.985000 14.880000 4.155000 ;
      RECT  0.115000  0.615000  0.380000 1.295000 ;
      RECT  0.115000  1.295000  1.510000 1.465000 ;
      RECT  0.115000  1.465000  0.365000 3.735000 ;
      RECT  0.545000  2.925000  1.495000 3.755000 ;
      RECT  0.570000  0.365000  1.160000 1.115000 ;
      RECT  1.180000  1.465000  1.510000 1.895000 ;
      RECT  1.340000  0.265000  2.290000 0.435000 ;
      RECT  1.340000  0.435000  1.510000 1.295000 ;
      RECT  1.675000  2.945000  2.005000 3.735000 ;
      RECT  1.690000  0.615000  1.940000 2.275000 ;
      RECT  1.690000  2.275000  2.835000 2.445000 ;
      RECT  1.690000  2.445000  2.005000 2.945000 ;
      RECT  2.120000  0.435000  2.290000 1.175000 ;
      RECT  2.120000  1.175000  3.185000 1.345000 ;
      RECT  2.235000  2.625000  2.485000 3.705000 ;
      RECT  2.470000  0.365000  3.005000 0.995000 ;
      RECT  2.665000  2.445000  2.835000 3.755000 ;
      RECT  3.015000  1.345000  3.185000 3.285000 ;
      RECT  3.015000  3.285000  5.005000 3.615000 ;
      RECT  3.185000  0.495000  3.535000 0.995000 ;
      RECT  3.365000  0.995000  3.535000 3.105000 ;
      RECT  3.715000  1.085000  3.885000 3.285000 ;
      RECT  4.065000  0.495000  4.315000 0.965000 ;
      RECT  4.065000  0.965000  6.315000 1.135000 ;
      RECT  4.065000  1.135000  4.235000 2.605000 ;
      RECT  4.065000  2.605000  4.395000 3.105000 ;
      RECT  4.415000  1.495000  4.655000 1.805000 ;
      RECT  4.415000  1.805000  6.985000 1.975000 ;
      RECT  4.415000  1.975000  4.655000 2.165000 ;
      RECT  4.835000  2.155000  6.635000 2.325000 ;
      RECT  4.835000  2.325000  5.005000 3.285000 ;
      RECT  4.855000  0.365000  5.805000 0.785000 ;
      RECT  5.135000  1.315000  5.865000 1.625000 ;
      RECT  5.185000  2.505000  6.285000 2.675000 ;
      RECT  5.185000  2.675000  5.425000 3.555000 ;
      RECT  5.605000  2.855000  5.935000 3.705000 ;
      RECT  5.985000  0.265000  6.315000 0.965000 ;
      RECT  6.115000  2.675000  6.895000 2.845000 ;
      RECT  6.465000  2.325000  8.960000 2.495000 ;
      RECT  6.565000  2.845000  6.895000 3.105000 ;
      RECT  6.800000  0.365000  7.750000 1.375000 ;
      RECT  6.815000  1.975000  8.450000 2.145000 ;
      RECT  7.075000  2.675000  8.025000 3.705000 ;
      RECT  8.280000  1.545000  8.785000 1.705000 ;
      RECT  8.280000  1.705000  9.310000 1.875000 ;
      RECT  8.280000  1.875000  8.450000 1.975000 ;
      RECT  8.630000  2.085000  8.960000 2.325000 ;
      RECT  8.695000  2.675000  9.310000 2.845000 ;
      RECT  8.695000  2.845000  8.865000 3.595000 ;
      RECT  8.695000  3.595000  9.825000 3.805000 ;
      RECT  9.025000  1.190000  9.660000 1.475000 ;
      RECT  9.045000  3.025000  9.660000 3.415000 ;
      RECT  9.140000  1.875000  9.310000 2.675000 ;
      RECT  9.490000  1.475000  9.660000 2.315000 ;
      RECT  9.490000  2.315000 12.210000 2.485000 ;
      RECT  9.490000  2.485000  9.660000 3.025000 ;
      RECT 10.010000  2.665000 10.960000 3.705000 ;
      RECT 10.305000  1.545000 10.635000 1.655000 ;
      RECT 10.305000  1.655000 12.560000 1.825000 ;
      RECT 10.305000  1.825000 10.635000 2.135000 ;
      RECT 11.300000  3.255000 11.550000 3.755000 ;
      RECT 11.340000  0.365000 11.930000 1.475000 ;
      RECT 11.380000  3.005000 12.560000 3.175000 ;
      RECT 11.380000  3.175000 11.550000 3.255000 ;
      RECT 11.410000  2.485000 12.210000 2.675000 ;
      RECT 11.410000  2.675000 11.740000 2.825000 ;
      RECT 11.730000  3.355000 12.680000 3.735000 ;
      RECT 11.880000  2.005000 12.210000 2.315000 ;
      RECT 12.120000  0.975000 12.450000 1.655000 ;
      RECT 12.390000  1.825000 12.560000 3.005000 ;
      RECT 12.745000  0.975000 13.075000 1.475000 ;
      RECT 12.865000  1.475000 13.075000 2.225000 ;
      RECT 12.865000  2.225000 14.240000 2.395000 ;
      RECT 12.865000  2.395000 13.115000 3.365000 ;
      RECT 13.255000  0.365000 14.205000 1.475000 ;
      RECT 13.295000  2.575000 14.240000 3.705000 ;
      RECT 13.910000  1.725000 14.240000 2.225000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.985000  0.325000 4.155000 ;
      RECT  0.575000  3.505000  0.745000 3.675000 ;
      RECT  0.600000  0.395000  0.770000 0.565000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.985000  0.805000 4.155000 ;
      RECT  0.935000  3.505000  1.105000 3.675000 ;
      RECT  0.960000  0.395000  1.130000 0.565000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.985000  1.285000 4.155000 ;
      RECT  1.295000  3.505000  1.465000 3.675000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.985000  1.765000 4.155000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.985000  2.245000 4.155000 ;
      RECT  2.265000  3.505000  2.435000 3.675000 ;
      RECT  2.470000  0.395000  2.640000 0.565000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.985000  2.725000 4.155000 ;
      RECT  2.830000  0.395000  3.000000 0.565000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.985000  3.205000 4.155000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.985000  3.685000 4.155000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.985000  4.165000 4.155000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.985000  4.645000 4.155000 ;
      RECT  4.885000  0.395000  5.055000 0.565000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.985000  5.125000 4.155000 ;
      RECT  5.245000  0.395000  5.415000 0.565000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.985000  5.605000 4.155000 ;
      RECT  5.605000  0.395000  5.775000 0.565000 ;
      RECT  5.635000  3.505000  5.805000 3.675000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.985000  6.085000 4.155000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.985000  6.565000 4.155000 ;
      RECT  6.830000  0.395000  7.000000 0.565000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.985000  7.045000 4.155000 ;
      RECT  7.105000  3.505000  7.275000 3.675000 ;
      RECT  7.190000  0.395000  7.360000 0.565000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.985000  7.525000 4.155000 ;
      RECT  7.465000  3.505000  7.635000 3.675000 ;
      RECT  7.550000  0.395000  7.720000 0.565000 ;
      RECT  7.825000  3.505000  7.995000 3.675000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.985000  8.005000 4.155000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.985000  8.485000 4.155000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.985000  8.965000 4.155000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.985000  9.445000 4.155000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.985000  9.925000 4.155000 ;
      RECT 10.040000  3.505000 10.210000 3.675000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.985000 10.405000 4.155000 ;
      RECT 10.400000  3.505000 10.570000 3.675000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.985000 10.885000 4.155000 ;
      RECT 10.760000  3.505000 10.930000 3.675000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.985000 11.365000 4.155000 ;
      RECT 11.370000  0.395000 11.540000 0.565000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.985000 11.845000 4.155000 ;
      RECT 11.730000  0.395000 11.900000 0.565000 ;
      RECT 11.760000  3.505000 11.930000 3.675000 ;
      RECT 12.120000  3.505000 12.290000 3.675000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.985000 12.325000 4.155000 ;
      RECT 12.480000  3.505000 12.650000 3.675000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.985000 12.805000 4.155000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.985000 13.285000 4.155000 ;
      RECT 13.285000  0.395000 13.455000 0.565000 ;
      RECT 13.320000  3.505000 13.490000 3.675000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.985000 13.765000 4.155000 ;
      RECT 13.645000  0.395000 13.815000 0.565000 ;
      RECT 13.680000  3.505000 13.850000 3.675000 ;
      RECT 14.005000  0.395000 14.175000 0.565000 ;
      RECT 14.040000  3.505000 14.210000 3.675000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.985000 14.245000 4.155000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.985000 14.725000 4.155000 ;
  END
END sky130_fd_sc_hvl__dfstp_1
MACRO sky130_fd_sc_hvl__dlclkp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__dlclkp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN GATE
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.610000 1.385000 0.940000 2.200000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.596250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.630000 0.515000 9.995000 1.215000 ;
        RECT 9.630000 1.895000 9.995000 3.735000 ;
        RECT 9.725000 1.215000 9.995000 1.895000 ;
    END
  END GCLK
  PIN CLK
    ANTENNAGATEAREA  1.170000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.360000 1.465000 3.690000 1.975000 ;
        RECT 8.235000 3.125000 8.600000 3.445000 ;
        RECT 8.350000 1.725000 8.680000 2.025000 ;
        RECT 8.350000 2.025000 8.600000 3.125000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 10.080000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 10.080000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 10.080000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 10.080000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 10.410000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 10.080000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.080000 0.085000 ;
      RECT 0.000000  3.985000 10.080000 4.155000 ;
      RECT 0.110000  2.200000  0.440000 3.445000 ;
      RECT 0.110000  3.445000  1.025000 3.555000 ;
      RECT 0.110000  3.555000  3.330000 3.815000 ;
      RECT 0.140000  0.365000  0.765000 0.625000 ;
      RECT 0.140000  0.625000  0.470000 1.170000 ;
      RECT 1.155000  0.365000  2.810000 0.535000 ;
      RECT 1.155000  0.535000  1.865000 0.670000 ;
      RECT 1.195000  3.165000  2.495000 3.385000 ;
      RECT 1.595000  1.555000  2.105000 1.885000 ;
      RECT 1.670000  0.840000  2.000000 1.555000 ;
      RECT 1.670000  1.885000  2.000000 2.995000 ;
      RECT 2.220000  0.705000  2.470000 1.080000 ;
      RECT 2.275000  1.080000  2.470000 2.145000 ;
      RECT 2.275000  2.145000  3.690000 2.315000 ;
      RECT 2.275000  2.315000  2.495000 3.165000 ;
      RECT 2.640000  0.535000  2.810000 1.125000 ;
      RECT 2.640000  1.125000  4.070000 1.295000 ;
      RECT 2.640000  1.295000  2.970000 1.965000 ;
      RECT 2.665000  3.445000  3.330000 3.555000 ;
      RECT 2.980000  0.255000  3.925000 0.535000 ;
      RECT 2.980000  0.535000  3.650000 0.625000 ;
      RECT 2.980000  0.625000  3.330000 0.955000 ;
      RECT 3.000000  2.485000  3.330000 3.445000 ;
      RECT 3.520000  2.315000  3.690000 3.385000 ;
      RECT 3.520000  3.385000  5.515000 3.555000 ;
      RECT 3.820000  0.705000  4.070000 1.125000 ;
      RECT 3.860000  1.295000  4.070000 3.005000 ;
      RECT 3.860000  3.005000  5.175000 3.215000 ;
      RECT 4.095000  0.255000  4.660000 0.535000 ;
      RECT 4.375000  0.535000  4.660000 1.195000 ;
      RECT 4.375000  1.195000  6.490000 1.365000 ;
      RECT 4.375000  1.365000  4.545000 2.330000 ;
      RECT 4.375000  2.330000  4.660000 2.660000 ;
      RECT 4.715000  1.615000  5.305000 1.945000 ;
      RECT 4.830000  0.255000  6.150000 0.625000 ;
      RECT 5.135000  1.945000  5.305000 2.425000 ;
      RECT 5.135000  2.425000  5.515000 2.595000 ;
      RECT 5.345000  2.595000  5.515000 3.385000 ;
      RECT 5.515000  1.535000  5.845000 1.875000 ;
      RECT 5.515000  1.875000  6.930000 2.085000 ;
      RECT 5.685000  3.445000  8.065000 3.615000 ;
      RECT 5.685000  3.615000  9.460000 3.815000 ;
      RECT 5.820000  0.625000  6.150000 1.025000 ;
      RECT 5.820000  2.330000  6.150000 3.445000 ;
      RECT 6.125000  1.365000  6.490000 1.655000 ;
      RECT 6.320000  0.355000  6.910000 0.670000 ;
      RECT 6.320000  0.670000  6.490000 1.195000 ;
      RECT 6.660000  0.840000  6.930000 1.615000 ;
      RECT 6.660000  1.615000  7.785000 1.825000 ;
      RECT 6.660000  1.825000  6.930000 1.875000 ;
      RECT 6.660000  2.085000  6.930000 2.660000 ;
      RECT 7.080000  0.255000  9.460000 0.625000 ;
      RECT 7.150000  0.885000  8.180000 1.215000 ;
      RECT 7.150000  2.225000  7.480000 3.445000 ;
      RECT 7.455000  1.385000  7.785000 1.615000 ;
      RECT 7.455000  1.825000  7.785000 2.055000 ;
      RECT 7.955000  1.215000  8.180000 1.385000 ;
      RECT 7.955000  1.385000  9.555000 1.555000 ;
      RECT 7.955000  1.555000  8.180000 2.955000 ;
      RECT 8.770000  0.625000  9.100000 1.215000 ;
      RECT 8.770000  2.195000  9.100000 3.445000 ;
      RECT 8.770000  3.445000  9.460000 3.615000 ;
      RECT 8.945000  1.555000  9.555000 1.725000 ;
    LAYER mcon ;
      RECT 0.140000  3.475000 0.310000 3.645000 ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.985000 0.325000 4.155000 ;
      RECT 0.175000  0.425000 0.345000 0.595000 ;
      RECT 0.500000  3.475000 0.670000 3.645000 ;
      RECT 0.535000  0.425000 0.705000 0.595000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.985000 0.805000 4.155000 ;
      RECT 0.860000  3.600000 1.030000 3.770000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.985000 1.285000 4.155000 ;
      RECT 1.220000  3.600000 1.390000 3.770000 ;
      RECT 1.580000  3.600000 1.750000 3.770000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.985000 1.765000 4.155000 ;
      RECT 1.995000  3.600000 2.165000 3.770000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.985000 2.245000 4.155000 ;
      RECT 2.355000  3.600000 2.525000 3.770000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.985000 2.725000 4.155000 ;
      RECT 2.715000  3.475000 2.885000 3.645000 ;
      RECT 2.995000  0.425000 3.165000 0.595000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.985000 3.205000 4.155000 ;
      RECT 3.075000  3.475000 3.245000 3.645000 ;
      RECT 3.355000  0.425000 3.525000 0.595000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.985000 3.685000 4.155000 ;
      RECT 3.715000  0.355000 3.885000 0.525000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.985000 4.165000 4.155000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.985000 4.645000 4.155000 ;
      RECT 4.870000  0.355000 5.040000 0.525000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.985000 5.125000 4.155000 ;
      RECT 5.230000  0.355000 5.400000 0.525000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.985000 5.605000 4.155000 ;
      RECT 5.590000  0.425000 5.760000 0.595000 ;
      RECT 5.715000  3.475000 5.885000 3.645000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.985000 6.085000 4.155000 ;
      RECT 5.950000  0.425000 6.120000 0.595000 ;
      RECT 6.075000  3.475000 6.245000 3.645000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.985000 6.565000 4.155000 ;
      RECT 6.435000  3.545000 6.605000 3.715000 ;
      RECT 6.795000  3.545000 6.965000 3.715000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.985000 7.045000 4.155000 ;
      RECT 7.100000  0.355000 7.270000 0.525000 ;
      RECT 7.155000  3.475000 7.325000 3.645000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.985000 7.525000 4.155000 ;
      RECT 7.460000  0.355000 7.630000 0.525000 ;
      RECT 7.515000  3.475000 7.685000 3.645000 ;
      RECT 7.820000  0.355000 7.990000 0.525000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.985000 8.005000 4.155000 ;
      RECT 8.180000  0.355000 8.350000 0.525000 ;
      RECT 8.195000  3.615000 8.365000 3.785000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.985000 8.485000 4.155000 ;
      RECT 8.540000  0.425000 8.710000 0.595000 ;
      RECT 8.555000  3.615000 8.725000 3.785000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.985000 8.965000 4.155000 ;
      RECT 8.900000  0.425000 9.070000 0.595000 ;
      RECT 8.915000  3.475000 9.085000 3.645000 ;
      RECT 9.260000  0.425000 9.430000 0.595000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.475000 9.445000 3.645000 ;
      RECT 9.275000  3.985000 9.445000 4.155000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000  3.985000 9.925000 4.155000 ;
  END
END sky130_fd_sc_hvl__dlclkp_1
MACRO sky130_fd_sc_hvl__dfxbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hvl__dfxbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.92000 BY  4.070000 ;
  SYMMETRY X Y ;
  SITE unithv ;
  PIN D
    ANTENNAGATEAREA  0.420000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.545000 3.350000 2.125000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.596250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.455000 0.675000 10.890000 1.465000 ;
        RECT 10.455000 2.195000 10.890000 3.735000 ;
        RECT 10.685000 1.465000 10.890000 2.195000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.626250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.460000 2.175000 13.810000 3.755000 ;
        RECT 13.480000 0.675000 13.810000 2.175000 ;
    END
  END Q_N
  PIN CLK
    ANTENNAGATEAREA  0.585000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.560000 1.550000 0.890000 2.220000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.255000 13.920000 0.625000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.115000 13.920000 0.115000 ;
      LAYER pwell ;
        RECT 0.000000 -0.085000 13.920000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.955000 13.920000 4.185000 ;
      LAYER nwell ;
        RECT -0.330000 1.885000 14.250000 4.485000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.445000 13.920000 3.815000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 13.920000 0.085000 ;
      RECT  0.000000  3.985000 13.920000 4.155000 ;
      RECT  0.110000  0.540000  0.440000 1.200000 ;
      RECT  0.110000  1.200000  1.545000 1.370000 ;
      RECT  0.110000  1.370000  0.380000 3.230000 ;
      RECT  0.570000  2.400000  1.160000 3.705000 ;
      RECT  0.620000  0.365000  1.570000 1.020000 ;
      RECT  1.215000  1.370000  1.545000 1.870000 ;
      RECT  1.340000  1.870000  1.510000 3.410000 ;
      RECT  1.340000  3.410000  2.290000 3.580000 ;
      RECT  1.690000  2.400000  1.940000 3.230000 ;
      RECT  1.750000  0.520000  1.920000 1.195000 ;
      RECT  1.750000  1.195000  3.340000 1.365000 ;
      RECT  1.750000  1.365000  1.940000 2.400000 ;
      RECT  2.100000  0.365000  2.990000 1.015000 ;
      RECT  2.120000  2.305000  3.350000 2.475000 ;
      RECT  2.120000  2.475000  2.290000 3.410000 ;
      RECT  2.470000  2.655000  3.000000 3.705000 ;
      RECT  3.170000  0.265000  4.980000 0.435000 ;
      RECT  3.170000  0.435000  3.340000 1.195000 ;
      RECT  3.180000  2.475000  3.350000 3.335000 ;
      RECT  3.180000  3.335000  5.085000 3.505000 ;
      RECT  3.520000  0.615000  3.850000 0.935000 ;
      RECT  3.530000  0.935000  3.700000 2.655000 ;
      RECT  3.530000  2.655000  3.770000 3.155000 ;
      RECT  3.880000  1.115000  4.120000 1.785000 ;
      RECT  3.950000  1.785000  4.120000 3.335000 ;
      RECT  4.300000  0.615000  4.630000 1.015000 ;
      RECT  4.300000  1.015000  4.470000 1.905000 ;
      RECT  4.300000  1.905000  6.540000 2.075000 ;
      RECT  4.300000  2.075000  4.550000 3.155000 ;
      RECT  4.650000  1.195000  4.980000 1.245000 ;
      RECT  4.650000  1.245000  6.485000 1.415000 ;
      RECT  4.650000  1.415000  4.980000 1.725000 ;
      RECT  4.755000  2.255000  5.085000 2.635000 ;
      RECT  4.755000  2.635000  6.565000 2.805000 ;
      RECT  4.755000  2.805000  5.085000 3.335000 ;
      RECT  4.810000  0.435000  4.980000 1.195000 ;
      RECT  5.185000  0.365000  6.135000 1.065000 ;
      RECT  5.265000  2.985000  6.215000 3.715000 ;
      RECT  5.435000  2.255000  5.765000 2.285000 ;
      RECT  5.435000  2.285000  6.915000 2.455000 ;
      RECT  6.210000  1.595000  6.540000 1.905000 ;
      RECT  6.210000  2.075000  6.540000 2.105000 ;
      RECT  6.315000  0.265000  7.345000 0.435000 ;
      RECT  6.315000  0.435000  6.485000 1.245000 ;
      RECT  6.395000  2.805000  6.565000 3.635000 ;
      RECT  6.395000  3.635000  8.245000 3.805000 ;
      RECT  6.665000  0.615000  6.995000 1.325000 ;
      RECT  6.745000  1.325000  6.915000 2.285000 ;
      RECT  6.745000  2.455000  6.915000 3.455000 ;
      RECT  7.095000  2.205000  7.425000 2.495000 ;
      RECT  7.095000  2.495000  7.265000 3.635000 ;
      RECT  7.175000  0.435000  7.345000 1.195000 ;
      RECT  7.175000  1.195000  7.445000 1.865000 ;
      RECT  7.445000  2.675000  7.795000 3.455000 ;
      RECT  7.540000  0.515000  8.595000 0.685000 ;
      RECT  7.540000  0.685000  7.795000 1.015000 ;
      RECT  7.625000  1.015000  7.795000 2.675000 ;
      RECT  7.975000  1.105000  8.245000 3.635000 ;
      RECT  8.425000  0.685000  8.595000 2.325000 ;
      RECT  8.425000  2.325000  9.725000 2.495000 ;
      RECT  8.505000  2.675000  9.455000 3.715000 ;
      RECT  8.775000  0.365000  9.725000 1.325000 ;
      RECT  8.775000  1.505000 10.235000 1.645000 ;
      RECT  8.775000  1.645000 10.505000 1.675000 ;
      RECT  8.775000  1.675000  9.105000 2.145000 ;
      RECT  9.395000  1.855000  9.725000 2.325000 ;
      RECT  9.905000  0.535000 10.235000 1.505000 ;
      RECT  9.905000  1.675000 10.505000 1.975000 ;
      RECT  9.905000  1.975000 10.235000 3.715000 ;
      RECT 11.070000  0.365000 11.625000 1.485000 ;
      RECT 11.070000  2.195000 11.605000 3.735000 ;
      RECT 11.785000  2.195000 12.115000 2.985000 ;
      RECT 11.805000  1.005000 12.135000 1.665000 ;
      RECT 11.805000  1.665000 13.300000 1.995000 ;
      RECT 11.805000  1.995000 12.115000 2.195000 ;
      RECT 12.295000  2.175000 13.245000 3.755000 ;
      RECT 12.315000  0.365000 13.265000 1.485000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.985000  0.325000 4.155000 ;
      RECT  0.600000  3.505000  0.770000 3.675000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.985000  0.805000 4.155000 ;
      RECT  0.650000  0.395000  0.820000 0.565000 ;
      RECT  0.960000  3.505000  1.130000 3.675000 ;
      RECT  1.010000  0.395000  1.180000 0.565000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.985000  1.285000 4.155000 ;
      RECT  1.370000  0.395000  1.540000 0.565000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.985000  1.765000 4.155000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.985000  2.245000 4.155000 ;
      RECT  2.100000  0.395000  2.270000 0.565000 ;
      RECT  2.460000  0.395000  2.630000 0.565000 ;
      RECT  2.470000  3.505000  2.640000 3.675000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.985000  2.725000 4.155000 ;
      RECT  2.820000  0.395000  2.990000 0.565000 ;
      RECT  2.830000  3.505000  3.000000 3.675000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.985000  3.205000 4.155000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.985000  3.685000 4.155000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.985000  4.165000 4.155000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.985000  4.645000 4.155000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.985000  5.125000 4.155000 ;
      RECT  5.215000  0.395000  5.385000 0.565000 ;
      RECT  5.295000  3.505000  5.465000 3.675000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.985000  5.605000 4.155000 ;
      RECT  5.575000  0.395000  5.745000 0.565000 ;
      RECT  5.655000  3.505000  5.825000 3.675000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.985000  6.085000 4.155000 ;
      RECT  5.935000  0.395000  6.105000 0.565000 ;
      RECT  6.015000  3.505000  6.185000 3.675000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.985000  6.565000 4.155000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.985000  7.045000 4.155000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.985000  7.525000 4.155000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.985000  8.005000 4.155000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.985000  8.485000 4.155000 ;
      RECT  8.535000  3.515000  8.705000 3.685000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.985000  8.965000 4.155000 ;
      RECT  8.805000  0.395000  8.975000 0.565000 ;
      RECT  8.895000  3.515000  9.065000 3.685000 ;
      RECT  9.165000  0.395000  9.335000 0.565000 ;
      RECT  9.255000  3.515000  9.425000 3.685000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.985000  9.445000 4.155000 ;
      RECT  9.525000  0.395000  9.695000 0.565000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.985000  9.925000 4.155000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.985000 10.405000 4.155000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.985000 10.885000 4.155000 ;
      RECT 11.070000  3.505000 11.240000 3.675000 ;
      RECT 11.080000  0.395000 11.250000 0.565000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.985000 11.365000 4.155000 ;
      RECT 11.430000  3.505000 11.600000 3.675000 ;
      RECT 11.440000  0.395000 11.610000 0.565000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.985000 11.845000 4.155000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.985000 12.325000 4.155000 ;
      RECT 12.325000  3.505000 12.495000 3.675000 ;
      RECT 12.345000  0.395000 12.515000 0.565000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.985000 12.805000 4.155000 ;
      RECT 12.685000  3.505000 12.855000 3.675000 ;
      RECT 12.705000  0.395000 12.875000 0.565000 ;
      RECT 13.045000  3.505000 13.215000 3.675000 ;
      RECT 13.065000  0.395000 13.235000 0.565000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.985000 13.285000 4.155000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.985000 13.765000 4.155000 ;
  END
END sky130_fd_sc_hvl__dfxbp_1
END LIBRARY