VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO raven_spi
  CLASS BLOCK ;
  FOREIGN raven_spi ;
  ORIGIN 0.000 0.000 ;
  SIZE 148.160 BY 169.200 ;
  PIN CSB
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 135.010 103.300 135.720 103.690 ;
      LAYER L1M1_PR_C ;
        RECT 135.510 103.330 135.680 103.500 ;
      LAYER met1 ;
        RECT 135.440 103.480 135.760 103.540 ;
        RECT 135.240 103.340 135.760 103.480 ;
        RECT 135.440 103.280 135.760 103.340 ;
      LAYER via ;
        RECT 135.470 103.280 135.730 103.540 ;
      LAYER met2 ;
        RECT 135.460 106.740 135.740 107.110 ;
        RECT 135.530 103.570 135.670 106.740 ;
        RECT 135.470 103.250 135.730 103.570 ;
      LAYER via2 ;
        RECT 135.460 106.790 135.740 107.070 ;
      LAYER met3 ;
        RECT 135.430 107.080 135.760 107.090 ;
        RECT 144.160 107.080 148.160 107.230 ;
        RECT 135.430 106.780 148.160 107.080 ;
        RECT 135.430 106.760 135.760 106.780 ;
        RECT 144.160 106.630 148.160 106.780 ;
    END
  END CSB
  PIN RST
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 11.170 119.580 11.880 119.970 ;
      LAYER L1M1_PR_C ;
        RECT 11.190 119.610 11.360 119.780 ;
      LAYER met1 ;
        RECT 11.120 119.760 11.440 119.820 ;
        RECT 10.920 119.620 11.440 119.760 ;
        RECT 11.120 119.560 11.440 119.620 ;
      LAYER via ;
        RECT 11.150 119.560 11.410 119.820 ;
      LAYER met2 ;
        RECT 11.150 119.530 11.410 119.850 ;
        RECT 11.210 117.470 11.350 119.530 ;
        RECT 11.140 117.100 11.420 117.470 ;
      LAYER via2 ;
        RECT 11.140 117.150 11.420 117.430 ;
      LAYER met3 ;
        RECT 0.000 117.440 4.000 117.590 ;
        RECT 11.110 117.440 11.440 117.450 ;
        RECT 0.000 117.140 11.440 117.440 ;
        RECT 0.000 116.990 4.000 117.140 ;
        RECT 11.110 117.120 11.440 117.140 ;
    END
  END RST
  PIN SCK
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 18.790 144.530 19.120 145.200 ;
        RECT 30.800 140.300 31.130 141.270 ;
        RECT 48.080 140.300 48.410 141.270 ;
        RECT 63.010 135.860 63.720 136.250 ;
        RECT 50.470 128.250 50.800 128.920 ;
        RECT 8.720 124.020 9.050 124.990 ;
        RECT 26.960 124.020 27.290 124.990 ;
        RECT 50.950 120.110 51.280 120.780 ;
        RECT 6.320 111.070 6.650 112.040 ;
        RECT 29.360 107.740 29.690 108.710 ;
        RECT 50.000 107.740 50.330 108.710 ;
        RECT 10.160 102.930 10.490 103.900 ;
        RECT 6.320 94.790 6.650 95.760 ;
        RECT 37.990 90.860 38.320 91.530 ;
        RECT 8.240 83.320 8.570 84.290 ;
        RECT 105.680 83.320 106.010 84.290 ;
        RECT 23.600 78.510 23.930 79.480 ;
        RECT 42.800 78.510 43.130 79.480 ;
        RECT 62.000 75.180 62.330 76.150 ;
        RECT 114.320 75.180 114.650 76.150 ;
        RECT 92.240 67.040 92.570 68.010 ;
        RECT 22.160 62.230 22.490 63.200 ;
        RECT 47.120 62.230 47.450 63.200 ;
        RECT 106.640 62.230 106.970 63.200 ;
        RECT 123.920 62.230 124.250 63.200 ;
        RECT 8.240 58.900 8.570 59.870 ;
        RECT 62.480 58.900 62.810 59.870 ;
        RECT 10.160 45.950 10.490 46.920 ;
        RECT 69.200 45.950 69.530 46.920 ;
        RECT 125.360 45.950 125.690 46.920 ;
        RECT 61.520 34.480 61.850 35.450 ;
        RECT 7.280 29.670 7.610 30.640 ;
        RECT 26.480 21.530 26.810 22.500 ;
        RECT 45.670 22.430 46.000 23.100 ;
        RECT 64.400 21.530 64.730 22.500 ;
        RECT 122.480 21.530 122.810 22.500 ;
        RECT 83.120 18.200 83.450 19.170 ;
        RECT 103.280 18.200 103.610 19.170 ;
      LAYER L1M1_PR_C ;
        RECT 18.870 144.770 19.040 144.940 ;
        RECT 30.870 140.330 31.040 140.500 ;
        RECT 48.150 140.330 48.320 140.500 ;
        RECT 63.030 135.890 63.200 136.060 ;
        RECT 50.550 128.490 50.720 128.660 ;
        RECT 8.790 124.790 8.960 124.960 ;
        RECT 27.030 124.790 27.200 124.960 ;
        RECT 51.030 120.350 51.200 120.520 ;
        RECT 6.390 111.840 6.560 112.010 ;
        RECT 29.430 108.510 29.600 108.680 ;
        RECT 50.070 108.510 50.240 108.680 ;
        RECT 10.230 103.700 10.400 103.870 ;
        RECT 6.390 95.560 6.560 95.730 ;
        RECT 38.070 91.120 38.240 91.290 ;
        RECT 8.310 84.090 8.480 84.260 ;
        RECT 105.750 83.350 105.920 83.520 ;
        RECT 23.670 78.540 23.840 78.710 ;
        RECT 42.870 78.540 43.040 78.710 ;
        RECT 62.070 75.210 62.240 75.380 ;
        RECT 114.390 75.210 114.560 75.380 ;
        RECT 92.310 67.070 92.480 67.240 ;
        RECT 22.230 62.260 22.400 62.430 ;
        RECT 47.190 63.000 47.360 63.170 ;
        RECT 106.710 62.630 106.880 62.800 ;
        RECT 123.990 62.260 124.160 62.430 ;
        RECT 8.310 58.930 8.480 59.100 ;
        RECT 62.550 58.930 62.720 59.100 ;
        RECT 10.230 45.980 10.400 46.150 ;
        RECT 69.270 45.980 69.440 46.150 ;
        RECT 125.430 45.980 125.600 46.150 ;
        RECT 61.590 35.250 61.760 35.420 ;
        RECT 7.350 30.440 7.520 30.610 ;
        RECT 45.750 22.670 45.920 22.840 ;
        RECT 26.550 22.300 26.720 22.470 ;
        RECT 64.470 21.560 64.640 21.730 ;
        RECT 122.550 21.560 122.720 21.730 ;
        RECT 83.190 18.600 83.360 18.770 ;
        RECT 103.350 18.600 103.520 18.770 ;
      LAYER met1 ;
        RECT 18.810 144.920 19.100 144.970 ;
        RECT 26.960 144.920 27.280 144.980 ;
        RECT 18.810 144.780 27.280 144.920 ;
        RECT 18.810 144.740 19.100 144.780 ;
        RECT 26.960 144.720 27.280 144.780 ;
        RECT 26.960 140.480 27.280 140.540 ;
        RECT 30.810 140.480 31.100 140.530 ;
        RECT 26.960 140.340 31.100 140.480 ;
        RECT 26.960 140.280 27.280 140.340 ;
        RECT 30.810 140.300 31.100 140.340 ;
        RECT 48.090 140.300 48.380 140.530 ;
        RECT 30.890 140.110 31.030 140.300 ;
        RECT 48.170 140.110 48.310 140.300 ;
        RECT 52.400 140.110 52.720 140.170 ;
        RECT 30.890 139.970 52.720 140.110 ;
        RECT 52.400 139.910 52.720 139.970 ;
        RECT 52.400 136.040 52.720 136.100 ;
        RECT 62.970 136.040 63.260 136.090 ;
        RECT 52.400 135.900 63.260 136.040 ;
        RECT 52.400 135.840 52.720 135.900 ;
        RECT 62.970 135.860 63.260 135.900 ;
        RECT 50.490 128.640 50.780 128.690 ;
        RECT 52.400 128.640 52.720 128.700 ;
        RECT 50.490 128.500 52.720 128.640 ;
        RECT 50.490 128.460 50.780 128.500 ;
        RECT 52.400 128.440 52.720 128.500 ;
        RECT 6.320 124.940 6.640 125.000 ;
        RECT 8.730 124.940 9.020 124.990 ;
        RECT 26.960 124.940 27.280 125.000 ;
        RECT 6.320 124.800 27.280 124.940 ;
        RECT 6.320 124.740 6.640 124.800 ;
        RECT 8.730 124.760 9.020 124.800 ;
        RECT 26.960 124.740 27.280 124.800 ;
        RECT 50.970 120.500 51.260 120.550 ;
        RECT 52.400 120.500 52.720 120.560 ;
        RECT 50.970 120.360 52.720 120.500 ;
        RECT 50.970 120.320 51.260 120.360 ;
        RECT 52.400 120.300 52.720 120.360 ;
        RECT 6.320 111.990 6.640 112.050 ;
        RECT 6.120 111.850 6.640 111.990 ;
        RECT 6.320 111.790 6.640 111.850 ;
        RECT 29.370 108.660 29.660 108.710 ;
        RECT 50.010 108.660 50.300 108.710 ;
        RECT 29.370 108.520 50.300 108.660 ;
        RECT 29.370 108.480 29.660 108.520 ;
        RECT 50.010 108.480 50.300 108.520 ;
        RECT 6.320 107.180 6.640 107.240 ;
        RECT 29.450 107.180 29.590 108.480 ;
        RECT 6.320 107.040 29.590 107.180 ;
        RECT 6.320 106.980 6.640 107.040 ;
        RECT 6.320 103.850 6.640 103.910 ;
        RECT 10.170 103.850 10.460 103.900 ;
        RECT 6.320 103.710 10.460 103.850 ;
        RECT 6.320 103.650 6.640 103.710 ;
        RECT 10.170 103.670 10.460 103.710 ;
        RECT 6.320 95.710 6.640 95.770 ;
        RECT 6.120 95.570 6.640 95.710 ;
        RECT 6.320 95.510 6.640 95.570 ;
        RECT 38.010 91.270 38.300 91.320 ;
        RECT 42.320 91.270 42.640 91.330 ;
        RECT 38.010 91.130 42.640 91.270 ;
        RECT 38.010 91.090 38.300 91.130 ;
        RECT 42.320 91.070 42.640 91.130 ;
        RECT 6.320 84.240 6.640 84.300 ;
        RECT 8.250 84.240 8.540 84.290 ;
        RECT 6.320 84.100 8.540 84.240 ;
        RECT 6.320 84.040 6.640 84.100 ;
        RECT 8.250 84.060 8.540 84.100 ;
        RECT 8.330 83.870 8.470 84.060 ;
        RECT 23.600 83.870 23.920 83.930 ;
        RECT 8.330 83.730 23.920 83.870 ;
        RECT 23.600 83.670 23.920 83.730 ;
        RECT 105.690 83.500 105.980 83.550 ;
        RECT 106.640 83.500 106.960 83.560 ;
        RECT 105.690 83.360 106.960 83.500 ;
        RECT 105.690 83.320 105.980 83.360 ;
        RECT 106.640 83.300 106.960 83.360 ;
        RECT 23.600 78.690 23.920 78.750 ;
        RECT 23.400 78.550 23.920 78.690 ;
        RECT 23.600 78.490 23.920 78.550 ;
        RECT 42.320 78.690 42.640 78.750 ;
        RECT 42.810 78.690 43.100 78.740 ;
        RECT 42.320 78.550 43.100 78.690 ;
        RECT 42.320 78.490 42.640 78.550 ;
        RECT 42.810 78.510 43.100 78.550 ;
        RECT 62.000 75.360 62.320 75.420 ;
        RECT 61.800 75.220 62.320 75.360 ;
        RECT 62.000 75.160 62.320 75.220 ;
        RECT 106.640 75.360 106.960 75.420 ;
        RECT 107.600 75.360 107.920 75.420 ;
        RECT 114.330 75.360 114.620 75.410 ;
        RECT 106.640 75.220 114.620 75.360 ;
        RECT 106.640 75.160 106.960 75.220 ;
        RECT 107.600 75.160 107.920 75.220 ;
        RECT 114.330 75.180 114.620 75.220 ;
        RECT 23.600 74.250 23.920 74.310 ;
        RECT 42.320 74.250 42.640 74.310 ;
        RECT 23.600 74.110 42.640 74.250 ;
        RECT 23.600 74.050 23.920 74.110 ;
        RECT 42.320 74.050 42.640 74.110 ;
        RECT 42.320 72.400 42.640 72.460 ;
        RECT 62.000 72.400 62.320 72.460 ;
        RECT 42.320 72.260 62.320 72.400 ;
        RECT 42.320 72.200 42.640 72.260 ;
        RECT 62.000 72.200 62.320 72.260 ;
        RECT 92.240 67.220 92.560 67.280 ;
        RECT 92.040 67.080 92.560 67.220 ;
        RECT 92.240 67.020 92.560 67.080 ;
        RECT 42.320 63.520 42.640 63.580 ;
        RECT 42.320 63.380 47.350 63.520 ;
        RECT 42.320 63.320 42.640 63.380 ;
        RECT 47.210 63.200 47.350 63.380 ;
        RECT 47.130 62.970 47.420 63.200 ;
        RECT 106.650 62.780 106.940 62.830 ;
        RECT 107.600 62.780 107.920 62.840 ;
        RECT 106.650 62.640 124.150 62.780 ;
        RECT 106.650 62.600 106.940 62.640 ;
        RECT 107.600 62.580 107.920 62.640 ;
        RECT 22.160 62.410 22.480 62.470 ;
        RECT 23.600 62.410 23.920 62.470 ;
        RECT 124.010 62.460 124.150 62.640 ;
        RECT 21.960 62.270 23.920 62.410 ;
        RECT 22.160 62.210 22.480 62.270 ;
        RECT 23.600 62.210 23.920 62.270 ;
        RECT 123.930 62.410 124.220 62.460 ;
        RECT 125.840 62.410 126.160 62.470 ;
        RECT 123.930 62.270 126.160 62.410 ;
        RECT 123.930 62.230 124.220 62.270 ;
        RECT 125.840 62.210 126.160 62.270 ;
        RECT 8.250 58.900 8.540 59.130 ;
        RECT 62.000 59.080 62.320 59.140 ;
        RECT 62.490 59.080 62.780 59.130 ;
        RECT 62.000 58.940 62.780 59.080 ;
        RECT 8.330 57.970 8.470 58.900 ;
        RECT 62.000 58.880 62.320 58.940 ;
        RECT 62.490 58.900 62.780 58.940 ;
        RECT 22.160 57.970 22.480 58.030 ;
        RECT 8.330 57.830 22.480 57.970 ;
        RECT 22.160 57.770 22.480 57.830 ;
        RECT 92.240 46.500 92.560 46.560 ;
        RECT 69.290 46.360 92.560 46.500 ;
        RECT 7.280 46.130 7.600 46.190 ;
        RECT 69.290 46.180 69.430 46.360 ;
        RECT 92.240 46.300 92.560 46.360 ;
        RECT 10.170 46.130 10.460 46.180 ;
        RECT 7.280 45.990 10.460 46.130 ;
        RECT 7.280 45.930 7.600 45.990 ;
        RECT 10.170 45.950 10.460 45.990 ;
        RECT 69.210 45.950 69.500 46.180 ;
        RECT 125.370 46.130 125.660 46.180 ;
        RECT 125.840 46.130 126.160 46.190 ;
        RECT 125.370 45.990 126.160 46.130 ;
        RECT 125.370 45.950 125.660 45.990 ;
        RECT 62.000 45.760 62.320 45.820 ;
        RECT 69.290 45.760 69.430 45.950 ;
        RECT 125.840 45.930 126.160 45.990 ;
        RECT 62.000 45.620 69.430 45.760 ;
        RECT 62.000 45.560 62.320 45.620 ;
        RECT 61.530 35.220 61.820 35.450 ;
        RECT 61.610 35.030 61.750 35.220 ;
        RECT 62.000 35.030 62.320 35.090 ;
        RECT 61.610 34.890 62.320 35.030 ;
        RECT 62.000 34.830 62.320 34.890 ;
        RECT 7.280 30.590 7.600 30.650 ;
        RECT 7.080 30.450 7.600 30.590 ;
        RECT 7.280 30.390 7.600 30.450 ;
        RECT 45.690 22.820 45.980 22.870 ;
        RECT 43.850 22.680 45.980 22.820 ;
        RECT 7.280 22.450 7.600 22.510 ;
        RECT 26.490 22.450 26.780 22.500 ;
        RECT 7.280 22.310 26.780 22.450 ;
        RECT 7.280 22.250 7.600 22.310 ;
        RECT 26.490 22.270 26.780 22.310 ;
        RECT 26.570 21.710 26.710 22.270 ;
        RECT 43.850 21.710 43.990 22.680 ;
        RECT 45.690 22.640 45.980 22.680 ;
        RECT 45.770 22.450 45.910 22.640 ;
        RECT 62.000 22.450 62.320 22.510 ;
        RECT 45.770 22.310 64.150 22.450 ;
        RECT 62.000 22.250 62.320 22.310 ;
        RECT 26.570 21.570 43.990 21.710 ;
        RECT 64.010 21.710 64.150 22.310 ;
        RECT 64.410 21.710 64.700 21.760 ;
        RECT 83.120 21.710 83.440 21.770 ;
        RECT 122.490 21.710 122.780 21.760 ;
        RECT 125.840 21.710 126.160 21.770 ;
        RECT 64.010 21.570 83.440 21.710 ;
        RECT 64.410 21.530 64.700 21.570 ;
        RECT 83.120 21.510 83.440 21.570 ;
        RECT 107.690 21.570 126.160 21.710 ;
        RECT 103.280 21.340 103.600 21.400 ;
        RECT 107.690 21.340 107.830 21.570 ;
        RECT 122.490 21.530 122.780 21.570 ;
        RECT 125.840 21.510 126.160 21.570 ;
        RECT 103.280 21.200 107.830 21.340 ;
        RECT 103.280 21.140 103.600 21.200 ;
        RECT 83.120 18.750 83.440 18.810 ;
        RECT 103.280 18.750 103.600 18.810 ;
        RECT 82.680 18.610 103.600 18.750 ;
        RECT 83.120 18.550 83.440 18.610 ;
        RECT 103.280 18.550 103.600 18.610 ;
      LAYER via ;
        RECT 26.990 144.720 27.250 144.980 ;
        RECT 26.990 140.280 27.250 140.540 ;
        RECT 52.430 139.910 52.690 140.170 ;
        RECT 52.430 135.840 52.690 136.100 ;
        RECT 52.430 128.440 52.690 128.700 ;
        RECT 6.350 124.740 6.610 125.000 ;
        RECT 26.990 124.740 27.250 125.000 ;
        RECT 52.430 120.300 52.690 120.560 ;
        RECT 6.350 111.790 6.610 112.050 ;
        RECT 6.350 106.980 6.610 107.240 ;
        RECT 6.350 103.650 6.610 103.910 ;
        RECT 6.350 95.510 6.610 95.770 ;
        RECT 42.350 91.070 42.610 91.330 ;
        RECT 6.350 84.040 6.610 84.300 ;
        RECT 23.630 83.670 23.890 83.930 ;
        RECT 106.670 83.300 106.930 83.560 ;
        RECT 23.630 78.490 23.890 78.750 ;
        RECT 42.350 78.490 42.610 78.750 ;
        RECT 62.030 75.160 62.290 75.420 ;
        RECT 106.670 75.160 106.930 75.420 ;
        RECT 107.630 75.160 107.890 75.420 ;
        RECT 23.630 74.050 23.890 74.310 ;
        RECT 42.350 74.050 42.610 74.310 ;
        RECT 42.350 72.200 42.610 72.460 ;
        RECT 62.030 72.200 62.290 72.460 ;
        RECT 92.270 67.020 92.530 67.280 ;
        RECT 42.350 63.320 42.610 63.580 ;
        RECT 107.630 62.580 107.890 62.840 ;
        RECT 22.190 62.210 22.450 62.470 ;
        RECT 23.630 62.210 23.890 62.470 ;
        RECT 125.870 62.210 126.130 62.470 ;
        RECT 62.030 58.880 62.290 59.140 ;
        RECT 22.190 57.770 22.450 58.030 ;
        RECT 7.310 45.930 7.570 46.190 ;
        RECT 92.270 46.300 92.530 46.560 ;
        RECT 62.030 45.560 62.290 45.820 ;
        RECT 125.870 45.930 126.130 46.190 ;
        RECT 62.030 34.830 62.290 35.090 ;
        RECT 7.310 30.390 7.570 30.650 ;
        RECT 7.310 22.250 7.570 22.510 ;
        RECT 62.030 22.250 62.290 22.510 ;
        RECT 83.150 21.510 83.410 21.770 ;
        RECT 103.310 21.140 103.570 21.400 ;
        RECT 125.870 21.510 126.130 21.770 ;
        RECT 83.150 18.550 83.410 18.810 ;
        RECT 103.310 18.550 103.570 18.810 ;
      LAYER met2 ;
        RECT 26.990 144.690 27.250 145.010 ;
        RECT 27.050 140.570 27.190 144.690 ;
        RECT 26.990 140.250 27.250 140.570 ;
        RECT 27.050 125.030 27.190 140.250 ;
        RECT 52.430 139.880 52.690 140.200 ;
        RECT 52.490 136.130 52.630 139.880 ;
        RECT 52.430 135.810 52.690 136.130 ;
        RECT 52.490 128.730 52.630 135.810 ;
        RECT 52.430 128.410 52.690 128.730 ;
        RECT 6.350 124.710 6.610 125.030 ;
        RECT 26.990 124.710 27.250 125.030 ;
        RECT 6.410 112.080 6.550 124.710 ;
        RECT 52.490 120.590 52.630 128.410 ;
        RECT 52.430 120.270 52.690 120.590 ;
        RECT 6.350 111.760 6.610 112.080 ;
        RECT 6.410 107.270 6.550 111.760 ;
        RECT 6.350 106.950 6.610 107.270 ;
        RECT 6.410 103.940 6.550 106.950 ;
        RECT 6.350 103.620 6.610 103.940 ;
        RECT 6.410 95.800 6.550 103.620 ;
        RECT 6.350 95.480 6.610 95.800 ;
        RECT 6.410 84.910 6.550 95.480 ;
        RECT 42.350 91.040 42.610 91.360 ;
        RECT 6.340 84.540 6.620 84.910 ;
        RECT 6.410 84.330 6.550 84.540 ;
        RECT 6.350 84.010 6.610 84.330 ;
        RECT 23.630 83.640 23.890 83.960 ;
        RECT 23.690 78.780 23.830 83.640 ;
        RECT 42.410 78.780 42.550 91.040 ;
        RECT 106.670 83.270 106.930 83.590 ;
        RECT 23.630 78.460 23.890 78.780 ;
        RECT 42.350 78.460 42.610 78.780 ;
        RECT 23.690 74.340 23.830 78.460 ;
        RECT 42.410 74.340 42.550 78.460 ;
        RECT 106.730 75.450 106.870 83.270 ;
        RECT 62.030 75.130 62.290 75.450 ;
        RECT 106.670 75.130 106.930 75.450 ;
        RECT 107.630 75.130 107.890 75.450 ;
        RECT 23.630 74.020 23.890 74.340 ;
        RECT 42.350 74.020 42.610 74.340 ;
        RECT 23.690 62.500 23.830 74.020 ;
        RECT 42.410 72.490 42.550 74.020 ;
        RECT 62.090 72.490 62.230 75.130 ;
        RECT 42.350 72.170 42.610 72.490 ;
        RECT 62.030 72.170 62.290 72.490 ;
        RECT 42.410 63.610 42.550 72.170 ;
        RECT 42.350 63.290 42.610 63.610 ;
        RECT 22.190 62.180 22.450 62.500 ;
        RECT 23.630 62.180 23.890 62.500 ;
        RECT 22.250 58.060 22.390 62.180 ;
        RECT 62.090 59.170 62.230 72.170 ;
        RECT 92.270 66.990 92.530 67.310 ;
        RECT 62.030 58.850 62.290 59.170 ;
        RECT 22.190 57.740 22.450 58.060 ;
        RECT 7.310 45.900 7.570 46.220 ;
        RECT 7.370 30.680 7.510 45.900 ;
        RECT 62.090 45.850 62.230 58.850 ;
        RECT 92.330 46.590 92.470 66.990 ;
        RECT 107.690 62.870 107.830 75.130 ;
        RECT 107.630 62.550 107.890 62.870 ;
        RECT 125.870 62.180 126.130 62.500 ;
        RECT 92.270 46.270 92.530 46.590 ;
        RECT 125.930 46.220 126.070 62.180 ;
        RECT 125.870 45.900 126.130 46.220 ;
        RECT 62.030 45.530 62.290 45.850 ;
        RECT 62.090 35.120 62.230 45.530 ;
        RECT 62.030 34.800 62.290 35.120 ;
        RECT 7.310 30.360 7.570 30.680 ;
        RECT 7.370 22.540 7.510 30.360 ;
        RECT 62.090 22.540 62.230 34.800 ;
        RECT 7.310 22.220 7.570 22.540 ;
        RECT 62.030 22.220 62.290 22.540 ;
        RECT 125.930 21.800 126.070 45.900 ;
        RECT 83.150 21.480 83.410 21.800 ;
        RECT 125.870 21.480 126.130 21.800 ;
        RECT 83.210 18.840 83.350 21.480 ;
        RECT 103.310 21.110 103.570 21.430 ;
        RECT 103.370 18.840 103.510 21.110 ;
        RECT 83.150 18.520 83.410 18.840 ;
        RECT 103.310 18.520 103.570 18.840 ;
      LAYER via2 ;
        RECT 6.340 84.590 6.620 84.870 ;
      LAYER met3 ;
        RECT 0.000 84.880 4.000 85.030 ;
        RECT 6.310 84.880 6.640 84.890 ;
        RECT 0.000 84.580 6.640 84.880 ;
        RECT 0.000 84.430 4.000 84.580 ;
        RECT 6.310 84.560 6.640 84.580 ;
    END
  END SCK
  PIN SDI
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 92.290 54.720 93.000 55.030 ;
        RECT 8.290 50.970 9.000 51.360 ;
        RECT 73.470 17.090 73.800 18.880 ;
      LAYER L1M1_PR_C ;
        RECT 92.790 54.860 92.960 55.030 ;
        RECT 8.790 51.160 8.960 51.330 ;
        RECT 73.590 18.600 73.760 18.770 ;
      LAYER met1 ;
        RECT 92.720 55.010 93.040 55.070 ;
        RECT 92.520 54.870 93.040 55.010 ;
        RECT 92.720 54.810 93.040 54.870 ;
        RECT 8.730 51.130 9.020 51.360 ;
        RECT 8.810 50.940 8.950 51.130 ;
        RECT 14.480 50.940 14.800 51.000 ;
        RECT 19.760 50.940 20.080 51.000 ;
        RECT 8.810 50.800 20.080 50.940 ;
        RECT 14.480 50.740 14.800 50.800 ;
        RECT 19.760 50.740 20.080 50.800 ;
        RECT 49.040 49.830 49.360 49.890 ;
        RECT 75.440 49.830 75.760 49.890 ;
        RECT 92.720 49.830 93.040 49.890 ;
        RECT 49.040 49.690 93.040 49.830 ;
        RECT 49.040 49.630 49.360 49.690 ;
        RECT 75.440 49.630 75.760 49.690 ;
        RECT 92.720 49.630 93.040 49.690 ;
        RECT 19.760 47.610 20.080 47.670 ;
        RECT 19.760 47.470 35.830 47.610 ;
        RECT 19.760 47.410 20.080 47.470 ;
        RECT 35.690 47.240 35.830 47.470 ;
        RECT 49.040 47.240 49.360 47.300 ;
        RECT 35.690 47.100 49.360 47.240 ;
        RECT 49.040 47.040 49.360 47.100 ;
        RECT 73.530 18.750 73.820 18.800 ;
        RECT 75.440 18.750 75.760 18.810 ;
        RECT 73.530 18.610 75.760 18.750 ;
        RECT 73.530 18.570 73.820 18.610 ;
        RECT 75.440 18.550 75.760 18.610 ;
      LAYER via ;
        RECT 92.750 54.810 93.010 55.070 ;
        RECT 14.510 50.740 14.770 51.000 ;
        RECT 19.790 50.740 20.050 51.000 ;
        RECT 49.070 49.630 49.330 49.890 ;
        RECT 75.470 49.630 75.730 49.890 ;
        RECT 92.750 49.630 93.010 49.890 ;
        RECT 19.790 47.410 20.050 47.670 ;
        RECT 49.070 47.040 49.330 47.300 ;
        RECT 75.470 18.550 75.730 18.810 ;
      LAYER met2 ;
        RECT 92.750 54.780 93.010 55.100 ;
        RECT 14.510 50.710 14.770 51.030 ;
        RECT 19.790 50.710 20.050 51.030 ;
        RECT 14.570 36.070 14.710 50.710 ;
        RECT 19.850 47.700 19.990 50.710 ;
        RECT 92.810 49.920 92.950 54.780 ;
        RECT 49.070 49.600 49.330 49.920 ;
        RECT 75.470 49.600 75.730 49.920 ;
        RECT 92.750 49.600 93.010 49.920 ;
        RECT 19.790 47.380 20.050 47.700 ;
        RECT 49.130 47.330 49.270 49.600 ;
        RECT 49.070 47.010 49.330 47.330 ;
        RECT 14.500 35.700 14.780 36.070 ;
        RECT 75.530 18.840 75.670 49.600 ;
        RECT 75.470 18.520 75.730 18.840 ;
      LAYER via2 ;
        RECT 14.500 35.750 14.780 36.030 ;
      LAYER met3 ;
        RECT 0.000 36.040 4.000 36.190 ;
        RECT 14.470 36.040 14.800 36.050 ;
        RECT 0.000 35.740 14.800 36.040 ;
        RECT 0.000 35.590 4.000 35.740 ;
        RECT 14.470 35.720 14.800 35.740 ;
    END
  END SDI
  PIN SDO
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 75.380 143.120 75.720 146.190 ;
        RECT 81.650 144.230 81.980 144.570 ;
      LAYER L1M1_PR_C ;
        RECT 75.510 144.770 75.680 144.940 ;
        RECT 81.750 144.400 81.920 144.570 ;
      LAYER met1 ;
        RECT 34.640 144.920 34.960 144.980 ;
        RECT 75.450 144.920 75.740 144.970 ;
        RECT 34.640 144.780 75.740 144.920 ;
        RECT 34.640 144.720 34.960 144.780 ;
        RECT 75.450 144.740 75.740 144.780 ;
        RECT 75.530 144.550 75.670 144.740 ;
        RECT 81.690 144.550 81.980 144.600 ;
        RECT 75.530 144.410 81.980 144.550 ;
        RECT 81.690 144.370 81.980 144.410 ;
      LAYER via ;
        RECT 34.670 144.720 34.930 144.980 ;
      LAYER met2 ;
        RECT 34.660 165.200 34.940 169.200 ;
        RECT 34.730 145.010 34.870 165.200 ;
        RECT 34.670 144.690 34.930 145.010 ;
    END
  END SDO
  PIN irq
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 104.850 87.040 105.450 87.430 ;
        RECT 120.020 81.730 120.360 84.800 ;
        RECT 95.650 70.740 96.360 71.130 ;
      LAYER L1M1_PR_C ;
        RECT 105.270 87.050 105.440 87.220 ;
        RECT 120.150 82.240 120.320 82.410 ;
        RECT 95.670 70.770 95.840 70.940 ;
      LAYER met1 ;
        RECT 105.210 87.200 105.500 87.250 ;
        RECT 104.330 87.060 105.500 87.200 ;
        RECT 100.880 86.830 101.200 86.890 ;
        RECT 104.330 86.830 104.470 87.060 ;
        RECT 105.210 87.020 105.500 87.060 ;
        RECT 100.880 86.690 104.470 86.830 ;
        RECT 100.880 86.630 101.200 86.690 ;
        RECT 100.880 82.390 101.200 82.450 ;
        RECT 120.090 82.390 120.380 82.440 ;
        RECT 100.880 82.250 120.380 82.390 ;
        RECT 100.880 82.190 101.200 82.250 ;
        RECT 120.090 82.210 120.380 82.250 ;
        RECT 98.480 71.290 98.800 71.350 ;
        RECT 95.690 71.150 98.800 71.290 ;
        RECT 93.680 70.920 94.000 70.980 ;
        RECT 95.690 70.970 95.830 71.150 ;
        RECT 98.480 71.090 98.800 71.150 ;
        RECT 95.610 70.920 95.900 70.970 ;
        RECT 93.680 70.780 95.900 70.920 ;
        RECT 93.680 70.720 94.000 70.780 ;
        RECT 95.610 70.740 95.900 70.780 ;
        RECT 93.200 18.380 93.520 18.440 ;
        RECT 97.040 18.380 97.360 18.440 ;
        RECT 93.200 18.240 97.360 18.380 ;
        RECT 93.200 18.180 93.520 18.240 ;
        RECT 97.040 18.180 97.360 18.240 ;
      LAYER via ;
        RECT 100.910 86.630 101.170 86.890 ;
        RECT 100.910 82.190 101.170 82.450 ;
        RECT 93.710 70.720 93.970 70.980 ;
        RECT 98.510 71.090 98.770 71.350 ;
        RECT 93.230 18.180 93.490 18.440 ;
        RECT 97.070 18.180 97.330 18.440 ;
      LAYER met2 ;
        RECT 100.910 86.600 101.170 86.920 ;
        RECT 100.970 82.480 101.110 86.600 ;
        RECT 100.910 82.160 101.170 82.480 ;
        RECT 98.510 71.290 98.770 71.380 ;
        RECT 100.970 71.290 101.110 82.160 ;
        RECT 98.510 71.150 101.110 71.290 ;
        RECT 98.510 71.060 98.770 71.150 ;
        RECT 93.710 70.690 93.970 71.010 ;
        RECT 93.770 50.200 93.910 70.690 ;
        RECT 93.290 50.060 93.910 50.200 ;
        RECT 93.290 18.470 93.430 50.060 ;
        RECT 93.230 18.150 93.490 18.470 ;
        RECT 97.070 18.150 97.330 18.470 ;
        RECT 97.130 4.000 97.270 18.150 ;
        RECT 97.060 0.000 97.340 4.000 ;
    END
  END irq
  PIN mask_rev[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 128.280 95.790 128.710 97.370 ;
        RECT 128.280 94.110 128.530 95.790 ;
      LAYER L1M1_PR_C ;
        RECT 128.310 94.450 128.480 94.620 ;
      LAYER met1 ;
        RECT 122.000 94.600 122.320 94.660 ;
        RECT 128.250 94.600 128.540 94.650 ;
        RECT 122.000 94.460 128.540 94.600 ;
        RECT 122.000 94.400 122.320 94.460 ;
        RECT 128.250 94.420 128.540 94.460 ;
        RECT 117.200 21.340 117.520 21.400 ;
        RECT 122.000 21.340 122.320 21.400 ;
        RECT 117.200 21.200 122.320 21.340 ;
        RECT 117.200 21.140 117.520 21.200 ;
        RECT 122.000 21.140 122.320 21.200 ;
      LAYER via ;
        RECT 122.030 94.400 122.290 94.660 ;
        RECT 117.230 21.140 117.490 21.400 ;
        RECT 122.030 21.140 122.290 21.400 ;
      LAYER met2 ;
        RECT 122.030 94.370 122.290 94.690 ;
        RECT 122.090 21.430 122.230 94.370 ;
        RECT 117.230 21.110 117.490 21.430 ;
        RECT 122.030 21.110 122.290 21.430 ;
        RECT 117.290 4.000 117.430 21.110 ;
        RECT 117.220 0.000 117.500 4.000 ;
    END
  END mask_rev[0]
  PIN mask_rev[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 12.600 136.490 13.030 138.070 ;
        RECT 12.600 134.810 12.850 136.490 ;
      LAYER L1M1_PR_C ;
        RECT 12.630 136.630 12.800 136.800 ;
      LAYER met1 ;
        RECT 7.280 151.210 7.600 151.270 ;
        RECT 13.520 151.210 13.840 151.270 ;
        RECT 7.280 151.070 13.840 151.210 ;
        RECT 7.280 151.010 7.600 151.070 ;
        RECT 13.520 151.010 13.840 151.070 ;
        RECT 7.280 136.780 7.600 136.840 ;
        RECT 12.570 136.780 12.860 136.830 ;
        RECT 7.280 136.640 12.860 136.780 ;
        RECT 7.280 136.580 7.600 136.640 ;
        RECT 12.570 136.600 12.860 136.640 ;
      LAYER via ;
        RECT 7.310 151.010 7.570 151.270 ;
        RECT 13.550 151.010 13.810 151.270 ;
        RECT 7.310 136.580 7.570 136.840 ;
      LAYER met2 ;
        RECT 13.540 165.200 13.820 169.200 ;
        RECT 13.610 151.300 13.750 165.200 ;
        RECT 7.310 150.980 7.570 151.300 ;
        RECT 13.550 150.980 13.810 151.300 ;
        RECT 7.370 136.870 7.510 150.980 ;
        RECT 7.310 136.550 7.570 136.870 ;
    END
  END mask_rev[1]
  PIN mask_rev[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 133.560 144.630 133.990 146.210 ;
        RECT 133.560 142.950 133.810 144.630 ;
      LAYER L1M1_PR_C ;
        RECT 133.590 145.510 133.760 145.680 ;
      LAYER met1 ;
        RECT 133.530 145.660 133.820 145.710 ;
        RECT 139.280 145.660 139.600 145.720 ;
        RECT 133.530 145.520 139.600 145.660 ;
        RECT 133.530 145.480 133.820 145.520 ;
        RECT 139.280 145.460 139.600 145.520 ;
      LAYER via ;
        RECT 139.310 145.460 139.570 145.720 ;
      LAYER met2 ;
        RECT 139.300 165.200 139.580 169.200 ;
        RECT 139.370 145.750 139.510 165.200 ;
        RECT 139.310 145.430 139.570 145.750 ;
    END
  END mask_rev[2]
  PIN mask_rev[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 102.360 144.630 102.790 146.210 ;
        RECT 102.360 142.950 102.610 144.630 ;
      LAYER L1M1_PR_C ;
        RECT 102.390 145.510 102.560 145.680 ;
      LAYER met1 ;
        RECT 102.330 145.660 102.620 145.710 ;
        RECT 107.600 145.660 107.920 145.720 ;
        RECT 102.330 145.520 107.920 145.660 ;
        RECT 102.330 145.480 102.620 145.520 ;
        RECT 107.600 145.460 107.920 145.520 ;
      LAYER via ;
        RECT 107.630 145.460 107.890 145.720 ;
      LAYER met2 ;
        RECT 107.620 165.200 107.900 169.200 ;
        RECT 107.690 145.750 107.830 165.200 ;
        RECT 107.630 145.430 107.890 145.750 ;
    END
  END mask_rev[3]
  PIN mask_rev_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 100.730 103.500 101.160 103.870 ;
        RECT 129.630 95.080 129.960 96.870 ;
      LAYER L1M1_PR_C ;
        RECT 100.950 103.700 101.120 103.870 ;
        RECT 129.750 96.670 129.920 96.840 ;
      LAYER met1 ;
        RECT 100.890 103.670 101.180 103.900 ;
        RECT 100.970 102.740 101.110 103.670 ;
        RECT 129.680 102.740 130.000 102.800 ;
        RECT 100.970 102.600 130.000 102.740 ;
        RECT 129.680 102.540 130.000 102.600 ;
        RECT 129.680 96.820 130.000 96.880 ;
        RECT 129.480 96.680 130.000 96.820 ;
        RECT 129.680 96.620 130.000 96.680 ;
      LAYER via ;
        RECT 129.710 102.540 129.970 102.800 ;
        RECT 129.710 96.620 129.970 96.880 ;
      LAYER met2 ;
        RECT 129.220 139.300 129.500 139.670 ;
        RECT 129.290 104.040 129.430 139.300 ;
        RECT 129.290 103.900 129.910 104.040 ;
        RECT 129.770 102.830 129.910 103.900 ;
        RECT 129.710 102.510 129.970 102.830 ;
        RECT 129.770 96.910 129.910 102.510 ;
        RECT 129.710 96.590 129.970 96.910 ;
      LAYER via2 ;
        RECT 129.220 139.350 129.500 139.630 ;
      LAYER met3 ;
        RECT 129.190 139.640 129.520 139.650 ;
        RECT 144.160 139.640 148.160 139.790 ;
        RECT 129.190 139.340 148.160 139.640 ;
        RECT 129.190 139.320 129.520 139.340 ;
        RECT 144.160 139.190 148.160 139.340 ;
    END
  END mask_rev_in[0]
  PIN mask_rev_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 13.950 135.780 14.280 137.570 ;
        RECT 77.210 127.680 78.120 128.010 ;
      LAYER L1M1_PR_C ;
        RECT 14.070 135.890 14.240 136.060 ;
        RECT 77.430 127.750 77.600 127.920 ;
      LAYER met1 ;
        RECT 14.010 136.040 14.300 136.090 ;
        RECT 20.240 136.040 20.560 136.100 ;
        RECT 14.010 135.900 20.560 136.040 ;
        RECT 14.010 135.860 14.300 135.900 ;
        RECT 20.240 135.840 20.560 135.900 ;
        RECT 18.320 129.010 18.640 129.070 ;
        RECT 20.240 129.010 20.560 129.070 ;
        RECT 18.320 128.870 77.590 129.010 ;
        RECT 18.320 128.810 18.640 128.870 ;
        RECT 20.240 128.810 20.560 128.870 ;
        RECT 77.450 127.950 77.590 128.870 ;
        RECT 77.370 127.720 77.660 127.950 ;
      LAYER via ;
        RECT 20.270 135.840 20.530 136.100 ;
        RECT 18.350 128.810 18.610 129.070 ;
        RECT 20.270 128.810 20.530 129.070 ;
      LAYER met2 ;
        RECT 20.270 135.810 20.530 136.130 ;
        RECT 20.330 129.100 20.470 135.810 ;
        RECT 18.350 128.780 18.610 129.100 ;
        RECT 20.270 128.780 20.530 129.100 ;
        RECT 18.410 68.630 18.550 128.780 ;
        RECT 18.340 68.260 18.620 68.630 ;
      LAYER via2 ;
        RECT 18.340 68.310 18.620 68.590 ;
      LAYER met3 ;
        RECT 0.000 68.600 4.000 68.750 ;
        RECT 18.310 68.600 18.640 68.610 ;
        RECT 0.000 68.300 18.640 68.600 ;
        RECT 0.000 68.150 4.000 68.300 ;
        RECT 18.310 68.280 18.640 68.300 ;
    END
  END mask_rev_in[1]
  PIN mask_rev_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 134.910 143.920 135.240 145.710 ;
        RECT 102.170 99.630 102.600 100.000 ;
      LAYER L1M1_PR_C ;
        RECT 135.030 144.030 135.200 144.200 ;
        RECT 102.390 99.630 102.560 99.800 ;
      LAYER met1 ;
        RECT 134.960 144.180 135.280 144.240 ;
        RECT 134.760 144.040 135.280 144.180 ;
        RECT 134.960 143.980 135.280 144.040 ;
        RECT 102.330 99.780 102.620 99.830 ;
        RECT 102.330 99.640 123.670 99.780 ;
        RECT 102.330 99.600 102.620 99.640 ;
        RECT 123.530 99.470 123.670 99.640 ;
        RECT 123.440 99.410 123.760 99.470 ;
        RECT 134.960 99.410 135.280 99.470 ;
        RECT 123.000 99.270 135.280 99.410 ;
        RECT 123.440 99.210 123.760 99.270 ;
        RECT 134.960 99.210 135.280 99.270 ;
      LAYER via ;
        RECT 134.990 143.980 135.250 144.240 ;
        RECT 123.470 99.210 123.730 99.470 ;
        RECT 134.990 99.210 135.250 99.470 ;
      LAYER met2 ;
        RECT 134.990 143.950 135.250 144.270 ;
        RECT 135.050 99.500 135.190 143.950 ;
        RECT 123.470 99.180 123.730 99.500 ;
        RECT 134.990 99.180 135.250 99.500 ;
        RECT 123.530 91.460 123.670 99.180 ;
        RECT 123.530 91.320 124.150 91.460 ;
        RECT 124.010 21.160 124.150 91.320 ;
        RECT 124.010 21.020 127.990 21.160 ;
        RECT 127.850 4.000 127.990 21.020 ;
        RECT 127.780 0.000 128.060 4.000 ;
    END
  END mask_rev_in[2]
  PIN mask_rev_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 103.710 143.920 104.040 145.710 ;
        RECT 73.570 132.460 73.980 133.130 ;
        RECT 78.390 131.820 78.560 132.730 ;
      LAYER L1M1_PR_C ;
        RECT 103.830 144.030 104.000 144.200 ;
        RECT 73.590 132.560 73.760 132.730 ;
        RECT 78.390 132.560 78.560 132.730 ;
      LAYER met1 ;
        RECT 103.760 144.180 104.080 144.240 ;
        RECT 103.560 144.040 104.080 144.180 ;
        RECT 103.760 143.980 104.080 144.040 ;
        RECT 72.560 132.710 72.880 132.770 ;
        RECT 73.530 132.710 73.820 132.760 ;
        RECT 78.330 132.710 78.620 132.760 ;
        RECT 72.560 132.570 78.620 132.710 ;
        RECT 72.560 132.510 72.880 132.570 ;
        RECT 73.530 132.530 73.820 132.570 ;
        RECT 78.330 132.530 78.620 132.570 ;
        RECT 78.330 131.970 78.620 132.020 ;
        RECT 78.330 131.830 84.310 131.970 ;
        RECT 78.330 131.790 78.620 131.830 ;
        RECT 84.170 131.230 84.310 131.830 ;
        RECT 103.760 131.230 104.080 131.290 ;
        RECT 84.170 131.090 104.080 131.230 ;
        RECT 103.760 131.030 104.080 131.090 ;
        RECT 20.720 104.590 21.040 104.650 ;
        RECT 72.560 104.590 72.880 104.650 ;
        RECT 20.720 104.450 72.880 104.590 ;
        RECT 20.720 104.390 21.040 104.450 ;
        RECT 72.560 104.390 72.880 104.450 ;
      LAYER via ;
        RECT 103.790 143.980 104.050 144.240 ;
        RECT 72.590 132.510 72.850 132.770 ;
        RECT 103.790 131.030 104.050 131.290 ;
        RECT 20.750 104.390 21.010 104.650 ;
        RECT 72.590 104.390 72.850 104.650 ;
      LAYER met2 ;
        RECT 103.790 143.950 104.050 144.270 ;
        RECT 72.590 132.480 72.850 132.800 ;
        RECT 72.650 104.680 72.790 132.480 ;
        RECT 103.850 131.320 103.990 143.950 ;
        RECT 103.790 131.000 104.050 131.320 ;
        RECT 20.750 104.360 21.010 104.680 ;
        RECT 72.590 104.360 72.850 104.680 ;
        RECT 20.810 101.190 20.950 104.360 ;
        RECT 20.740 100.820 21.020 101.190 ;
      LAYER via2 ;
        RECT 20.740 100.870 21.020 101.150 ;
      LAYER met3 ;
        RECT 0.000 101.160 4.000 101.310 ;
        RECT 20.710 101.160 21.040 101.170 ;
        RECT 0.000 100.860 21.040 101.160 ;
        RECT 0.000 100.710 4.000 100.860 ;
        RECT 20.710 100.840 21.040 100.860 ;
    END
  END mask_rev_in[3]
  PIN mfgr_id[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 45.690 145.630 46.270 146.270 ;
        RECT 45.690 144.220 45.960 145.630 ;
        RECT 45.200 143.950 45.960 144.220 ;
        RECT 45.200 142.950 45.530 143.950 ;
      LAYER L1M1_PR_C ;
        RECT 45.750 145.510 45.920 145.680 ;
      LAYER met1 ;
        RECT 45.200 145.660 45.520 145.720 ;
        RECT 45.690 145.660 45.980 145.710 ;
        RECT 45.200 145.520 45.980 145.660 ;
        RECT 45.200 145.460 45.520 145.520 ;
        RECT 45.690 145.480 45.980 145.520 ;
      LAYER via ;
        RECT 45.230 145.460 45.490 145.720 ;
      LAYER met2 ;
        RECT 45.220 165.200 45.500 169.200 ;
        RECT 45.290 145.750 45.430 165.200 ;
        RECT 45.230 145.430 45.490 145.750 ;
    END
  END mfgr_id[0]
  PIN mfgr_id[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 22.680 22.540 22.930 23.880 ;
        RECT 22.220 22.290 22.930 22.540 ;
        RECT 22.220 21.420 22.470 22.290 ;
        RECT 21.890 20.780 22.470 21.420 ;
      LAYER L1M1_PR_C ;
        RECT 22.230 21.190 22.400 21.360 ;
      LAYER met1 ;
        RECT 22.170 21.340 22.460 21.390 ;
        RECT 23.120 21.340 23.440 21.400 ;
        RECT 22.170 21.200 23.440 21.340 ;
        RECT 22.170 21.160 22.460 21.200 ;
        RECT 23.120 21.140 23.440 21.200 ;
      LAYER via ;
        RECT 23.150 21.140 23.410 21.400 ;
      LAYER met2 ;
        RECT 23.150 21.110 23.410 21.430 ;
        RECT 23.210 4.000 23.350 21.110 ;
        RECT 23.140 0.000 23.420 4.000 ;
    END
  END mfgr_id[10]
  PIN mfgr_id[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 137.360 59.550 137.690 60.550 ;
        RECT 137.360 59.280 138.120 59.550 ;
        RECT 137.850 57.870 138.120 59.280 ;
        RECT 137.850 57.230 138.430 57.870 ;
      LAYER L1M1_PR_C ;
        RECT 137.910 59.300 138.080 59.470 ;
      LAYER met1 ;
        RECT 137.840 59.450 138.160 59.510 ;
        RECT 137.640 59.310 138.160 59.450 ;
        RECT 137.840 59.250 138.160 59.310 ;
      LAYER via ;
        RECT 137.870 59.250 138.130 59.510 ;
      LAYER met2 ;
        RECT 137.860 59.380 138.140 59.750 ;
        RECT 137.870 59.220 138.130 59.380 ;
      LAYER via2 ;
        RECT 137.860 59.430 138.140 59.710 ;
      LAYER met3 ;
        RECT 137.830 59.720 138.160 59.730 ;
        RECT 144.160 59.720 148.160 59.870 ;
        RECT 137.830 59.420 148.160 59.720 ;
        RECT 137.830 59.400 138.160 59.420 ;
        RECT 144.160 59.270 148.160 59.420 ;
    END
  END mfgr_id[11]
  PIN mfgr_id[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 65.090 149.520 65.670 150.160 ;
        RECT 65.420 148.650 65.670 149.520 ;
        RECT 65.420 148.400 66.130 148.650 ;
        RECT 65.880 147.060 66.130 148.400 ;
      LAYER L1M1_PR_C ;
        RECT 65.430 149.580 65.600 149.750 ;
      LAYER met1 ;
        RECT 65.370 149.730 65.660 149.780 ;
        RECT 66.320 149.730 66.640 149.790 ;
        RECT 65.370 149.590 66.640 149.730 ;
        RECT 65.370 149.550 65.660 149.590 ;
        RECT 66.320 149.530 66.640 149.590 ;
      LAYER via ;
        RECT 66.350 149.530 66.610 149.790 ;
      LAYER met2 ;
        RECT 66.340 165.200 66.620 169.200 ;
        RECT 66.410 149.820 66.550 165.200 ;
        RECT 66.350 149.500 66.610 149.820 ;
    END
  END mfgr_id[1]
  PIN mfgr_id[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 135.480 87.660 135.730 89.000 ;
        RECT 135.020 87.410 135.730 87.660 ;
        RECT 135.020 86.540 135.270 87.410 ;
        RECT 134.690 85.900 135.270 86.540 ;
      LAYER L1M1_PR_C ;
        RECT 135.510 88.530 135.680 88.700 ;
      LAYER met1 ;
        RECT 135.440 88.680 135.760 88.740 ;
        RECT 135.240 88.540 135.760 88.680 ;
        RECT 135.440 88.480 135.760 88.540 ;
      LAYER via ;
        RECT 135.470 88.480 135.730 88.740 ;
      LAYER met2 ;
        RECT 135.460 90.460 135.740 90.830 ;
        RECT 135.530 88.770 135.670 90.460 ;
        RECT 135.470 88.450 135.730 88.770 ;
      LAYER via2 ;
        RECT 135.460 90.510 135.740 90.790 ;
      LAYER met3 ;
        RECT 135.430 90.800 135.760 90.810 ;
        RECT 144.160 90.800 148.160 90.950 ;
        RECT 135.430 90.500 148.160 90.800 ;
        RECT 135.430 90.480 135.760 90.500 ;
        RECT 144.160 90.350 148.160 90.500 ;
    END
  END mfgr_id[2]
  PIN mfgr_id[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 128.730 145.630 129.310 146.270 ;
        RECT 128.730 144.220 129.000 145.630 ;
        RECT 128.240 143.950 129.000 144.220 ;
        RECT 128.240 142.950 128.570 143.950 ;
      LAYER L1M1_PR_C ;
        RECT 128.790 145.510 128.960 145.680 ;
      LAYER met1 ;
        RECT 128.720 145.660 129.040 145.720 ;
        RECT 128.520 145.520 129.040 145.660 ;
        RECT 128.720 145.460 129.040 145.520 ;
      LAYER via ;
        RECT 128.750 145.460 129.010 145.720 ;
      LAYER met2 ;
        RECT 128.740 165.200 129.020 169.200 ;
        RECT 128.810 145.750 128.950 165.200 ;
        RECT 128.750 145.430 129.010 145.750 ;
    END
  END mfgr_id[3]
  PIN mfgr_id[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 138.840 38.820 139.090 40.160 ;
        RECT 138.380 38.570 139.090 38.820 ;
        RECT 138.380 37.700 138.630 38.570 ;
        RECT 138.050 37.060 138.630 37.700 ;
      LAYER L1M1_PR_C ;
        RECT 138.870 39.690 139.040 39.860 ;
      LAYER met1 ;
        RECT 138.800 39.840 139.120 39.900 ;
        RECT 138.600 39.700 139.120 39.840 ;
        RECT 138.800 39.640 139.120 39.700 ;
      LAYER via ;
        RECT 138.830 39.640 139.090 39.900 ;
      LAYER met2 ;
        RECT 138.820 43.100 139.100 43.470 ;
        RECT 138.890 39.930 139.030 43.100 ;
        RECT 138.830 39.610 139.090 39.930 ;
      LAYER via2 ;
        RECT 138.820 43.150 139.100 43.430 ;
      LAYER met3 ;
        RECT 138.790 43.440 139.120 43.450 ;
        RECT 144.160 43.440 148.160 43.590 ;
        RECT 138.790 43.140 148.160 43.440 ;
        RECT 138.790 43.120 139.120 43.140 ;
        RECT 144.160 42.990 148.160 43.140 ;
    END
  END mfgr_id[4]
  PIN mfgr_id[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 11.600 132.810 11.930 133.810 ;
        RECT 11.600 132.540 12.360 132.810 ;
        RECT 12.090 131.130 12.360 132.540 ;
        RECT 12.090 130.490 12.670 131.130 ;
      LAYER L1M1_PR_C ;
        RECT 11.670 133.300 11.840 133.470 ;
      LAYER met1 ;
        RECT 11.600 133.450 11.920 133.510 ;
        RECT 11.400 133.310 11.920 133.450 ;
        RECT 11.600 133.250 11.920 133.310 ;
      LAYER via ;
        RECT 11.630 133.250 11.890 133.510 ;
      LAYER met2 ;
        RECT 11.620 133.380 11.900 133.750 ;
        RECT 11.630 133.220 11.890 133.380 ;
      LAYER via2 ;
        RECT 11.620 133.430 11.900 133.710 ;
      LAYER met3 ;
        RECT 0.000 133.720 4.000 133.870 ;
        RECT 11.590 133.720 11.920 133.730 ;
        RECT 0.000 133.420 11.920 133.720 ;
        RECT 0.000 133.270 4.000 133.420 ;
        RECT 11.590 133.400 11.920 133.420 ;
    END
  END mfgr_id[5]
  PIN mfgr_id[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 75.170 149.520 75.750 150.160 ;
        RECT 75.500 148.650 75.750 149.520 ;
        RECT 75.500 148.400 76.210 148.650 ;
        RECT 75.960 147.060 76.210 148.400 ;
      LAYER L1M1_PR_C ;
        RECT 75.510 149.580 75.680 149.750 ;
      LAYER met1 ;
        RECT 75.450 149.730 75.740 149.780 ;
        RECT 76.880 149.730 77.200 149.790 ;
        RECT 75.450 149.590 77.200 149.730 ;
        RECT 75.450 149.550 75.740 149.590 ;
        RECT 76.880 149.530 77.200 149.590 ;
      LAYER via ;
        RECT 76.910 149.530 77.170 149.790 ;
      LAYER met2 ;
        RECT 76.900 165.200 77.180 169.200 ;
        RECT 76.970 149.820 77.110 165.200 ;
        RECT 76.910 149.500 77.170 149.820 ;
    END
  END mfgr_id[6]
  PIN mfgr_id[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 135.440 26.990 135.770 27.990 ;
        RECT 135.440 26.720 136.200 26.990 ;
        RECT 135.930 25.310 136.200 26.720 ;
        RECT 135.930 24.670 136.510 25.310 ;
      LAYER L1M1_PR_C ;
        RECT 135.990 26.740 136.160 26.910 ;
      LAYER met1 ;
        RECT 135.920 26.890 136.240 26.950 ;
        RECT 135.720 26.750 136.240 26.890 ;
        RECT 135.920 26.690 136.240 26.750 ;
      LAYER via ;
        RECT 135.950 26.690 136.210 26.950 ;
      LAYER met2 ;
        RECT 135.940 26.820 136.220 27.190 ;
        RECT 135.950 26.660 136.210 26.820 ;
      LAYER via2 ;
        RECT 135.940 26.870 136.220 27.150 ;
      LAYER met3 ;
        RECT 135.910 27.160 136.240 27.170 ;
        RECT 144.160 27.160 148.160 27.310 ;
        RECT 135.910 26.860 148.160 27.160 ;
        RECT 135.910 26.840 136.240 26.860 ;
        RECT 144.160 26.710 148.160 26.860 ;
    END
  END mfgr_id[7]
  PIN mfgr_id[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 23.120 149.090 23.450 150.090 ;
        RECT 23.120 148.820 23.880 149.090 ;
        RECT 23.610 147.410 23.880 148.820 ;
        RECT 23.610 146.770 24.190 147.410 ;
      LAYER L1M1_PR_C ;
        RECT 23.190 149.580 23.360 149.750 ;
      LAYER met1 ;
        RECT 23.130 149.730 23.420 149.780 ;
        RECT 24.080 149.730 24.400 149.790 ;
        RECT 23.130 149.590 24.400 149.730 ;
        RECT 23.130 149.550 23.420 149.590 ;
        RECT 24.080 149.530 24.400 149.590 ;
      LAYER via ;
        RECT 24.110 149.530 24.370 149.790 ;
      LAYER met2 ;
        RECT 24.100 165.200 24.380 169.200 ;
        RECT 24.170 149.820 24.310 165.200 ;
        RECT 24.110 149.500 24.370 149.820 ;
    END
  END mfgr_id[8]
  PIN mfgr_id[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 16.880 18.850 17.210 19.850 ;
        RECT 16.880 18.580 17.640 18.850 ;
        RECT 17.370 17.170 17.640 18.580 ;
        RECT 17.370 16.530 17.950 17.170 ;
      LAYER L1M1_PR_C ;
        RECT 17.430 18.600 17.600 18.770 ;
      LAYER met1 ;
        RECT 17.370 18.750 17.660 18.800 ;
        RECT 37.040 18.750 37.360 18.810 ;
        RECT 54.800 18.750 55.120 18.810 ;
        RECT 17.370 18.610 37.360 18.750 ;
        RECT 17.370 18.570 17.660 18.610 ;
        RECT 37.040 18.550 37.360 18.610 ;
        RECT 38.570 18.610 55.120 18.750 ;
        RECT 38.570 18.440 38.710 18.610 ;
        RECT 54.800 18.550 55.120 18.610 ;
        RECT 38.480 18.180 38.800 18.440 ;
      LAYER via ;
        RECT 37.070 18.550 37.330 18.810 ;
        RECT 54.830 18.550 55.090 18.810 ;
        RECT 38.510 18.180 38.770 18.440 ;
      LAYER met2 ;
        RECT 37.070 18.520 37.330 18.840 ;
        RECT 54.830 18.520 55.090 18.840 ;
        RECT 37.130 18.010 37.270 18.520 ;
        RECT 38.510 18.150 38.770 18.470 ;
        RECT 38.570 18.010 38.710 18.150 ;
        RECT 37.130 17.870 38.710 18.010 ;
        RECT 54.890 4.000 55.030 18.520 ;
        RECT 54.820 0.000 55.100 4.000 ;
    END
  END mfgr_id[9]
  PIN pll_bias_ena
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 11.640 144.640 11.890 145.980 ;
        RECT 11.180 144.390 11.890 144.640 ;
        RECT 11.180 143.520 11.430 144.390 ;
        RECT 10.850 142.880 11.430 143.520 ;
      LAYER L1M1_PR_C ;
        RECT 11.190 143.660 11.360 143.830 ;
      LAYER met1 ;
        RECT 2.960 143.810 3.280 143.870 ;
        RECT 11.130 143.810 11.420 143.860 ;
        RECT 2.960 143.670 11.420 143.810 ;
        RECT 2.960 143.610 3.280 143.670 ;
        RECT 11.130 143.630 11.420 143.670 ;
      LAYER via ;
        RECT 2.990 143.610 3.250 143.870 ;
      LAYER met2 ;
        RECT 2.980 165.200 3.260 169.200 ;
        RECT 3.050 143.900 3.190 165.200 ;
        RECT 2.990 143.580 3.250 143.900 ;
    END
  END pll_bias_ena
  PIN pll_bypass
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 96.130 75.490 96.860 75.820 ;
        RECT 104.370 75.370 104.970 75.760 ;
        RECT 128.660 73.590 129.000 76.660 ;
      LAYER L1M1_PR_C ;
        RECT 96.150 75.580 96.320 75.750 ;
        RECT 104.790 75.580 104.960 75.750 ;
        RECT 128.790 74.100 128.960 74.270 ;
      LAYER met1 ;
        RECT 96.090 75.550 96.380 75.780 ;
        RECT 104.720 75.730 105.040 75.790 ;
        RECT 97.610 75.590 105.040 75.730 ;
        RECT 96.170 75.360 96.310 75.550 ;
        RECT 97.610 75.360 97.750 75.590 ;
        RECT 104.720 75.530 105.040 75.590 ;
        RECT 96.170 75.220 97.750 75.360 ;
        RECT 104.720 74.250 105.040 74.310 ;
        RECT 128.720 74.250 129.040 74.310 ;
        RECT 104.720 74.110 129.040 74.250 ;
        RECT 104.720 74.050 105.040 74.110 ;
        RECT 128.720 74.050 129.040 74.110 ;
      LAYER via ;
        RECT 104.750 75.530 105.010 75.790 ;
        RECT 104.750 74.050 105.010 74.310 ;
        RECT 128.750 74.050 129.010 74.310 ;
      LAYER met2 ;
        RECT 104.750 75.500 105.010 75.820 ;
        RECT 104.810 74.340 104.950 75.500 ;
        RECT 104.750 74.020 105.010 74.340 ;
        RECT 128.750 74.020 129.010 74.340 ;
        RECT 128.810 39.660 128.950 74.020 ;
        RECT 128.330 39.520 128.950 39.660 ;
        RECT 128.330 10.910 128.470 39.520 ;
        RECT 128.260 10.540 128.540 10.910 ;
      LAYER via2 ;
        RECT 128.260 10.590 128.540 10.870 ;
      LAYER met3 ;
        RECT 128.230 10.880 128.560 10.890 ;
        RECT 144.160 10.880 148.160 11.030 ;
        RECT 128.230 10.580 148.160 10.880 ;
        RECT 128.230 10.560 128.560 10.580 ;
        RECT 144.160 10.430 148.160 10.580 ;
    END
  END pll_bypass
  PIN pll_cp_ena
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 64.820 118.680 65.170 121.650 ;
        RECT 67.810 119.580 68.520 119.970 ;
      LAYER L1M1_PR_C ;
        RECT 64.950 119.610 65.120 119.780 ;
        RECT 68.310 119.610 68.480 119.780 ;
      LAYER met1 ;
        RECT 94.160 120.500 94.480 120.560 ;
        RECT 90.890 120.360 94.480 120.500 ;
        RECT 81.290 119.990 88.630 120.130 ;
        RECT 64.890 119.760 65.180 119.810 ;
        RECT 68.250 119.760 68.540 119.810 ;
        RECT 64.890 119.620 76.630 119.760 ;
        RECT 64.890 119.580 65.180 119.620 ;
        RECT 68.250 119.580 68.540 119.620 ;
        RECT 76.490 119.020 76.630 119.620 ;
        RECT 81.290 119.020 81.430 119.990 ;
        RECT 88.490 119.760 88.630 119.990 ;
        RECT 90.890 119.760 91.030 120.360 ;
        RECT 94.160 120.300 94.480 120.360 ;
        RECT 88.490 119.620 91.030 119.760 ;
        RECT 76.490 118.880 81.430 119.020 ;
      LAYER via ;
        RECT 94.190 120.300 94.450 120.560 ;
      LAYER met2 ;
        RECT 97.060 165.200 97.340 169.200 ;
        RECT 97.130 151.400 97.270 165.200 ;
        RECT 94.730 151.260 97.270 151.400 ;
        RECT 94.730 121.060 94.870 151.260 ;
        RECT 94.250 120.920 94.870 121.060 ;
        RECT 94.250 120.590 94.390 120.920 ;
        RECT 94.190 120.270 94.450 120.590 ;
    END
  END pll_cp_ena
  PIN pll_trim[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 77.410 111.400 78.140 111.730 ;
        RECT 43.700 106.150 44.040 109.220 ;
        RECT 34.690 103.260 35.850 103.500 ;
      LAYER L1M1_PR_C ;
        RECT 77.430 111.470 77.600 111.640 ;
        RECT 43.830 106.660 44.000 106.830 ;
        RECT 34.710 103.330 34.880 103.500 ;
      LAYER met1 ;
        RECT 77.370 111.440 77.660 111.670 ;
        RECT 72.080 111.250 72.400 111.310 ;
        RECT 77.450 111.250 77.590 111.440 ;
        RECT 72.080 111.110 77.590 111.250 ;
        RECT 72.080 111.050 72.400 111.110 ;
        RECT 72.080 107.550 72.400 107.610 ;
        RECT 43.850 107.410 72.400 107.550 ;
        RECT 33.200 106.810 33.520 106.870 ;
        RECT 43.850 106.860 43.990 107.410 ;
        RECT 72.080 107.350 72.400 107.410 ;
        RECT 43.770 106.810 44.060 106.860 ;
        RECT 33.200 106.670 44.060 106.810 ;
        RECT 33.200 106.610 33.520 106.670 ;
        RECT 43.770 106.630 44.060 106.670 ;
        RECT 34.650 103.300 34.940 103.530 ;
        RECT 33.200 103.110 33.520 103.170 ;
        RECT 34.730 103.110 34.870 103.300 ;
        RECT 33.200 102.970 34.870 103.110 ;
        RECT 33.200 102.910 33.520 102.970 ;
        RECT 21.200 56.120 21.520 56.180 ;
        RECT 31.280 56.120 31.600 56.180 ;
        RECT 21.200 55.980 31.600 56.120 ;
        RECT 21.200 55.920 21.520 55.980 ;
        RECT 31.280 55.920 31.600 55.980 ;
      LAYER via ;
        RECT 72.110 111.050 72.370 111.310 ;
        RECT 33.230 106.610 33.490 106.870 ;
        RECT 72.110 107.350 72.370 107.610 ;
        RECT 33.230 102.910 33.490 103.170 ;
        RECT 21.230 55.920 21.490 56.180 ;
        RECT 31.310 55.920 31.570 56.180 ;
      LAYER met2 ;
        RECT 72.110 111.020 72.370 111.340 ;
        RECT 72.170 107.640 72.310 111.020 ;
        RECT 72.110 107.320 72.370 107.640 ;
        RECT 33.230 106.580 33.490 106.900 ;
        RECT 33.290 103.200 33.430 106.580 ;
        RECT 33.230 102.880 33.490 103.200 ;
        RECT 33.290 67.150 33.430 102.880 ;
        RECT 31.300 66.780 31.580 67.150 ;
        RECT 33.220 66.780 33.500 67.150 ;
        RECT 31.370 56.210 31.510 66.780 ;
        RECT 21.230 55.890 21.490 56.210 ;
        RECT 31.310 55.890 31.570 56.210 ;
        RECT 21.290 52.350 21.430 55.890 ;
        RECT 21.220 51.980 21.500 52.350 ;
      LAYER via2 ;
        RECT 31.300 66.830 31.580 67.110 ;
        RECT 33.220 66.830 33.500 67.110 ;
        RECT 21.220 52.030 21.500 52.310 ;
      LAYER met3 ;
        RECT 31.270 67.120 31.600 67.130 ;
        RECT 33.190 67.120 33.520 67.130 ;
        RECT 31.270 66.820 33.520 67.120 ;
        RECT 31.270 66.800 31.600 66.820 ;
        RECT 33.190 66.800 33.520 66.820 ;
        RECT 0.000 52.320 4.000 52.470 ;
        RECT 21.190 52.320 21.520 52.330 ;
        RECT 0.000 52.020 21.520 52.320 ;
        RECT 0.000 51.870 4.000 52.020 ;
        RECT 21.190 52.000 21.520 52.020 ;
    END
  END pll_trim[0]
  PIN pll_trim[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 64.340 106.150 64.680 109.220 ;
        RECT 61.570 103.300 62.280 103.690 ;
      LAYER L1M1_PR_C ;
        RECT 64.470 106.660 64.640 106.830 ;
        RECT 61.590 103.330 61.760 103.500 ;
      LAYER met1 ;
        RECT 61.040 106.810 61.360 106.870 ;
        RECT 64.410 106.810 64.700 106.860 ;
        RECT 61.040 106.670 64.700 106.810 ;
        RECT 61.040 106.610 61.360 106.670 ;
        RECT 64.410 106.630 64.700 106.670 ;
        RECT 61.040 103.480 61.360 103.540 ;
        RECT 61.530 103.480 61.820 103.530 ;
        RECT 61.040 103.340 61.820 103.480 ;
        RECT 61.040 103.280 61.360 103.340 ;
        RECT 61.530 103.300 61.820 103.340 ;
        RECT 62.960 50.570 63.280 50.630 ;
        RECT 63.440 50.570 63.760 50.630 ;
        RECT 62.960 50.430 63.760 50.570 ;
        RECT 62.960 50.370 63.280 50.430 ;
        RECT 63.440 50.370 63.760 50.430 ;
        RECT 62.960 25.410 63.280 25.470 ;
        RECT 75.920 25.410 76.240 25.470 ;
        RECT 62.960 25.270 76.240 25.410 ;
        RECT 62.960 25.210 63.280 25.270 ;
        RECT 75.920 25.210 76.240 25.270 ;
      LAYER via ;
        RECT 61.070 106.610 61.330 106.870 ;
        RECT 61.070 103.280 61.330 103.540 ;
        RECT 62.990 50.370 63.250 50.630 ;
        RECT 63.470 50.370 63.730 50.630 ;
        RECT 62.990 25.210 63.250 25.470 ;
        RECT 75.950 25.210 76.210 25.470 ;
      LAYER met2 ;
        RECT 61.070 106.580 61.330 106.900 ;
        RECT 61.130 103.570 61.270 106.580 ;
        RECT 61.070 103.250 61.330 103.570 ;
        RECT 61.130 101.190 61.270 103.250 ;
        RECT 61.060 100.820 61.340 101.190 ;
        RECT 63.460 100.820 63.740 101.190 ;
        RECT 63.530 50.660 63.670 100.820 ;
        RECT 62.990 50.340 63.250 50.660 ;
        RECT 63.470 50.340 63.730 50.660 ;
        RECT 63.050 25.500 63.190 50.340 ;
        RECT 62.990 25.180 63.250 25.500 ;
        RECT 75.950 25.180 76.210 25.500 ;
        RECT 76.010 4.000 76.150 25.180 ;
        RECT 75.940 0.000 76.220 4.000 ;
      LAYER via2 ;
        RECT 61.060 100.870 61.340 101.150 ;
        RECT 63.460 100.870 63.740 101.150 ;
      LAYER met3 ;
        RECT 61.030 101.160 61.360 101.170 ;
        RECT 63.430 101.160 63.760 101.170 ;
        RECT 61.030 100.860 63.760 101.160 ;
        RECT 61.030 100.840 61.360 100.860 ;
        RECT 63.430 100.840 63.760 100.860 ;
    END
  END pll_trim[1]
  PIN pll_trim[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 45.140 138.710 45.480 141.780 ;
        RECT 38.050 127.680 39.210 127.920 ;
        RECT 92.570 111.400 93.480 111.730 ;
      LAYER L1M1_PR_C ;
        RECT 45.270 141.070 45.440 141.240 ;
        RECT 39.030 127.750 39.200 127.920 ;
        RECT 92.790 111.470 92.960 111.640 ;
      LAYER met1 ;
        RECT 92.720 143.810 93.040 143.870 ;
        RECT 129.200 143.810 129.520 143.870 ;
        RECT 92.720 143.670 129.520 143.810 ;
        RECT 92.720 143.610 93.040 143.670 ;
        RECT 129.200 143.610 129.520 143.670 ;
        RECT 43.280 141.220 43.600 141.280 ;
        RECT 45.210 141.220 45.500 141.270 ;
        RECT 92.720 141.220 93.040 141.280 ;
        RECT 43.280 141.080 93.040 141.220 ;
        RECT 43.280 141.020 43.600 141.080 ;
        RECT 45.210 141.040 45.500 141.080 ;
        RECT 92.720 141.020 93.040 141.080 ;
        RECT 43.280 128.270 43.600 128.330 ;
        RECT 39.050 128.130 43.600 128.270 ;
        RECT 39.050 127.950 39.190 128.130 ;
        RECT 43.280 128.070 43.600 128.130 ;
        RECT 38.970 127.720 39.260 127.950 ;
        RECT 92.720 111.620 93.040 111.680 ;
        RECT 92.520 111.480 93.040 111.620 ;
        RECT 92.720 111.420 93.040 111.480 ;
      LAYER via ;
        RECT 92.750 143.610 93.010 143.870 ;
        RECT 129.230 143.610 129.490 143.870 ;
        RECT 43.310 141.020 43.570 141.280 ;
        RECT 92.750 141.020 93.010 141.280 ;
        RECT 43.310 128.070 43.570 128.330 ;
        RECT 92.750 111.420 93.010 111.680 ;
      LAYER met2 ;
        RECT 129.220 155.580 129.500 155.950 ;
        RECT 129.290 143.900 129.430 155.580 ;
        RECT 92.750 143.580 93.010 143.900 ;
        RECT 129.230 143.580 129.490 143.900 ;
        RECT 92.810 141.310 92.950 143.580 ;
        RECT 43.310 140.990 43.570 141.310 ;
        RECT 92.750 140.990 93.010 141.310 ;
        RECT 43.370 128.360 43.510 140.990 ;
        RECT 43.310 128.040 43.570 128.360 ;
        RECT 92.810 111.710 92.950 140.990 ;
        RECT 92.750 111.390 93.010 111.710 ;
      LAYER via2 ;
        RECT 129.220 155.630 129.500 155.910 ;
      LAYER met3 ;
        RECT 129.190 155.920 129.520 155.930 ;
        RECT 144.160 155.920 148.160 156.070 ;
        RECT 129.190 155.620 148.160 155.920 ;
        RECT 129.190 155.600 129.520 155.620 ;
        RECT 144.160 155.470 148.160 155.620 ;
    END
  END pll_trim[2]
  PIN pll_trim[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 62.420 138.710 62.760 141.780 ;
        RECT 48.990 124.420 49.320 124.660 ;
        RECT 87.900 119.560 88.200 119.890 ;
      LAYER L1M1_PR_C ;
        RECT 62.550 139.590 62.720 139.760 ;
        RECT 49.110 124.420 49.280 124.590 ;
        RECT 87.990 119.610 88.160 119.780 ;
      LAYER met1 ;
        RECT 87.440 140.110 87.760 140.170 ;
        RECT 62.570 139.970 87.760 140.110 ;
        RECT 62.570 139.800 62.710 139.970 ;
        RECT 87.440 139.910 87.760 139.970 ;
        RECT 62.480 139.740 62.800 139.800 ;
        RECT 62.280 139.600 62.800 139.740 ;
        RECT 62.480 139.540 62.800 139.600 ;
        RECT 49.050 124.570 49.340 124.620 ;
        RECT 62.480 124.570 62.800 124.630 ;
        RECT 49.050 124.430 62.800 124.570 ;
        RECT 49.050 124.390 49.340 124.430 ;
        RECT 62.480 124.370 62.800 124.430 ;
        RECT 87.440 119.760 87.760 119.820 ;
        RECT 87.930 119.760 88.220 119.810 ;
        RECT 87.440 119.620 88.220 119.760 ;
        RECT 87.440 119.560 87.760 119.620 ;
        RECT 87.930 119.580 88.220 119.620 ;
      LAYER via ;
        RECT 87.470 139.910 87.730 140.170 ;
        RECT 62.510 139.540 62.770 139.800 ;
        RECT 62.510 124.370 62.770 124.630 ;
        RECT 87.470 119.560 87.730 119.820 ;
      LAYER met2 ;
        RECT 87.460 165.200 87.740 169.200 ;
        RECT 87.530 140.200 87.670 165.200 ;
        RECT 87.470 139.880 87.730 140.200 ;
        RECT 62.510 139.510 62.770 139.830 ;
        RECT 62.570 124.660 62.710 139.510 ;
        RECT 62.510 124.340 62.770 124.660 ;
        RECT 87.530 119.850 87.670 139.880 ;
        RECT 87.470 119.530 87.730 119.850 ;
    END
  END pll_trim[3]
  PIN pll_vco_ena
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 64.340 126.820 64.690 129.790 ;
        RECT 67.350 127.750 67.520 129.400 ;
        RECT 67.810 127.720 68.520 128.110 ;
      LAYER L1M1_PR_C ;
        RECT 64.470 127.750 64.640 127.920 ;
        RECT 67.350 129.230 67.520 129.400 ;
        RECT 67.830 127.750 68.000 127.920 ;
      LAYER met1 ;
        RECT 67.290 129.380 67.580 129.430 ;
        RECT 67.290 129.240 78.550 129.380 ;
        RECT 67.290 129.200 67.580 129.240 ;
        RECT 78.410 129.010 78.550 129.240 ;
        RECT 78.410 128.870 101.590 129.010 ;
        RECT 101.450 128.640 101.590 128.870 ;
        RECT 117.680 128.640 118.000 128.700 ;
        RECT 101.450 128.500 118.000 128.640 ;
        RECT 117.680 128.440 118.000 128.500 ;
        RECT 64.410 127.900 64.700 127.950 ;
        RECT 67.290 127.900 67.580 127.950 ;
        RECT 67.770 127.900 68.060 127.950 ;
        RECT 64.410 127.760 68.060 127.900 ;
        RECT 64.410 127.720 64.700 127.760 ;
        RECT 67.290 127.720 67.580 127.760 ;
        RECT 67.770 127.720 68.060 127.760 ;
      LAYER via ;
        RECT 117.710 128.440 117.970 128.700 ;
      LAYER met2 ;
        RECT 118.180 165.200 118.460 169.200 ;
        RECT 118.250 135.860 118.390 165.200 ;
        RECT 117.770 135.720 118.390 135.860 ;
        RECT 117.770 128.730 117.910 135.720 ;
        RECT 117.710 128.410 117.970 128.730 ;
    END
  END pll_vco_ena
  PIN prod_id[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 135.440 75.830 135.770 76.830 ;
        RECT 135.440 75.560 136.200 75.830 ;
        RECT 135.930 74.150 136.200 75.560 ;
        RECT 135.930 73.510 136.510 74.150 ;
      LAYER L1M1_PR_C ;
        RECT 135.990 75.580 136.160 75.750 ;
      LAYER met1 ;
        RECT 135.920 75.730 136.240 75.790 ;
        RECT 135.720 75.590 136.240 75.730 ;
        RECT 135.920 75.530 136.240 75.590 ;
      LAYER via ;
        RECT 135.950 75.530 136.210 75.790 ;
      LAYER met2 ;
        RECT 135.940 75.660 136.220 76.030 ;
        RECT 135.950 75.500 136.210 75.660 ;
      LAYER via2 ;
        RECT 135.940 75.710 136.220 75.990 ;
      LAYER met3 ;
        RECT 135.910 76.000 136.240 76.010 ;
        RECT 144.160 76.000 148.160 76.150 ;
        RECT 135.910 75.700 148.160 76.000 ;
        RECT 135.910 75.680 136.240 75.700 ;
        RECT 144.160 75.550 148.160 75.700 ;
    END
  END prod_id[0]
  PIN prod_id[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 20.450 19.280 21.030 19.920 ;
        RECT 20.780 18.410 21.030 19.280 ;
        RECT 20.780 18.160 21.490 18.410 ;
        RECT 21.240 16.820 21.490 18.160 ;
      LAYER L1M1_PR_C ;
        RECT 21.270 17.860 21.440 18.030 ;
      LAYER met1 ;
        RECT 21.210 18.010 21.500 18.060 ;
        RECT 44.240 18.010 44.560 18.070 ;
        RECT 21.210 17.870 37.750 18.010 ;
        RECT 21.210 17.830 21.500 17.870 ;
        RECT 37.610 17.270 37.750 17.870 ;
        RECT 38.570 17.870 44.560 18.010 ;
        RECT 38.570 17.270 38.710 17.870 ;
        RECT 44.240 17.810 44.560 17.870 ;
        RECT 37.610 17.130 38.710 17.270 ;
      LAYER via ;
        RECT 44.270 17.810 44.530 18.070 ;
      LAYER met2 ;
        RECT 44.270 17.780 44.530 18.100 ;
        RECT 44.330 4.000 44.470 17.780 ;
        RECT 44.260 0.000 44.540 4.000 ;
    END
  END prod_id[1]
  PIN prod_id[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 18.810 23.530 19.390 24.170 ;
        RECT 18.810 22.120 19.080 23.530 ;
        RECT 18.320 21.850 19.080 22.120 ;
        RECT 18.320 20.850 18.650 21.850 ;
      LAYER L1M1_PR_C ;
        RECT 18.870 22.670 19.040 22.840 ;
      LAYER met1 ;
        RECT 18.810 22.820 19.100 22.870 ;
        RECT 33.680 22.820 34.000 22.880 ;
        RECT 18.810 22.680 34.000 22.820 ;
        RECT 18.810 22.640 19.100 22.680 ;
        RECT 33.680 22.620 34.000 22.680 ;
      LAYER via ;
        RECT 33.710 22.620 33.970 22.880 ;
      LAYER met2 ;
        RECT 33.710 22.590 33.970 22.910 ;
        RECT 33.770 4.000 33.910 22.590 ;
        RECT 33.700 0.000 33.980 4.000 ;
    END
  END prod_id[2]
  PIN prod_id[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 135.440 18.850 135.770 19.850 ;
        RECT 135.440 18.580 136.200 18.850 ;
        RECT 135.930 17.170 136.200 18.580 ;
        RECT 135.930 16.530 136.510 17.170 ;
      LAYER L1M1_PR_C ;
        RECT 135.990 17.120 136.160 17.290 ;
      LAYER met1 ;
        RECT 135.930 17.270 136.220 17.320 ;
        RECT 138.320 17.270 138.640 17.330 ;
        RECT 135.930 17.130 138.640 17.270 ;
        RECT 135.930 17.090 136.220 17.130 ;
        RECT 138.320 17.070 138.640 17.130 ;
      LAYER via ;
        RECT 138.350 17.070 138.610 17.330 ;
      LAYER met2 ;
        RECT 138.350 17.040 138.610 17.360 ;
        RECT 138.410 4.000 138.550 17.040 ;
        RECT 138.340 0.000 138.620 4.000 ;
    END
  END prod_id[3]
  PIN prod_id[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 121.040 18.850 121.370 19.850 ;
        RECT 121.040 18.580 121.800 18.850 ;
        RECT 121.530 17.170 121.800 18.580 ;
        RECT 121.530 16.530 122.110 17.170 ;
      LAYER L1M1_PR_C ;
        RECT 121.590 17.490 121.760 17.660 ;
      LAYER met1 ;
        RECT 106.640 17.640 106.960 17.700 ;
        RECT 121.530 17.640 121.820 17.690 ;
        RECT 106.640 17.500 121.820 17.640 ;
        RECT 106.640 17.440 106.960 17.500 ;
        RECT 121.530 17.460 121.820 17.500 ;
      LAYER via ;
        RECT 106.670 17.440 106.930 17.700 ;
      LAYER met2 ;
        RECT 106.670 17.410 106.930 17.730 ;
        RECT 106.730 4.000 106.870 17.410 ;
        RECT 106.660 0.000 106.940 4.000 ;
    END
  END prod_id[4]
  PIN prod_id[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 125.360 18.850 125.690 19.850 ;
        RECT 125.360 18.580 126.120 18.850 ;
        RECT 125.850 17.170 126.120 18.580 ;
        RECT 125.850 16.530 126.430 17.170 ;
      LAYER L1M1_PR_C ;
        RECT 125.910 17.860 126.080 18.030 ;
      LAYER met1 ;
        RECT 86.480 18.010 86.800 18.070 ;
        RECT 125.850 18.010 126.140 18.060 ;
        RECT 86.480 17.870 126.140 18.010 ;
        RECT 86.480 17.810 86.800 17.870 ;
        RECT 125.850 17.830 126.140 17.870 ;
      LAYER via ;
        RECT 86.510 17.810 86.770 18.070 ;
      LAYER met2 ;
        RECT 86.510 17.780 86.770 18.100 ;
        RECT 86.570 4.000 86.710 17.780 ;
        RECT 86.500 0.000 86.780 4.000 ;
    END
  END prod_id[5]
  PIN prod_id[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 12.560 18.850 12.890 19.850 ;
        RECT 12.560 18.580 13.320 18.850 ;
        RECT 13.050 17.170 13.320 18.580 ;
        RECT 13.050 16.530 13.630 17.170 ;
      LAYER L1M1_PR_C ;
        RECT 13.110 17.120 13.280 17.290 ;
      LAYER met1 ;
        RECT 13.040 17.270 13.360 17.330 ;
        RECT 12.840 17.130 13.360 17.270 ;
        RECT 13.040 17.070 13.360 17.130 ;
        RECT 13.040 15.050 13.360 15.110 ;
        RECT 65.360 15.050 65.680 15.110 ;
        RECT 13.040 14.910 65.680 15.050 ;
        RECT 13.040 14.850 13.360 14.910 ;
        RECT 65.360 14.850 65.680 14.910 ;
      LAYER via ;
        RECT 13.070 17.070 13.330 17.330 ;
        RECT 13.070 14.850 13.330 15.110 ;
        RECT 65.390 14.850 65.650 15.110 ;
      LAYER met2 ;
        RECT 13.070 17.040 13.330 17.360 ;
        RECT 13.130 15.140 13.270 17.040 ;
        RECT 13.070 14.820 13.330 15.140 ;
        RECT 65.390 14.820 65.650 15.140 ;
        RECT 65.450 4.000 65.590 14.820 ;
        RECT 65.380 0.000 65.660 4.000 ;
    END
  END prod_id[6]
  PIN prod_id[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 12.090 23.530 12.670 24.170 ;
        RECT 12.090 22.120 12.360 23.530 ;
        RECT 11.600 21.850 12.360 22.120 ;
        RECT 11.600 20.850 11.930 21.850 ;
      LAYER L1M1_PR_C ;
        RECT 11.670 21.560 11.840 21.730 ;
      LAYER met1 ;
        RECT 11.600 21.710 11.920 21.770 ;
        RECT 11.400 21.570 11.920 21.710 ;
        RECT 11.600 21.510 11.920 21.570 ;
      LAYER via ;
        RECT 11.630 21.510 11.890 21.770 ;
      LAYER met2 ;
        RECT 11.630 21.480 11.890 21.800 ;
        RECT 11.690 19.790 11.830 21.480 ;
        RECT 11.620 19.420 11.900 19.790 ;
      LAYER via2 ;
        RECT 11.620 19.470 11.900 19.750 ;
      LAYER met3 ;
        RECT 0.000 19.760 4.000 19.910 ;
        RECT 11.590 19.760 11.920 19.770 ;
        RECT 0.000 19.460 11.920 19.760 ;
        RECT 0.000 19.310 4.000 19.460 ;
        RECT 11.590 19.440 11.920 19.460 ;
    END
  END prod_id[7]
  PIN reg_ena
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 46.210 107.950 46.920 108.340 ;
        RECT 51.860 89.990 52.210 92.960 ;
      LAYER L1M1_PR_C ;
        RECT 46.230 108.140 46.400 108.310 ;
        RECT 51.990 90.380 52.160 90.550 ;
      LAYER met1 ;
        RECT 46.160 108.290 46.480 108.350 ;
        RECT 45.960 108.150 46.480 108.290 ;
        RECT 46.160 108.090 46.480 108.150 ;
        RECT 46.160 90.530 46.480 90.590 ;
        RECT 51.930 90.530 52.220 90.580 ;
        RECT 46.160 90.390 52.220 90.530 ;
        RECT 46.160 90.330 46.480 90.390 ;
        RECT 51.930 90.350 52.220 90.390 ;
        RECT 12.560 15.420 12.880 15.480 ;
        RECT 46.160 15.420 46.480 15.480 ;
        RECT 12.560 15.280 46.480 15.420 ;
        RECT 12.560 15.220 12.880 15.280 ;
        RECT 46.160 15.220 46.480 15.280 ;
      LAYER via ;
        RECT 46.190 108.090 46.450 108.350 ;
        RECT 46.190 90.330 46.450 90.590 ;
        RECT 12.590 15.220 12.850 15.480 ;
        RECT 46.190 15.220 46.450 15.480 ;
      LAYER met2 ;
        RECT 46.190 108.060 46.450 108.380 ;
        RECT 46.250 90.620 46.390 108.060 ;
        RECT 46.190 90.300 46.450 90.620 ;
        RECT 46.250 15.510 46.390 90.300 ;
        RECT 12.590 15.190 12.850 15.510 ;
        RECT 46.190 15.190 46.450 15.510 ;
        RECT 12.650 4.000 12.790 15.190 ;
        RECT 12.580 0.000 12.860 4.000 ;
    END
  END reg_ena
  PIN reset
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 83.550 83.720 83.880 83.960 ;
        RECT 74.610 78.900 75.210 79.290 ;
        RECT 76.340 73.590 76.680 76.660 ;
      LAYER L1M1_PR_C ;
        RECT 83.670 83.720 83.840 83.890 ;
        RECT 75.030 78.910 75.200 79.080 ;
        RECT 76.470 75.950 76.640 76.120 ;
      LAYER met1 ;
        RECT 55.760 151.210 56.080 151.270 ;
        RECT 75.920 151.210 76.240 151.270 ;
        RECT 55.760 151.070 76.240 151.210 ;
        RECT 55.760 151.010 56.080 151.070 ;
        RECT 75.920 151.010 76.240 151.070 ;
        RECT 75.920 86.460 76.240 86.520 ;
        RECT 83.600 86.460 83.920 86.520 ;
        RECT 75.920 86.320 83.920 86.460 ;
        RECT 75.920 86.260 76.240 86.320 ;
        RECT 83.600 86.260 83.920 86.320 ;
        RECT 83.600 83.870 83.920 83.930 ;
        RECT 83.400 83.730 83.920 83.870 ;
        RECT 83.600 83.670 83.920 83.730 ;
        RECT 74.970 79.060 75.260 79.110 ;
        RECT 75.920 79.060 76.240 79.120 ;
        RECT 74.970 78.920 76.240 79.060 ;
        RECT 74.970 78.880 75.260 78.920 ;
        RECT 75.920 78.860 76.240 78.920 ;
        RECT 75.920 76.100 76.240 76.160 ;
        RECT 76.410 76.100 76.700 76.150 ;
        RECT 75.920 75.960 76.700 76.100 ;
        RECT 75.920 75.900 76.240 75.960 ;
        RECT 76.410 75.920 76.700 75.960 ;
      LAYER via ;
        RECT 55.790 151.010 56.050 151.270 ;
        RECT 75.950 151.010 76.210 151.270 ;
        RECT 75.950 86.260 76.210 86.520 ;
        RECT 83.630 86.260 83.890 86.520 ;
        RECT 83.630 83.670 83.890 83.930 ;
        RECT 75.950 78.860 76.210 79.120 ;
        RECT 75.950 75.900 76.210 76.160 ;
      LAYER met2 ;
        RECT 55.780 165.200 56.060 169.200 ;
        RECT 55.850 151.300 55.990 165.200 ;
        RECT 55.790 150.980 56.050 151.300 ;
        RECT 75.950 150.980 76.210 151.300 ;
        RECT 76.010 86.550 76.150 150.980 ;
        RECT 75.950 86.230 76.210 86.550 ;
        RECT 83.630 86.230 83.890 86.550 ;
        RECT 76.010 79.150 76.150 86.230 ;
        RECT 83.690 83.960 83.830 86.230 ;
        RECT 83.630 83.640 83.890 83.960 ;
        RECT 75.950 78.830 76.210 79.150 ;
        RECT 76.010 76.190 76.150 78.830 ;
        RECT 75.950 75.870 76.210 76.190 ;
    END
  END reset
  PIN sdo_enb
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 125.780 98.130 126.130 101.100 ;
      LAYER L1M1_PR_C ;
        RECT 125.910 100.370 126.080 100.540 ;
      LAYER met1 ;
        RECT 125.840 100.520 126.160 100.580 ;
        RECT 125.640 100.380 126.160 100.520 ;
        RECT 125.840 100.320 126.160 100.380 ;
      LAYER via ;
        RECT 125.870 100.320 126.130 100.580 ;
      LAYER met2 ;
        RECT 125.860 123.020 126.140 123.390 ;
        RECT 125.930 100.610 126.070 123.020 ;
        RECT 125.870 100.290 126.130 100.610 ;
      LAYER via2 ;
        RECT 125.860 123.070 126.140 123.350 ;
      LAYER met3 ;
        RECT 125.830 123.360 126.160 123.370 ;
        RECT 144.160 123.360 148.160 123.510 ;
        RECT 125.830 123.060 148.160 123.360 ;
        RECT 125.830 123.040 126.160 123.060 ;
        RECT 144.160 122.910 148.160 123.060 ;
    END
  END sdo_enb
  PIN trap
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 78.370 70.700 78.720 70.940 ;
      LAYER L1M1_PR_C ;
        RECT 78.390 70.770 78.560 70.940 ;
      LAYER met1 ;
        RECT 77.360 70.920 77.680 70.980 ;
        RECT 78.330 70.920 78.620 70.970 ;
        RECT 77.360 70.780 78.620 70.920 ;
        RECT 77.360 70.720 77.680 70.780 ;
        RECT 78.330 70.740 78.620 70.780 ;
        RECT 2.960 19.120 3.280 19.180 ;
        RECT 26.960 19.120 27.280 19.180 ;
        RECT 2.960 18.980 27.280 19.120 ;
        RECT 2.960 18.920 3.280 18.980 ;
        RECT 26.960 18.920 27.280 18.980 ;
        RECT 26.960 15.790 27.280 15.850 ;
        RECT 40.880 15.790 41.200 15.850 ;
        RECT 26.960 15.650 41.200 15.790 ;
        RECT 26.960 15.590 27.280 15.650 ;
        RECT 40.880 15.590 41.200 15.650 ;
        RECT 77.360 14.680 77.680 14.740 ;
        RECT 45.290 14.540 77.680 14.680 ;
        RECT 40.880 14.310 41.200 14.370 ;
        RECT 45.290 14.310 45.430 14.540 ;
        RECT 77.360 14.480 77.680 14.540 ;
        RECT 40.880 14.170 45.430 14.310 ;
        RECT 40.880 14.110 41.200 14.170 ;
      LAYER via ;
        RECT 77.390 70.720 77.650 70.980 ;
        RECT 2.990 18.920 3.250 19.180 ;
        RECT 26.990 18.920 27.250 19.180 ;
        RECT 26.990 15.590 27.250 15.850 ;
        RECT 40.910 15.590 41.170 15.850 ;
        RECT 40.910 14.110 41.170 14.370 ;
        RECT 77.390 14.480 77.650 14.740 ;
      LAYER met2 ;
        RECT 77.390 70.690 77.650 71.010 ;
        RECT 2.990 18.890 3.250 19.210 ;
        RECT 26.990 18.890 27.250 19.210 ;
        RECT 3.050 4.000 3.190 18.890 ;
        RECT 27.050 15.880 27.190 18.890 ;
        RECT 26.990 15.560 27.250 15.880 ;
        RECT 40.910 15.560 41.170 15.880 ;
        RECT 40.970 14.400 41.110 15.560 ;
        RECT 77.450 14.770 77.590 70.690 ;
        RECT 77.390 14.450 77.650 14.770 ;
        RECT 40.910 14.080 41.170 14.400 ;
        RECT 2.980 0.000 3.260 4.000 ;
    END
  END trap
  PIN xtal_ena
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 32.660 143.100 33.010 146.070 ;
        RECT 35.170 135.860 35.880 136.250 ;
      LAYER L1M1_PR_C ;
        RECT 32.790 145.510 32.960 145.680 ;
        RECT 35.190 135.890 35.360 136.060 ;
      LAYER met1 ;
        RECT 21.200 145.660 21.520 145.720 ;
        RECT 32.730 145.660 33.020 145.710 ;
        RECT 35.120 145.660 35.440 145.720 ;
        RECT 21.200 145.520 35.440 145.660 ;
        RECT 21.200 145.460 21.520 145.520 ;
        RECT 32.730 145.480 33.020 145.520 ;
        RECT 35.120 145.460 35.440 145.520 ;
        RECT 35.120 136.040 35.440 136.100 ;
        RECT 34.920 135.900 35.440 136.040 ;
        RECT 35.120 135.840 35.440 135.900 ;
      LAYER via ;
        RECT 21.230 145.460 21.490 145.720 ;
        RECT 35.150 145.460 35.410 145.720 ;
        RECT 35.150 135.840 35.410 136.100 ;
      LAYER met2 ;
        RECT 21.220 149.660 21.500 150.030 ;
        RECT 21.290 145.750 21.430 149.660 ;
        RECT 21.230 145.430 21.490 145.750 ;
        RECT 35.150 145.430 35.410 145.750 ;
        RECT 35.210 136.130 35.350 145.430 ;
        RECT 35.150 135.810 35.410 136.130 ;
      LAYER via2 ;
        RECT 21.220 149.710 21.500 149.990 ;
      LAYER met3 ;
        RECT 0.000 150.000 4.000 150.150 ;
        RECT 21.190 150.000 21.520 150.010 ;
        RECT 0.000 149.700 21.520 150.000 ;
        RECT 0.000 149.550 4.000 149.700 ;
        RECT 21.190 149.680 21.520 149.700 ;
    END
  END xtal_ena
  PIN VPWR
    DIRECTION INOUT ;
    PORT
      LAYER li1 ;
        RECT 6.470 146.860 6.640 147.030 ;
        RECT 6.910 146.860 7.080 147.030 ;
        RECT 7.320 146.860 7.490 147.030 ;
        RECT 7.750 146.860 7.920 147.030 ;
        RECT 8.190 146.860 8.360 147.030 ;
        RECT 8.600 146.860 8.770 147.030 ;
        RECT 10.310 146.860 10.480 147.030 ;
        RECT 10.750 146.860 10.920 147.030 ;
        RECT 11.160 146.860 11.330 147.030 ;
        RECT 11.590 146.860 11.760 147.030 ;
        RECT 12.030 146.860 12.200 147.030 ;
        RECT 12.440 146.860 12.610 147.030 ;
        RECT 14.150 146.860 14.320 147.030 ;
        RECT 14.590 146.860 14.760 147.030 ;
        RECT 15.000 146.860 15.170 147.030 ;
        RECT 15.430 146.860 15.600 147.030 ;
        RECT 15.870 146.860 16.040 147.030 ;
        RECT 16.280 146.860 16.450 147.030 ;
        RECT 17.990 146.860 18.160 147.030 ;
        RECT 18.430 146.860 18.600 147.030 ;
        RECT 18.840 146.860 19.010 147.030 ;
        RECT 19.270 146.860 19.440 147.030 ;
        RECT 19.710 146.860 19.880 147.030 ;
        RECT 20.120 146.860 20.290 147.030 ;
        RECT 22.360 146.910 22.530 147.080 ;
        RECT 22.720 146.910 22.890 147.080 ;
        RECT 25.190 146.860 25.360 147.030 ;
        RECT 25.630 146.860 25.800 147.030 ;
        RECT 26.040 146.860 26.210 147.030 ;
        RECT 26.470 146.860 26.640 147.030 ;
        RECT 26.910 146.860 27.080 147.030 ;
        RECT 27.320 146.860 27.490 147.030 ;
        RECT 29.030 146.860 29.200 147.030 ;
        RECT 29.470 146.860 29.640 147.030 ;
        RECT 29.880 146.860 30.050 147.030 ;
        RECT 30.310 146.860 30.480 147.030 ;
        RECT 30.750 146.860 30.920 147.030 ;
        RECT 31.160 146.860 31.330 147.030 ;
        RECT 32.870 146.860 33.040 147.030 ;
        RECT 33.310 146.860 33.480 147.030 ;
        RECT 33.720 146.860 33.890 147.030 ;
        RECT 34.150 146.860 34.320 147.030 ;
        RECT 34.590 146.860 34.760 147.030 ;
        RECT 35.000 146.860 35.170 147.030 ;
        RECT 36.710 146.860 36.880 147.030 ;
        RECT 37.150 146.860 37.320 147.030 ;
        RECT 37.560 146.860 37.730 147.030 ;
        RECT 37.990 146.860 38.160 147.030 ;
        RECT 38.430 146.860 38.600 147.030 ;
        RECT 38.840 146.860 39.010 147.030 ;
        RECT 40.550 146.860 40.720 147.030 ;
        RECT 40.990 146.860 41.160 147.030 ;
        RECT 41.400 146.860 41.570 147.030 ;
        RECT 41.830 146.860 42.000 147.030 ;
        RECT 42.270 146.860 42.440 147.030 ;
        RECT 42.680 146.860 42.850 147.030 ;
        RECT 44.390 146.860 44.560 147.030 ;
        RECT 44.830 146.860 45.000 147.030 ;
        RECT 45.240 146.860 45.410 147.030 ;
        RECT 45.670 146.860 45.840 147.030 ;
        RECT 46.110 146.860 46.280 147.030 ;
        RECT 46.520 146.860 46.690 147.030 ;
        RECT 48.230 146.860 48.400 147.030 ;
        RECT 48.670 146.860 48.840 147.030 ;
        RECT 49.080 146.860 49.250 147.030 ;
        RECT 49.510 146.860 49.680 147.030 ;
        RECT 49.950 146.860 50.120 147.030 ;
        RECT 50.360 146.860 50.530 147.030 ;
        RECT 52.070 146.860 52.240 147.030 ;
        RECT 52.510 146.860 52.680 147.030 ;
        RECT 52.920 146.860 53.090 147.030 ;
        RECT 53.350 146.860 53.520 147.030 ;
        RECT 53.790 146.860 53.960 147.030 ;
        RECT 54.200 146.860 54.370 147.030 ;
        RECT 55.910 146.860 56.080 147.030 ;
        RECT 56.350 146.860 56.520 147.030 ;
        RECT 56.760 146.860 56.930 147.030 ;
        RECT 57.190 146.860 57.360 147.030 ;
        RECT 57.630 146.860 57.800 147.030 ;
        RECT 58.040 146.860 58.210 147.030 ;
        RECT 59.750 146.860 59.920 147.030 ;
        RECT 60.190 146.860 60.360 147.030 ;
        RECT 60.600 146.860 60.770 147.030 ;
        RECT 61.030 146.860 61.200 147.030 ;
        RECT 61.470 146.860 61.640 147.030 ;
        RECT 61.880 146.860 62.050 147.030 ;
        RECT 63.380 146.860 63.550 147.030 ;
        RECT 63.740 146.860 63.910 147.030 ;
        RECT 64.180 146.860 64.350 147.030 ;
        RECT 65.080 146.910 65.250 147.080 ;
        RECT 65.440 146.910 65.610 147.080 ;
        RECT 67.910 146.860 68.080 147.030 ;
        RECT 68.350 146.860 68.520 147.030 ;
        RECT 68.760 146.860 68.930 147.030 ;
        RECT 69.190 146.860 69.360 147.030 ;
        RECT 69.630 146.860 69.800 147.030 ;
        RECT 70.040 146.860 70.210 147.030 ;
        RECT 71.750 146.860 71.920 147.030 ;
        RECT 72.190 146.860 72.360 147.030 ;
        RECT 72.600 146.860 72.770 147.030 ;
        RECT 73.030 146.860 73.200 147.030 ;
        RECT 73.470 146.860 73.640 147.030 ;
        RECT 73.880 146.860 74.050 147.030 ;
        RECT 75.160 146.910 75.330 147.080 ;
        RECT 75.520 146.910 75.690 147.080 ;
        RECT 77.990 146.860 78.160 147.030 ;
        RECT 78.430 146.860 78.600 147.030 ;
        RECT 78.840 146.860 79.010 147.030 ;
        RECT 79.270 146.860 79.440 147.030 ;
        RECT 79.710 146.860 79.880 147.030 ;
        RECT 80.120 146.860 80.290 147.030 ;
        RECT 81.830 146.860 82.000 147.030 ;
        RECT 82.270 146.860 82.440 147.030 ;
        RECT 82.680 146.860 82.850 147.030 ;
        RECT 83.110 146.860 83.280 147.030 ;
        RECT 83.550 146.860 83.720 147.030 ;
        RECT 83.960 146.860 84.130 147.030 ;
        RECT 85.670 146.860 85.840 147.030 ;
        RECT 86.110 146.860 86.280 147.030 ;
        RECT 86.520 146.860 86.690 147.030 ;
        RECT 86.950 146.860 87.120 147.030 ;
        RECT 87.390 146.860 87.560 147.030 ;
        RECT 87.800 146.860 87.970 147.030 ;
        RECT 89.510 146.860 89.680 147.030 ;
        RECT 89.950 146.860 90.120 147.030 ;
        RECT 90.360 146.860 90.530 147.030 ;
        RECT 90.790 146.860 90.960 147.030 ;
        RECT 91.230 146.860 91.400 147.030 ;
        RECT 91.640 146.860 91.810 147.030 ;
        RECT 93.350 146.860 93.520 147.030 ;
        RECT 93.790 146.860 93.960 147.030 ;
        RECT 94.200 146.860 94.370 147.030 ;
        RECT 94.630 146.860 94.800 147.030 ;
        RECT 95.070 146.860 95.240 147.030 ;
        RECT 95.480 146.860 95.650 147.030 ;
        RECT 97.190 146.860 97.360 147.030 ;
        RECT 97.630 146.860 97.800 147.030 ;
        RECT 98.040 146.860 98.210 147.030 ;
        RECT 98.470 146.860 98.640 147.030 ;
        RECT 98.910 146.860 99.080 147.030 ;
        RECT 99.320 146.860 99.490 147.030 ;
        RECT 101.030 146.860 101.200 147.030 ;
        RECT 101.470 146.860 101.640 147.030 ;
        RECT 101.880 146.860 102.050 147.030 ;
        RECT 102.310 146.860 102.480 147.030 ;
        RECT 102.750 146.860 102.920 147.030 ;
        RECT 103.160 146.860 103.330 147.030 ;
        RECT 104.870 146.860 105.040 147.030 ;
        RECT 105.310 146.860 105.480 147.030 ;
        RECT 105.720 146.860 105.890 147.030 ;
        RECT 106.150 146.860 106.320 147.030 ;
        RECT 106.590 146.860 106.760 147.030 ;
        RECT 107.000 146.860 107.170 147.030 ;
        RECT 108.710 146.860 108.880 147.030 ;
        RECT 109.150 146.860 109.320 147.030 ;
        RECT 109.560 146.860 109.730 147.030 ;
        RECT 109.990 146.860 110.160 147.030 ;
        RECT 110.430 146.860 110.600 147.030 ;
        RECT 110.840 146.860 111.010 147.030 ;
        RECT 112.550 146.860 112.720 147.030 ;
        RECT 112.990 146.860 113.160 147.030 ;
        RECT 113.400 146.860 113.570 147.030 ;
        RECT 113.830 146.860 114.000 147.030 ;
        RECT 114.270 146.860 114.440 147.030 ;
        RECT 114.680 146.860 114.850 147.030 ;
        RECT 116.390 146.860 116.560 147.030 ;
        RECT 116.830 146.860 117.000 147.030 ;
        RECT 117.240 146.860 117.410 147.030 ;
        RECT 117.670 146.860 117.840 147.030 ;
        RECT 118.110 146.860 118.280 147.030 ;
        RECT 118.520 146.860 118.690 147.030 ;
        RECT 120.230 146.860 120.400 147.030 ;
        RECT 120.670 146.860 120.840 147.030 ;
        RECT 121.080 146.860 121.250 147.030 ;
        RECT 121.510 146.860 121.680 147.030 ;
        RECT 121.950 146.860 122.120 147.030 ;
        RECT 122.360 146.860 122.530 147.030 ;
        RECT 124.070 146.860 124.240 147.030 ;
        RECT 124.510 146.860 124.680 147.030 ;
        RECT 124.920 146.860 125.090 147.030 ;
        RECT 125.350 146.860 125.520 147.030 ;
        RECT 125.790 146.860 125.960 147.030 ;
        RECT 126.200 146.860 126.370 147.030 ;
        RECT 127.910 146.860 128.080 147.030 ;
        RECT 128.350 146.860 128.520 147.030 ;
        RECT 128.760 146.860 128.930 147.030 ;
        RECT 129.190 146.860 129.360 147.030 ;
        RECT 129.630 146.860 129.800 147.030 ;
        RECT 130.040 146.860 130.210 147.030 ;
        RECT 131.750 146.860 131.920 147.030 ;
        RECT 132.190 146.860 132.360 147.030 ;
        RECT 132.600 146.860 132.770 147.030 ;
        RECT 133.030 146.860 133.200 147.030 ;
        RECT 133.470 146.860 133.640 147.030 ;
        RECT 133.880 146.860 134.050 147.030 ;
        RECT 135.590 146.860 135.760 147.030 ;
        RECT 136.030 146.860 136.200 147.030 ;
        RECT 136.440 146.860 136.610 147.030 ;
        RECT 136.870 146.860 137.040 147.030 ;
        RECT 137.310 146.860 137.480 147.030 ;
        RECT 137.720 146.860 137.890 147.030 ;
        RECT 139.220 146.860 139.390 147.030 ;
        RECT 139.580 146.860 139.750 147.030 ;
        RECT 140.020 146.860 140.190 147.030 ;
        RECT 5.920 146.430 6.090 146.610 ;
        RECT 6.400 146.430 6.570 146.610 ;
        RECT 6.880 146.430 7.050 146.610 ;
        RECT 7.360 146.430 7.530 146.610 ;
        RECT 7.840 146.430 8.010 146.610 ;
        RECT 8.320 146.430 8.490 146.610 ;
        RECT 8.800 146.430 8.970 146.610 ;
        RECT 9.280 146.430 9.450 146.610 ;
        RECT 9.760 146.430 9.930 146.610 ;
        RECT 10.240 146.430 10.410 146.610 ;
        RECT 10.720 146.430 10.890 146.610 ;
        RECT 11.200 146.430 11.370 146.610 ;
        RECT 11.680 146.430 11.850 146.610 ;
        RECT 12.160 146.430 12.330 146.610 ;
        RECT 12.640 146.430 12.810 146.610 ;
        RECT 13.120 146.430 13.290 146.610 ;
        RECT 13.600 146.430 13.770 146.610 ;
        RECT 14.080 146.430 14.250 146.610 ;
        RECT 14.560 146.430 14.730 146.610 ;
        RECT 15.040 146.430 15.210 146.610 ;
        RECT 15.520 146.430 15.690 146.610 ;
        RECT 16.000 146.430 16.170 146.610 ;
        RECT 16.480 146.430 16.650 146.610 ;
        RECT 16.960 146.430 17.130 146.610 ;
        RECT 17.440 146.430 17.610 146.610 ;
      LAYER li1 ;
        RECT 17.760 146.600 18.240 146.610 ;
      LAYER li1 ;
        RECT 17.920 146.430 18.090 146.600 ;
        RECT 18.400 146.430 18.570 146.610 ;
        RECT 18.880 146.430 19.050 146.610 ;
        RECT 19.360 146.430 19.530 146.610 ;
        RECT 19.840 146.430 20.010 146.610 ;
        RECT 20.320 146.430 20.490 146.610 ;
        RECT 20.800 146.430 20.970 146.610 ;
        RECT 21.280 146.430 21.450 146.610 ;
        RECT 21.760 146.430 21.930 146.610 ;
        RECT 22.240 146.430 22.410 146.610 ;
        RECT 22.720 146.430 22.890 146.610 ;
        RECT 23.200 146.430 23.370 146.610 ;
        RECT 23.680 146.430 23.850 146.610 ;
        RECT 24.160 146.430 24.330 146.610 ;
        RECT 24.640 146.430 24.810 146.610 ;
        RECT 25.120 146.430 25.290 146.610 ;
        RECT 25.600 146.430 25.770 146.610 ;
        RECT 26.080 146.430 26.250 146.610 ;
        RECT 26.560 146.430 26.730 146.610 ;
        RECT 27.040 146.430 27.210 146.610 ;
        RECT 27.520 146.430 27.690 146.610 ;
        RECT 28.000 146.430 28.170 146.610 ;
        RECT 28.480 146.430 28.650 146.610 ;
        RECT 28.960 146.430 29.130 146.610 ;
        RECT 29.440 146.430 29.610 146.610 ;
        RECT 29.920 146.430 30.090 146.610 ;
        RECT 30.400 146.430 30.570 146.610 ;
        RECT 30.880 146.430 31.050 146.610 ;
        RECT 31.360 146.430 31.530 146.610 ;
        RECT 31.840 146.430 32.010 146.610 ;
        RECT 32.320 146.430 32.490 146.610 ;
        RECT 32.800 146.430 32.970 146.610 ;
        RECT 33.280 146.430 33.450 146.610 ;
        RECT 33.760 146.430 33.930 146.610 ;
        RECT 34.240 146.430 34.410 146.610 ;
        RECT 34.720 146.430 34.890 146.610 ;
        RECT 35.200 146.430 35.370 146.610 ;
        RECT 35.680 146.430 35.850 146.610 ;
      LAYER li1 ;
        RECT 36.000 146.600 36.480 146.610 ;
      LAYER li1 ;
        RECT 36.160 146.430 36.330 146.600 ;
        RECT 36.640 146.430 36.810 146.610 ;
        RECT 37.120 146.430 37.290 146.610 ;
        RECT 37.600 146.430 37.770 146.610 ;
        RECT 38.080 146.430 38.250 146.610 ;
        RECT 38.560 146.430 38.730 146.610 ;
        RECT 39.040 146.430 39.210 146.610 ;
        RECT 39.520 146.430 39.690 146.610 ;
        RECT 40.000 146.430 40.170 146.610 ;
        RECT 40.480 146.430 40.650 146.610 ;
        RECT 40.960 146.430 41.130 146.610 ;
        RECT 41.440 146.430 41.610 146.610 ;
        RECT 41.920 146.430 42.090 146.610 ;
        RECT 42.400 146.430 42.570 146.610 ;
        RECT 42.880 146.430 43.050 146.610 ;
        RECT 43.360 146.430 43.530 146.610 ;
      LAYER li1 ;
        RECT 43.680 146.600 44.160 146.610 ;
      LAYER li1 ;
        RECT 43.840 146.430 44.010 146.600 ;
        RECT 44.320 146.430 44.490 146.610 ;
        RECT 44.800 146.430 44.970 146.610 ;
        RECT 45.280 146.430 45.450 146.610 ;
        RECT 45.760 146.430 45.930 146.610 ;
        RECT 46.240 146.430 46.410 146.610 ;
        RECT 46.720 146.430 46.890 146.610 ;
        RECT 47.200 146.430 47.370 146.610 ;
        RECT 47.680 146.430 47.850 146.610 ;
        RECT 48.160 146.430 48.330 146.610 ;
        RECT 48.640 146.430 48.810 146.610 ;
        RECT 49.120 146.430 49.290 146.610 ;
        RECT 49.600 146.430 49.770 146.610 ;
        RECT 50.080 146.430 50.250 146.610 ;
        RECT 50.560 146.430 50.730 146.610 ;
        RECT 51.040 146.430 51.210 146.610 ;
        RECT 51.520 146.430 51.690 146.610 ;
        RECT 52.000 146.430 52.170 146.610 ;
        RECT 52.480 146.430 52.650 146.610 ;
        RECT 52.960 146.430 53.130 146.610 ;
        RECT 53.440 146.430 53.610 146.610 ;
        RECT 53.920 146.430 54.090 146.610 ;
        RECT 54.400 146.430 54.570 146.610 ;
        RECT 54.880 146.430 55.050 146.610 ;
        RECT 55.360 146.430 55.530 146.610 ;
        RECT 55.840 146.430 56.010 146.610 ;
        RECT 56.320 146.430 56.490 146.610 ;
        RECT 56.800 146.430 56.970 146.610 ;
        RECT 57.280 146.430 57.450 146.610 ;
        RECT 57.760 146.430 57.930 146.610 ;
        RECT 58.240 146.430 58.410 146.610 ;
        RECT 58.720 146.430 58.890 146.610 ;
        RECT 59.200 146.430 59.370 146.610 ;
        RECT 59.680 146.430 59.850 146.610 ;
        RECT 60.160 146.430 60.330 146.610 ;
        RECT 60.640 146.430 60.810 146.610 ;
        RECT 61.120 146.430 61.290 146.610 ;
        RECT 61.600 146.430 61.770 146.610 ;
        RECT 62.080 146.430 62.250 146.610 ;
        RECT 62.560 146.430 62.730 146.610 ;
        RECT 63.040 146.430 63.210 146.610 ;
        RECT 63.520 146.430 63.690 146.610 ;
        RECT 64.000 146.430 64.170 146.610 ;
        RECT 64.480 146.430 64.650 146.610 ;
        RECT 64.960 146.430 65.130 146.610 ;
        RECT 65.440 146.430 65.610 146.610 ;
        RECT 65.920 146.430 66.090 146.610 ;
        RECT 66.400 146.430 66.570 146.610 ;
        RECT 66.880 146.430 67.050 146.610 ;
        RECT 67.360 146.430 67.530 146.610 ;
        RECT 67.840 146.430 68.010 146.610 ;
        RECT 68.320 146.430 68.490 146.610 ;
        RECT 68.800 146.430 68.970 146.610 ;
        RECT 69.280 146.430 69.450 146.610 ;
        RECT 69.760 146.430 69.930 146.610 ;
        RECT 70.240 146.430 70.410 146.610 ;
        RECT 70.720 146.430 70.890 146.610 ;
        RECT 71.200 146.430 71.370 146.610 ;
        RECT 71.680 146.430 71.850 146.610 ;
        RECT 72.160 146.430 72.330 146.610 ;
        RECT 72.640 146.430 72.810 146.610 ;
        RECT 73.120 146.430 73.290 146.610 ;
        RECT 73.600 146.430 73.770 146.610 ;
        RECT 74.080 146.430 74.250 146.610 ;
        RECT 74.560 146.430 74.730 146.610 ;
        RECT 75.040 146.430 75.210 146.610 ;
        RECT 75.520 146.430 75.690 146.610 ;
        RECT 76.000 146.430 76.170 146.610 ;
        RECT 76.480 146.430 76.650 146.610 ;
        RECT 76.960 146.430 77.130 146.610 ;
        RECT 77.440 146.430 77.610 146.610 ;
        RECT 77.920 146.430 78.090 146.610 ;
        RECT 78.400 146.430 78.570 146.610 ;
        RECT 78.880 146.430 79.050 146.610 ;
        RECT 79.360 146.430 79.530 146.610 ;
        RECT 79.840 146.430 80.010 146.610 ;
        RECT 80.320 146.430 80.490 146.610 ;
        RECT 80.800 146.430 80.970 146.610 ;
        RECT 81.280 146.430 81.450 146.610 ;
        RECT 81.760 146.430 81.930 146.610 ;
        RECT 82.240 146.430 82.410 146.610 ;
        RECT 82.720 146.430 82.890 146.610 ;
        RECT 83.200 146.430 83.370 146.610 ;
        RECT 83.680 146.430 83.850 146.610 ;
        RECT 84.160 146.430 84.330 146.610 ;
        RECT 84.640 146.430 84.810 146.610 ;
        RECT 85.120 146.430 85.290 146.610 ;
      LAYER li1 ;
        RECT 85.440 146.600 85.920 146.610 ;
      LAYER li1 ;
        RECT 85.600 146.430 85.770 146.600 ;
        RECT 86.080 146.430 86.250 146.610 ;
        RECT 86.560 146.430 86.730 146.610 ;
        RECT 87.040 146.430 87.210 146.610 ;
        RECT 87.520 146.430 87.690 146.610 ;
        RECT 88.000 146.430 88.170 146.610 ;
        RECT 88.480 146.430 88.650 146.610 ;
        RECT 88.960 146.430 89.130 146.610 ;
        RECT 89.440 146.430 89.610 146.610 ;
        RECT 89.920 146.430 90.090 146.610 ;
        RECT 90.400 146.430 90.570 146.610 ;
        RECT 90.880 146.430 91.050 146.610 ;
        RECT 91.360 146.430 91.530 146.610 ;
        RECT 91.840 146.430 92.010 146.610 ;
        RECT 92.320 146.430 92.490 146.610 ;
        RECT 92.800 146.430 92.970 146.610 ;
        RECT 93.280 146.430 93.450 146.610 ;
        RECT 93.760 146.430 93.930 146.610 ;
        RECT 94.240 146.430 94.410 146.610 ;
        RECT 94.720 146.430 94.890 146.610 ;
        RECT 95.200 146.430 95.370 146.610 ;
        RECT 95.680 146.430 95.850 146.610 ;
        RECT 96.160 146.430 96.330 146.610 ;
        RECT 96.640 146.430 96.810 146.610 ;
        RECT 97.120 146.430 97.290 146.610 ;
        RECT 97.600 146.430 97.770 146.610 ;
        RECT 98.080 146.430 98.250 146.610 ;
        RECT 98.560 146.430 98.730 146.610 ;
        RECT 99.040 146.430 99.210 146.610 ;
        RECT 99.520 146.430 99.690 146.610 ;
        RECT 100.000 146.430 100.170 146.610 ;
        RECT 100.480 146.430 100.650 146.610 ;
        RECT 100.960 146.430 101.130 146.610 ;
        RECT 101.440 146.430 101.610 146.610 ;
        RECT 101.920 146.430 102.090 146.610 ;
        RECT 102.400 146.430 102.570 146.610 ;
        RECT 102.880 146.430 103.050 146.610 ;
        RECT 103.360 146.430 103.530 146.610 ;
        RECT 103.840 146.430 104.010 146.610 ;
        RECT 104.320 146.430 104.490 146.610 ;
        RECT 104.800 146.430 104.970 146.610 ;
        RECT 105.280 146.430 105.450 146.610 ;
        RECT 105.760 146.430 105.930 146.610 ;
        RECT 106.240 146.430 106.410 146.610 ;
        RECT 106.720 146.430 106.890 146.610 ;
        RECT 107.200 146.430 107.370 146.610 ;
        RECT 107.680 146.430 107.850 146.610 ;
        RECT 108.160 146.430 108.330 146.610 ;
        RECT 108.640 146.430 108.810 146.610 ;
        RECT 109.120 146.430 109.290 146.610 ;
        RECT 109.600 146.430 109.770 146.610 ;
        RECT 110.080 146.430 110.250 146.610 ;
        RECT 110.560 146.430 110.730 146.610 ;
        RECT 111.040 146.430 111.210 146.610 ;
        RECT 111.520 146.430 111.690 146.610 ;
        RECT 112.000 146.430 112.170 146.610 ;
        RECT 112.480 146.430 112.650 146.610 ;
        RECT 112.960 146.430 113.130 146.610 ;
        RECT 113.440 146.430 113.610 146.610 ;
        RECT 113.920 146.430 114.090 146.610 ;
        RECT 114.400 146.430 114.570 146.610 ;
        RECT 114.880 146.430 115.050 146.610 ;
        RECT 115.360 146.430 115.530 146.610 ;
        RECT 115.840 146.430 116.010 146.610 ;
        RECT 116.320 146.430 116.490 146.610 ;
        RECT 116.800 146.430 116.970 146.610 ;
        RECT 117.280 146.430 117.450 146.610 ;
        RECT 117.760 146.430 117.930 146.610 ;
        RECT 118.240 146.430 118.410 146.610 ;
        RECT 118.720 146.430 118.890 146.610 ;
        RECT 119.200 146.430 119.370 146.610 ;
        RECT 119.680 146.430 119.850 146.610 ;
        RECT 120.160 146.430 120.330 146.610 ;
        RECT 120.640 146.430 120.810 146.610 ;
        RECT 121.120 146.430 121.290 146.610 ;
        RECT 121.600 146.430 121.770 146.610 ;
        RECT 122.080 146.430 122.250 146.610 ;
        RECT 122.560 146.430 122.730 146.610 ;
        RECT 123.040 146.430 123.210 146.610 ;
        RECT 123.520 146.430 123.690 146.610 ;
        RECT 124.000 146.430 124.170 146.610 ;
        RECT 124.480 146.430 124.650 146.610 ;
        RECT 124.960 146.430 125.130 146.610 ;
        RECT 125.440 146.430 125.610 146.610 ;
        RECT 125.920 146.430 126.090 146.610 ;
        RECT 126.400 146.430 126.570 146.610 ;
        RECT 126.880 146.430 127.050 146.610 ;
        RECT 127.360 146.430 127.530 146.610 ;
        RECT 127.840 146.430 128.010 146.610 ;
        RECT 128.320 146.430 128.490 146.610 ;
        RECT 128.800 146.430 128.970 146.610 ;
        RECT 129.280 146.430 129.450 146.610 ;
        RECT 129.760 146.430 129.930 146.610 ;
        RECT 130.240 146.430 130.410 146.610 ;
        RECT 130.720 146.430 130.890 146.610 ;
        RECT 131.200 146.430 131.370 146.610 ;
        RECT 131.680 146.430 131.850 146.610 ;
        RECT 132.160 146.430 132.330 146.610 ;
        RECT 132.640 146.430 132.810 146.610 ;
        RECT 133.120 146.430 133.290 146.610 ;
        RECT 133.600 146.430 133.770 146.610 ;
        RECT 134.080 146.430 134.250 146.610 ;
        RECT 134.560 146.430 134.730 146.610 ;
        RECT 135.040 146.430 135.210 146.610 ;
        RECT 135.520 146.430 135.690 146.610 ;
        RECT 136.000 146.430 136.170 146.610 ;
        RECT 136.480 146.430 136.650 146.610 ;
        RECT 136.960 146.430 137.130 146.610 ;
        RECT 137.440 146.430 137.610 146.610 ;
        RECT 137.920 146.430 138.090 146.610 ;
        RECT 138.400 146.430 138.570 146.610 ;
        RECT 138.880 146.430 139.050 146.610 ;
        RECT 139.360 146.430 139.530 146.610 ;
        RECT 139.840 146.430 140.010 146.610 ;
        RECT 140.320 146.430 140.490 146.610 ;
        RECT 140.800 146.430 140.970 146.610 ;
        RECT 141.280 146.430 141.450 146.610 ;
      LAYER li1 ;
        RECT 141.600 146.430 142.080 146.610 ;
      LAYER li1 ;
        RECT 6.470 146.010 6.640 146.180 ;
        RECT 6.910 146.010 7.080 146.180 ;
        RECT 7.320 146.010 7.490 146.180 ;
        RECT 7.750 146.010 7.920 146.180 ;
        RECT 8.190 146.010 8.360 146.180 ;
        RECT 8.600 146.010 8.770 146.180 ;
        RECT 10.840 145.960 11.010 146.130 ;
        RECT 11.200 145.960 11.370 146.130 ;
        RECT 13.670 146.010 13.840 146.180 ;
        RECT 14.110 146.010 14.280 146.180 ;
        RECT 14.520 146.010 14.690 146.180 ;
        RECT 14.950 146.010 15.120 146.180 ;
        RECT 15.390 146.010 15.560 146.180 ;
        RECT 15.800 146.010 15.970 146.180 ;
        RECT 18.820 145.960 18.990 146.130 ;
        RECT 19.180 145.960 19.350 146.130 ;
        RECT 19.540 145.960 19.710 146.130 ;
        RECT 20.510 145.960 20.680 146.130 ;
        RECT 23.880 145.960 24.050 146.130 ;
        RECT 25.350 145.960 25.520 146.130 ;
        RECT 25.710 145.960 25.880 146.130 ;
        RECT 26.070 145.960 26.240 146.130 ;
        RECT 28.280 145.960 28.450 146.130 ;
        RECT 28.640 145.960 28.810 146.130 ;
        RECT 29.000 145.960 29.170 146.130 ;
        RECT 30.000 145.960 30.170 146.130 ;
        RECT 30.360 145.960 30.530 146.130 ;
        RECT 30.720 145.960 30.890 146.130 ;
        RECT 31.560 145.960 31.730 146.130 ;
        RECT 31.920 145.960 32.090 146.130 ;
        RECT 32.280 145.960 32.450 146.130 ;
        RECT 33.620 146.010 33.790 146.180 ;
        RECT 33.980 146.010 34.150 146.180 ;
        RECT 34.420 146.010 34.590 146.180 ;
        RECT 37.220 145.960 37.390 146.130 ;
        RECT 37.580 145.960 37.750 146.130 ;
        RECT 39.590 146.010 39.760 146.180 ;
        RECT 40.030 146.010 40.200 146.180 ;
        RECT 40.440 146.010 40.610 146.180 ;
        RECT 40.870 146.010 41.040 146.180 ;
        RECT 41.310 146.010 41.480 146.180 ;
        RECT 41.720 146.010 41.890 146.180 ;
        RECT 44.440 145.960 44.610 146.130 ;
        RECT 44.800 145.960 44.970 146.130 ;
        RECT 47.270 146.010 47.440 146.180 ;
        RECT 47.710 146.010 47.880 146.180 ;
        RECT 48.120 146.010 48.290 146.180 ;
        RECT 48.550 146.010 48.720 146.180 ;
        RECT 48.990 146.010 49.160 146.180 ;
        RECT 49.400 146.010 49.570 146.180 ;
        RECT 51.140 145.960 51.310 146.130 ;
        RECT 51.500 145.960 51.670 146.130 ;
        RECT 53.510 146.010 53.680 146.180 ;
        RECT 53.950 146.010 54.120 146.180 ;
        RECT 54.360 146.010 54.530 146.180 ;
        RECT 54.790 146.010 54.960 146.180 ;
        RECT 55.230 146.010 55.400 146.180 ;
        RECT 55.640 146.010 55.810 146.180 ;
        RECT 57.350 146.010 57.520 146.180 ;
        RECT 57.790 146.010 57.960 146.180 ;
        RECT 58.200 146.010 58.370 146.180 ;
        RECT 58.630 146.010 58.800 146.180 ;
        RECT 59.070 146.010 59.240 146.180 ;
        RECT 59.480 146.010 59.650 146.180 ;
        RECT 61.140 145.960 61.310 146.130 ;
        RECT 61.500 145.960 61.670 146.130 ;
        RECT 63.530 145.960 63.700 146.130 ;
        RECT 65.960 145.960 66.130 146.130 ;
        RECT 66.320 145.960 66.490 146.130 ;
        RECT 66.680 145.960 66.850 146.130 ;
        RECT 68.300 145.960 68.470 146.130 ;
        RECT 68.660 145.960 68.830 146.130 ;
        RECT 69.020 145.960 69.190 146.130 ;
        RECT 71.000 145.960 71.170 146.130 ;
        RECT 71.360 145.960 71.530 146.130 ;
        RECT 71.720 145.960 71.890 146.130 ;
        RECT 72.750 145.960 72.920 146.130 ;
        RECT 73.110 145.960 73.280 146.130 ;
        RECT 73.470 145.960 73.640 146.130 ;
        RECT 74.280 145.960 74.450 146.130 ;
        RECT 74.640 145.960 74.810 146.130 ;
        RECT 75.000 145.960 75.170 146.130 ;
        RECT 76.340 146.010 76.510 146.180 ;
        RECT 76.700 146.010 76.870 146.180 ;
        RECT 77.140 146.010 77.310 146.180 ;
        RECT 77.880 145.960 78.050 146.130 ;
        RECT 78.240 145.960 78.410 146.130 ;
        RECT 78.600 145.960 78.770 146.130 ;
        RECT 79.440 145.960 79.610 146.130 ;
        RECT 79.800 145.960 79.970 146.130 ;
        RECT 80.160 145.960 80.330 146.130 ;
        RECT 81.080 145.960 81.250 146.130 ;
        RECT 81.440 145.960 81.610 146.130 ;
        RECT 81.800 145.960 81.970 146.130 ;
        RECT 83.060 146.010 83.230 146.180 ;
        RECT 83.420 146.010 83.590 146.180 ;
        RECT 83.860 146.010 84.030 146.180 ;
        RECT 86.660 145.960 86.830 146.130 ;
        RECT 87.020 145.960 87.190 146.130 ;
        RECT 89.030 146.010 89.200 146.180 ;
        RECT 89.470 146.010 89.640 146.180 ;
        RECT 89.880 146.010 90.050 146.180 ;
        RECT 90.310 146.010 90.480 146.180 ;
        RECT 90.750 146.010 90.920 146.180 ;
        RECT 91.160 146.010 91.330 146.180 ;
        RECT 92.870 146.010 93.040 146.180 ;
        RECT 93.310 146.010 93.480 146.180 ;
        RECT 93.720 146.010 93.890 146.180 ;
        RECT 94.150 146.010 94.320 146.180 ;
        RECT 94.590 146.010 94.760 146.180 ;
        RECT 95.000 146.010 95.170 146.180 ;
        RECT 96.500 146.010 96.670 146.180 ;
        RECT 96.860 146.010 97.030 146.180 ;
        RECT 97.300 146.010 97.470 146.180 ;
        RECT 98.660 145.960 98.830 146.130 ;
        RECT 99.020 145.960 99.190 146.130 ;
        RECT 100.820 146.010 100.990 146.180 ;
        RECT 101.180 146.010 101.350 146.180 ;
        RECT 101.620 146.010 101.790 146.180 ;
        RECT 102.980 145.960 103.150 146.130 ;
        RECT 103.340 145.960 103.510 146.130 ;
        RECT 105.140 146.010 105.310 146.180 ;
        RECT 105.500 146.010 105.670 146.180 ;
        RECT 105.940 146.010 106.110 146.180 ;
        RECT 107.300 145.960 107.470 146.130 ;
        RECT 107.660 145.960 107.830 146.130 ;
        RECT 109.670 146.010 109.840 146.180 ;
        RECT 110.110 146.010 110.280 146.180 ;
        RECT 110.520 146.010 110.690 146.180 ;
        RECT 110.950 146.010 111.120 146.180 ;
        RECT 111.390 146.010 111.560 146.180 ;
        RECT 111.800 146.010 111.970 146.180 ;
        RECT 113.510 146.010 113.680 146.180 ;
        RECT 113.950 146.010 114.120 146.180 ;
        RECT 114.360 146.010 114.530 146.180 ;
        RECT 114.790 146.010 114.960 146.180 ;
        RECT 115.230 146.010 115.400 146.180 ;
        RECT 115.640 146.010 115.810 146.180 ;
        RECT 117.350 146.010 117.520 146.180 ;
        RECT 117.790 146.010 117.960 146.180 ;
        RECT 118.200 146.010 118.370 146.180 ;
        RECT 118.630 146.010 118.800 146.180 ;
        RECT 119.070 146.010 119.240 146.180 ;
        RECT 119.480 146.010 119.650 146.180 ;
        RECT 121.190 146.010 121.360 146.180 ;
        RECT 121.630 146.010 121.800 146.180 ;
        RECT 122.040 146.010 122.210 146.180 ;
        RECT 122.470 146.010 122.640 146.180 ;
        RECT 122.910 146.010 123.080 146.180 ;
        RECT 123.320 146.010 123.490 146.180 ;
        RECT 124.820 146.010 124.990 146.180 ;
        RECT 125.180 146.010 125.350 146.180 ;
        RECT 125.620 146.010 125.790 146.180 ;
        RECT 127.480 145.960 127.650 146.130 ;
        RECT 127.840 145.960 128.010 146.130 ;
        RECT 130.310 146.010 130.480 146.180 ;
        RECT 130.750 146.010 130.920 146.180 ;
        RECT 131.160 146.010 131.330 146.180 ;
        RECT 131.590 146.010 131.760 146.180 ;
        RECT 132.030 146.010 132.200 146.180 ;
        RECT 132.440 146.010 132.610 146.180 ;
        RECT 134.180 145.960 134.350 146.130 ;
        RECT 134.540 145.960 134.710 146.130 ;
        RECT 136.550 146.010 136.720 146.180 ;
        RECT 136.990 146.010 137.160 146.180 ;
        RECT 137.400 146.010 137.570 146.180 ;
        RECT 137.830 146.010 138.000 146.180 ;
        RECT 138.270 146.010 138.440 146.180 ;
        RECT 138.680 146.010 138.850 146.180 ;
        RECT 140.180 146.010 140.350 146.180 ;
        RECT 140.540 146.010 140.710 146.180 ;
        RECT 140.980 146.010 141.150 146.180 ;
        RECT 6.470 138.720 6.640 138.890 ;
        RECT 6.910 138.720 7.080 138.890 ;
        RECT 7.320 138.720 7.490 138.890 ;
        RECT 7.750 138.720 7.920 138.890 ;
        RECT 8.190 138.720 8.360 138.890 ;
        RECT 8.600 138.720 8.770 138.890 ;
        RECT 10.310 138.720 10.480 138.890 ;
        RECT 10.750 138.720 10.920 138.890 ;
        RECT 11.160 138.720 11.330 138.890 ;
        RECT 11.590 138.720 11.760 138.890 ;
        RECT 12.030 138.720 12.200 138.890 ;
        RECT 12.440 138.720 12.610 138.890 ;
        RECT 14.150 138.720 14.320 138.890 ;
        RECT 14.590 138.720 14.760 138.890 ;
        RECT 15.000 138.720 15.170 138.890 ;
        RECT 15.430 138.720 15.600 138.890 ;
        RECT 15.870 138.720 16.040 138.890 ;
        RECT 16.280 138.720 16.450 138.890 ;
        RECT 17.990 138.720 18.160 138.890 ;
        RECT 18.430 138.720 18.600 138.890 ;
        RECT 18.840 138.720 19.010 138.890 ;
        RECT 19.270 138.720 19.440 138.890 ;
        RECT 19.710 138.720 19.880 138.890 ;
        RECT 20.120 138.720 20.290 138.890 ;
        RECT 21.830 138.720 22.000 138.890 ;
        RECT 22.270 138.720 22.440 138.890 ;
        RECT 22.680 138.720 22.850 138.890 ;
        RECT 23.110 138.720 23.280 138.890 ;
        RECT 23.550 138.720 23.720 138.890 ;
        RECT 23.960 138.720 24.130 138.890 ;
        RECT 25.670 138.720 25.840 138.890 ;
        RECT 26.110 138.720 26.280 138.890 ;
        RECT 26.520 138.720 26.690 138.890 ;
        RECT 26.950 138.720 27.120 138.890 ;
        RECT 27.390 138.720 27.560 138.890 ;
        RECT 27.800 138.720 27.970 138.890 ;
        RECT 30.900 138.770 31.070 138.940 ;
        RECT 31.260 138.770 31.430 138.940 ;
        RECT 33.290 138.770 33.460 138.940 ;
        RECT 35.720 138.770 35.890 138.940 ;
        RECT 36.080 138.770 36.250 138.940 ;
        RECT 36.440 138.770 36.610 138.940 ;
        RECT 38.060 138.770 38.230 138.940 ;
        RECT 38.420 138.770 38.590 138.940 ;
        RECT 38.780 138.770 38.950 138.940 ;
        RECT 40.760 138.770 40.930 138.940 ;
        RECT 41.120 138.770 41.290 138.940 ;
        RECT 41.480 138.770 41.650 138.940 ;
        RECT 42.510 138.770 42.680 138.940 ;
        RECT 42.870 138.770 43.040 138.940 ;
        RECT 43.230 138.770 43.400 138.940 ;
        RECT 44.040 138.770 44.210 138.940 ;
        RECT 44.400 138.770 44.570 138.940 ;
        RECT 44.760 138.770 44.930 138.940 ;
        RECT 46.100 138.720 46.270 138.890 ;
        RECT 46.460 138.720 46.630 138.890 ;
        RECT 46.900 138.720 47.070 138.890 ;
        RECT 48.180 138.770 48.350 138.940 ;
        RECT 48.540 138.770 48.710 138.940 ;
        RECT 50.570 138.770 50.740 138.940 ;
        RECT 53.000 138.770 53.170 138.940 ;
        RECT 53.360 138.770 53.530 138.940 ;
        RECT 53.720 138.770 53.890 138.940 ;
        RECT 55.340 138.770 55.510 138.940 ;
        RECT 55.700 138.770 55.870 138.940 ;
        RECT 56.060 138.770 56.230 138.940 ;
        RECT 58.040 138.770 58.210 138.940 ;
        RECT 58.400 138.770 58.570 138.940 ;
        RECT 58.760 138.770 58.930 138.940 ;
        RECT 59.790 138.770 59.960 138.940 ;
        RECT 60.150 138.770 60.320 138.940 ;
        RECT 60.510 138.770 60.680 138.940 ;
        RECT 61.320 138.770 61.490 138.940 ;
        RECT 61.680 138.770 61.850 138.940 ;
        RECT 62.040 138.770 62.210 138.940 ;
        RECT 63.380 138.720 63.550 138.890 ;
        RECT 63.740 138.720 63.910 138.890 ;
        RECT 64.180 138.720 64.350 138.890 ;
        RECT 65.540 138.770 65.710 138.940 ;
        RECT 65.900 138.770 66.070 138.940 ;
        RECT 67.910 138.720 68.080 138.890 ;
        RECT 68.350 138.720 68.520 138.890 ;
        RECT 68.760 138.720 68.930 138.890 ;
        RECT 69.190 138.720 69.360 138.890 ;
        RECT 69.630 138.720 69.800 138.890 ;
        RECT 70.040 138.720 70.210 138.890 ;
        RECT 71.160 138.770 71.330 138.940 ;
        RECT 71.520 138.770 71.690 138.940 ;
        RECT 72.980 138.720 73.150 138.890 ;
        RECT 73.340 138.720 73.510 138.890 ;
        RECT 73.780 138.720 73.950 138.890 ;
        RECT 75.140 138.770 75.310 138.940 ;
        RECT 75.500 138.770 75.670 138.940 ;
        RECT 77.300 138.720 77.470 138.890 ;
        RECT 77.660 138.720 77.830 138.890 ;
        RECT 78.100 138.720 78.270 138.890 ;
        RECT 79.380 138.770 79.550 138.940 ;
        RECT 79.740 138.770 79.910 138.940 ;
        RECT 81.770 138.770 81.940 138.940 ;
        RECT 84.200 138.770 84.370 138.940 ;
        RECT 84.560 138.770 84.730 138.940 ;
        RECT 84.920 138.770 85.090 138.940 ;
        RECT 86.540 138.770 86.710 138.940 ;
        RECT 86.900 138.770 87.070 138.940 ;
        RECT 87.260 138.770 87.430 138.940 ;
        RECT 89.240 138.770 89.410 138.940 ;
        RECT 89.600 138.770 89.770 138.940 ;
        RECT 89.960 138.770 90.130 138.940 ;
        RECT 90.990 138.770 91.160 138.940 ;
        RECT 91.350 138.770 91.520 138.940 ;
        RECT 91.710 138.770 91.880 138.940 ;
        RECT 92.520 138.770 92.690 138.940 ;
        RECT 92.880 138.770 93.050 138.940 ;
        RECT 93.240 138.770 93.410 138.940 ;
        RECT 94.790 138.720 94.960 138.890 ;
        RECT 95.230 138.720 95.400 138.890 ;
        RECT 95.640 138.720 95.810 138.890 ;
        RECT 96.070 138.720 96.240 138.890 ;
        RECT 96.510 138.720 96.680 138.890 ;
        RECT 96.920 138.720 97.090 138.890 ;
        RECT 98.580 138.770 98.750 138.940 ;
        RECT 98.940 138.770 99.110 138.940 ;
        RECT 100.970 138.770 101.140 138.940 ;
        RECT 103.400 138.770 103.570 138.940 ;
        RECT 103.760 138.770 103.930 138.940 ;
        RECT 104.120 138.770 104.290 138.940 ;
        RECT 105.740 138.770 105.910 138.940 ;
        RECT 106.100 138.770 106.270 138.940 ;
        RECT 106.460 138.770 106.630 138.940 ;
        RECT 108.440 138.770 108.610 138.940 ;
        RECT 108.800 138.770 108.970 138.940 ;
        RECT 109.160 138.770 109.330 138.940 ;
        RECT 110.190 138.770 110.360 138.940 ;
        RECT 110.550 138.770 110.720 138.940 ;
        RECT 110.910 138.770 111.080 138.940 ;
        RECT 111.720 138.770 111.890 138.940 ;
        RECT 112.080 138.770 112.250 138.940 ;
        RECT 112.440 138.770 112.610 138.940 ;
        RECT 113.990 138.720 114.160 138.890 ;
        RECT 114.430 138.720 114.600 138.890 ;
        RECT 114.840 138.720 115.010 138.890 ;
        RECT 115.270 138.720 115.440 138.890 ;
        RECT 115.710 138.720 115.880 138.890 ;
        RECT 116.120 138.720 116.290 138.890 ;
        RECT 117.830 138.720 118.000 138.890 ;
        RECT 118.270 138.720 118.440 138.890 ;
        RECT 118.680 138.720 118.850 138.890 ;
        RECT 119.110 138.720 119.280 138.890 ;
        RECT 119.550 138.720 119.720 138.890 ;
        RECT 119.960 138.720 120.130 138.890 ;
        RECT 121.670 138.720 121.840 138.890 ;
        RECT 122.110 138.720 122.280 138.890 ;
        RECT 122.520 138.720 122.690 138.890 ;
        RECT 122.950 138.720 123.120 138.890 ;
        RECT 123.390 138.720 123.560 138.890 ;
        RECT 123.800 138.720 123.970 138.890 ;
        RECT 125.510 138.720 125.680 138.890 ;
        RECT 125.950 138.720 126.120 138.890 ;
        RECT 126.360 138.720 126.530 138.890 ;
        RECT 126.790 138.720 126.960 138.890 ;
        RECT 127.230 138.720 127.400 138.890 ;
        RECT 127.640 138.720 127.810 138.890 ;
        RECT 129.350 138.720 129.520 138.890 ;
        RECT 129.790 138.720 129.960 138.890 ;
        RECT 130.200 138.720 130.370 138.890 ;
        RECT 130.630 138.720 130.800 138.890 ;
        RECT 131.070 138.720 131.240 138.890 ;
        RECT 131.480 138.720 131.650 138.890 ;
        RECT 133.190 138.720 133.360 138.890 ;
        RECT 133.630 138.720 133.800 138.890 ;
        RECT 134.040 138.720 134.210 138.890 ;
        RECT 134.470 138.720 134.640 138.890 ;
        RECT 134.910 138.720 135.080 138.890 ;
        RECT 135.320 138.720 135.490 138.890 ;
        RECT 137.030 138.720 137.200 138.890 ;
        RECT 137.470 138.720 137.640 138.890 ;
        RECT 137.880 138.720 138.050 138.890 ;
        RECT 138.310 138.720 138.480 138.890 ;
        RECT 138.750 138.720 138.920 138.890 ;
        RECT 139.160 138.720 139.330 138.890 ;
        RECT 140.660 138.720 140.830 138.890 ;
        RECT 141.020 138.720 141.190 138.890 ;
        RECT 141.460 138.720 141.630 138.890 ;
        RECT 5.920 138.290 6.090 138.470 ;
        RECT 6.400 138.290 6.570 138.470 ;
        RECT 6.880 138.290 7.050 138.470 ;
        RECT 7.360 138.290 7.530 138.470 ;
        RECT 7.840 138.290 8.010 138.470 ;
        RECT 8.320 138.290 8.490 138.470 ;
        RECT 8.800 138.290 8.970 138.470 ;
        RECT 9.280 138.290 9.450 138.470 ;
        RECT 9.760 138.290 9.930 138.470 ;
        RECT 10.240 138.290 10.410 138.470 ;
        RECT 10.720 138.290 10.890 138.470 ;
        RECT 11.200 138.290 11.370 138.470 ;
        RECT 11.680 138.290 11.850 138.470 ;
        RECT 12.160 138.290 12.330 138.470 ;
        RECT 12.640 138.290 12.810 138.470 ;
        RECT 13.120 138.290 13.290 138.470 ;
        RECT 13.600 138.290 13.770 138.470 ;
        RECT 14.080 138.290 14.250 138.470 ;
        RECT 14.560 138.290 14.730 138.470 ;
        RECT 15.040 138.290 15.210 138.470 ;
        RECT 15.520 138.290 15.690 138.470 ;
        RECT 16.000 138.290 16.170 138.470 ;
        RECT 16.480 138.290 16.650 138.470 ;
        RECT 16.960 138.290 17.130 138.470 ;
        RECT 17.440 138.290 17.610 138.470 ;
        RECT 17.920 138.290 18.090 138.470 ;
        RECT 18.400 138.290 18.570 138.470 ;
        RECT 18.880 138.290 19.050 138.470 ;
        RECT 19.360 138.290 19.530 138.470 ;
        RECT 19.840 138.290 20.010 138.470 ;
        RECT 20.320 138.290 20.490 138.470 ;
        RECT 20.800 138.290 20.970 138.470 ;
        RECT 21.280 138.290 21.450 138.470 ;
        RECT 21.760 138.290 21.930 138.470 ;
        RECT 22.240 138.290 22.410 138.470 ;
        RECT 22.720 138.290 22.890 138.470 ;
        RECT 23.200 138.290 23.370 138.470 ;
        RECT 23.680 138.290 23.850 138.470 ;
        RECT 24.160 138.290 24.330 138.470 ;
        RECT 24.640 138.290 24.810 138.470 ;
        RECT 25.120 138.290 25.290 138.470 ;
        RECT 25.600 138.290 25.770 138.470 ;
        RECT 26.080 138.290 26.250 138.470 ;
        RECT 26.560 138.290 26.730 138.470 ;
        RECT 27.040 138.290 27.210 138.470 ;
        RECT 27.520 138.290 27.690 138.470 ;
        RECT 28.000 138.290 28.170 138.470 ;
        RECT 28.480 138.290 28.650 138.470 ;
        RECT 28.960 138.290 29.130 138.470 ;
        RECT 29.440 138.290 29.610 138.470 ;
        RECT 29.920 138.460 30.090 138.470 ;
      LAYER li1 ;
        RECT 30.240 138.460 30.720 138.470 ;
        RECT 29.760 138.290 30.240 138.460 ;
      LAYER li1 ;
        RECT 30.400 138.290 30.570 138.460 ;
        RECT 30.880 138.290 31.050 138.470 ;
        RECT 31.360 138.290 31.530 138.470 ;
        RECT 31.840 138.290 32.010 138.470 ;
        RECT 32.320 138.290 32.490 138.470 ;
        RECT 32.800 138.290 32.970 138.470 ;
        RECT 33.280 138.290 33.450 138.470 ;
        RECT 33.760 138.290 33.930 138.470 ;
        RECT 34.240 138.290 34.410 138.470 ;
        RECT 34.720 138.290 34.890 138.470 ;
        RECT 35.200 138.290 35.370 138.470 ;
        RECT 35.680 138.290 35.850 138.470 ;
        RECT 36.160 138.290 36.330 138.470 ;
        RECT 36.640 138.290 36.810 138.470 ;
        RECT 37.120 138.290 37.290 138.470 ;
        RECT 37.600 138.290 37.770 138.470 ;
        RECT 38.080 138.290 38.250 138.470 ;
        RECT 38.560 138.290 38.730 138.470 ;
        RECT 39.040 138.290 39.210 138.470 ;
        RECT 39.520 138.290 39.690 138.470 ;
        RECT 40.000 138.290 40.170 138.470 ;
        RECT 40.480 138.290 40.650 138.470 ;
        RECT 40.960 138.290 41.130 138.470 ;
        RECT 41.440 138.290 41.610 138.470 ;
        RECT 41.920 138.290 42.090 138.470 ;
        RECT 42.400 138.290 42.570 138.470 ;
        RECT 42.880 138.290 43.050 138.470 ;
        RECT 43.360 138.290 43.530 138.470 ;
        RECT 43.840 138.290 44.010 138.470 ;
        RECT 44.320 138.290 44.490 138.470 ;
        RECT 44.800 138.290 44.970 138.470 ;
        RECT 45.280 138.290 45.450 138.470 ;
        RECT 45.760 138.290 45.930 138.470 ;
        RECT 46.240 138.290 46.410 138.470 ;
        RECT 46.720 138.290 46.890 138.470 ;
        RECT 47.200 138.290 47.370 138.470 ;
        RECT 47.680 138.290 47.850 138.470 ;
        RECT 48.160 138.290 48.330 138.470 ;
        RECT 48.640 138.290 48.810 138.470 ;
        RECT 49.120 138.290 49.290 138.470 ;
        RECT 49.600 138.290 49.770 138.470 ;
        RECT 50.080 138.290 50.250 138.470 ;
        RECT 50.560 138.290 50.730 138.470 ;
        RECT 51.040 138.290 51.210 138.470 ;
        RECT 51.520 138.290 51.690 138.470 ;
        RECT 52.000 138.290 52.170 138.470 ;
        RECT 52.480 138.290 52.650 138.470 ;
        RECT 52.960 138.290 53.130 138.470 ;
        RECT 53.440 138.290 53.610 138.470 ;
        RECT 53.920 138.290 54.090 138.470 ;
        RECT 54.400 138.290 54.570 138.470 ;
        RECT 54.880 138.290 55.050 138.470 ;
        RECT 55.360 138.290 55.530 138.470 ;
        RECT 55.840 138.290 56.010 138.470 ;
        RECT 56.320 138.290 56.490 138.470 ;
        RECT 56.800 138.290 56.970 138.470 ;
        RECT 57.280 138.290 57.450 138.470 ;
        RECT 57.760 138.290 57.930 138.470 ;
        RECT 58.240 138.290 58.410 138.470 ;
        RECT 58.720 138.290 58.890 138.470 ;
        RECT 59.200 138.290 59.370 138.470 ;
        RECT 59.680 138.290 59.850 138.470 ;
        RECT 60.160 138.290 60.330 138.470 ;
        RECT 60.640 138.290 60.810 138.470 ;
        RECT 61.120 138.290 61.290 138.470 ;
        RECT 61.600 138.290 61.770 138.470 ;
        RECT 62.080 138.290 62.250 138.470 ;
      LAYER li1 ;
        RECT 62.400 138.460 62.880 138.470 ;
      LAYER li1 ;
        RECT 62.560 138.290 62.730 138.460 ;
        RECT 63.040 138.290 63.210 138.470 ;
        RECT 63.520 138.290 63.690 138.470 ;
        RECT 64.000 138.290 64.170 138.470 ;
        RECT 64.480 138.290 64.650 138.470 ;
        RECT 64.960 138.290 65.130 138.470 ;
        RECT 65.440 138.290 65.610 138.470 ;
        RECT 65.920 138.290 66.090 138.470 ;
        RECT 66.400 138.290 66.570 138.470 ;
        RECT 66.880 138.290 67.050 138.470 ;
        RECT 67.360 138.290 67.530 138.470 ;
        RECT 67.840 138.290 68.010 138.470 ;
        RECT 68.320 138.290 68.490 138.470 ;
        RECT 68.800 138.290 68.970 138.470 ;
        RECT 69.280 138.290 69.450 138.470 ;
        RECT 69.760 138.290 69.930 138.470 ;
        RECT 70.240 138.290 70.410 138.470 ;
        RECT 70.720 138.290 70.890 138.470 ;
        RECT 71.200 138.290 71.370 138.470 ;
        RECT 71.680 138.290 71.850 138.470 ;
        RECT 72.160 138.290 72.330 138.470 ;
        RECT 72.640 138.290 72.810 138.470 ;
        RECT 73.120 138.290 73.290 138.470 ;
        RECT 73.600 138.290 73.770 138.470 ;
        RECT 74.080 138.290 74.250 138.470 ;
        RECT 74.560 138.290 74.730 138.470 ;
      LAYER li1 ;
        RECT 74.880 138.460 75.360 138.470 ;
      LAYER li1 ;
        RECT 75.040 138.290 75.210 138.460 ;
        RECT 75.520 138.290 75.690 138.470 ;
        RECT 76.000 138.290 76.170 138.470 ;
        RECT 76.480 138.290 76.650 138.470 ;
        RECT 76.960 138.290 77.130 138.470 ;
        RECT 77.440 138.290 77.610 138.470 ;
        RECT 77.920 138.290 78.090 138.470 ;
        RECT 78.400 138.290 78.570 138.470 ;
        RECT 78.880 138.290 79.050 138.470 ;
        RECT 79.360 138.290 79.530 138.470 ;
        RECT 79.840 138.290 80.010 138.470 ;
        RECT 80.320 138.290 80.490 138.470 ;
        RECT 80.800 138.290 80.970 138.470 ;
        RECT 81.280 138.290 81.450 138.470 ;
        RECT 81.760 138.290 81.930 138.470 ;
        RECT 82.240 138.290 82.410 138.470 ;
        RECT 82.720 138.290 82.890 138.470 ;
        RECT 83.200 138.290 83.370 138.470 ;
        RECT 83.680 138.290 83.850 138.470 ;
        RECT 84.160 138.290 84.330 138.470 ;
        RECT 84.640 138.290 84.810 138.470 ;
        RECT 85.120 138.290 85.290 138.470 ;
        RECT 85.600 138.290 85.770 138.470 ;
        RECT 86.080 138.290 86.250 138.470 ;
        RECT 86.560 138.290 86.730 138.470 ;
        RECT 87.040 138.290 87.210 138.470 ;
        RECT 87.520 138.290 87.690 138.470 ;
        RECT 88.000 138.290 88.170 138.470 ;
        RECT 88.480 138.290 88.650 138.470 ;
        RECT 88.960 138.290 89.130 138.470 ;
        RECT 89.440 138.290 89.610 138.470 ;
        RECT 89.920 138.290 90.090 138.470 ;
        RECT 90.400 138.290 90.570 138.470 ;
        RECT 90.880 138.290 91.050 138.470 ;
        RECT 91.360 138.290 91.530 138.470 ;
        RECT 91.840 138.290 92.010 138.470 ;
        RECT 92.320 138.290 92.490 138.470 ;
        RECT 92.800 138.290 92.970 138.470 ;
        RECT 93.280 138.290 93.450 138.470 ;
        RECT 93.760 138.290 93.930 138.470 ;
        RECT 94.240 138.290 94.410 138.470 ;
        RECT 94.720 138.290 94.890 138.470 ;
        RECT 95.200 138.290 95.370 138.470 ;
        RECT 95.680 138.290 95.850 138.470 ;
        RECT 96.160 138.290 96.330 138.470 ;
        RECT 96.640 138.290 96.810 138.470 ;
        RECT 97.120 138.290 97.290 138.470 ;
        RECT 97.600 138.290 97.770 138.470 ;
      LAYER li1 ;
        RECT 97.920 138.460 98.400 138.470 ;
      LAYER li1 ;
        RECT 98.080 138.290 98.250 138.460 ;
        RECT 98.560 138.290 98.730 138.470 ;
        RECT 99.040 138.290 99.210 138.470 ;
        RECT 99.520 138.290 99.690 138.470 ;
        RECT 100.000 138.290 100.170 138.470 ;
        RECT 100.480 138.290 100.650 138.470 ;
        RECT 100.960 138.290 101.130 138.470 ;
        RECT 101.440 138.290 101.610 138.470 ;
        RECT 101.920 138.290 102.090 138.470 ;
        RECT 102.400 138.290 102.570 138.470 ;
        RECT 102.880 138.290 103.050 138.470 ;
        RECT 103.360 138.290 103.530 138.470 ;
        RECT 103.840 138.290 104.010 138.470 ;
        RECT 104.320 138.290 104.490 138.470 ;
        RECT 104.800 138.290 104.970 138.470 ;
        RECT 105.280 138.290 105.450 138.470 ;
        RECT 105.760 138.290 105.930 138.470 ;
        RECT 106.240 138.290 106.410 138.470 ;
        RECT 106.720 138.290 106.890 138.470 ;
        RECT 107.200 138.290 107.370 138.470 ;
        RECT 107.680 138.290 107.850 138.470 ;
        RECT 108.160 138.290 108.330 138.470 ;
        RECT 108.640 138.290 108.810 138.470 ;
        RECT 109.120 138.290 109.290 138.470 ;
      LAYER li1 ;
        RECT 109.440 138.460 109.920 138.470 ;
      LAYER li1 ;
        RECT 109.600 138.290 109.770 138.460 ;
        RECT 110.080 138.290 110.250 138.470 ;
        RECT 110.560 138.290 110.730 138.470 ;
        RECT 111.040 138.290 111.210 138.470 ;
        RECT 111.520 138.290 111.690 138.470 ;
        RECT 112.000 138.290 112.170 138.470 ;
        RECT 112.480 138.290 112.650 138.470 ;
        RECT 112.960 138.290 113.130 138.470 ;
        RECT 113.440 138.290 113.610 138.470 ;
        RECT 113.920 138.290 114.090 138.470 ;
        RECT 114.400 138.290 114.570 138.470 ;
        RECT 114.880 138.290 115.050 138.470 ;
        RECT 115.360 138.290 115.530 138.470 ;
        RECT 115.840 138.290 116.010 138.470 ;
        RECT 116.320 138.290 116.490 138.470 ;
        RECT 116.800 138.290 116.970 138.470 ;
        RECT 117.280 138.290 117.450 138.470 ;
        RECT 117.760 138.290 117.930 138.470 ;
        RECT 118.240 138.290 118.410 138.470 ;
        RECT 118.720 138.290 118.890 138.470 ;
        RECT 119.200 138.290 119.370 138.470 ;
        RECT 119.680 138.290 119.850 138.470 ;
        RECT 120.160 138.290 120.330 138.470 ;
        RECT 120.640 138.290 120.810 138.470 ;
        RECT 121.120 138.290 121.290 138.470 ;
        RECT 121.600 138.290 121.770 138.470 ;
        RECT 122.080 138.290 122.250 138.470 ;
        RECT 122.560 138.290 122.730 138.470 ;
        RECT 123.040 138.290 123.210 138.470 ;
        RECT 123.520 138.290 123.690 138.470 ;
        RECT 124.000 138.290 124.170 138.470 ;
        RECT 124.480 138.290 124.650 138.470 ;
        RECT 124.960 138.290 125.130 138.470 ;
        RECT 125.440 138.290 125.610 138.470 ;
        RECT 125.920 138.290 126.090 138.470 ;
        RECT 126.400 138.290 126.570 138.470 ;
        RECT 126.880 138.290 127.050 138.470 ;
        RECT 127.360 138.290 127.530 138.470 ;
        RECT 127.840 138.290 128.010 138.470 ;
        RECT 128.320 138.290 128.490 138.470 ;
        RECT 128.800 138.290 128.970 138.470 ;
        RECT 129.280 138.290 129.450 138.470 ;
        RECT 129.760 138.290 129.930 138.470 ;
        RECT 130.240 138.290 130.410 138.470 ;
        RECT 130.720 138.290 130.890 138.470 ;
        RECT 131.200 138.290 131.370 138.470 ;
        RECT 131.680 138.290 131.850 138.470 ;
        RECT 132.160 138.290 132.330 138.470 ;
        RECT 132.640 138.290 132.810 138.470 ;
        RECT 133.120 138.290 133.290 138.470 ;
        RECT 133.600 138.290 133.770 138.470 ;
        RECT 134.080 138.290 134.250 138.470 ;
        RECT 134.560 138.290 134.730 138.470 ;
        RECT 135.040 138.290 135.210 138.470 ;
        RECT 135.520 138.290 135.690 138.470 ;
        RECT 136.000 138.290 136.170 138.470 ;
        RECT 136.480 138.290 136.650 138.470 ;
        RECT 136.960 138.290 137.130 138.470 ;
        RECT 137.440 138.290 137.610 138.470 ;
        RECT 137.920 138.290 138.090 138.470 ;
        RECT 138.400 138.290 138.570 138.470 ;
        RECT 138.880 138.290 139.050 138.470 ;
        RECT 139.360 138.290 139.530 138.470 ;
        RECT 139.840 138.290 140.010 138.470 ;
        RECT 140.320 138.290 140.490 138.470 ;
        RECT 140.800 138.290 140.970 138.470 ;
        RECT 141.280 138.290 141.450 138.470 ;
      LAYER li1 ;
        RECT 141.600 138.460 142.080 138.470 ;
      LAYER li1 ;
        RECT 141.760 138.290 141.930 138.460 ;
        RECT 6.470 137.870 6.640 138.040 ;
        RECT 6.910 137.870 7.080 138.040 ;
        RECT 7.320 137.870 7.490 138.040 ;
        RECT 7.750 137.870 7.920 138.040 ;
        RECT 8.190 137.870 8.360 138.040 ;
        RECT 8.600 137.870 8.770 138.040 ;
        RECT 10.100 137.870 10.270 138.040 ;
        RECT 10.460 137.870 10.630 138.040 ;
        RECT 10.900 137.870 11.070 138.040 ;
        RECT 13.220 137.820 13.390 137.990 ;
        RECT 13.580 137.820 13.750 137.990 ;
        RECT 15.590 137.870 15.760 138.040 ;
        RECT 16.030 137.870 16.200 138.040 ;
        RECT 16.440 137.870 16.610 138.040 ;
        RECT 16.870 137.870 17.040 138.040 ;
        RECT 17.310 137.870 17.480 138.040 ;
        RECT 17.720 137.870 17.890 138.040 ;
        RECT 19.430 137.870 19.600 138.040 ;
        RECT 19.870 137.870 20.040 138.040 ;
        RECT 20.280 137.870 20.450 138.040 ;
        RECT 20.710 137.870 20.880 138.040 ;
        RECT 21.150 137.870 21.320 138.040 ;
        RECT 21.560 137.870 21.730 138.040 ;
        RECT 23.270 137.870 23.440 138.040 ;
        RECT 23.710 137.870 23.880 138.040 ;
        RECT 24.120 137.870 24.290 138.040 ;
        RECT 24.550 137.870 24.720 138.040 ;
        RECT 24.990 137.870 25.160 138.040 ;
        RECT 25.400 137.870 25.570 138.040 ;
        RECT 27.110 137.870 27.280 138.040 ;
        RECT 27.550 137.870 27.720 138.040 ;
        RECT 27.960 137.870 28.130 138.040 ;
        RECT 28.390 137.870 28.560 138.040 ;
        RECT 28.830 137.870 29.000 138.040 ;
        RECT 29.240 137.870 29.410 138.040 ;
        RECT 31.460 137.820 31.630 137.990 ;
        RECT 31.820 137.820 31.990 137.990 ;
        RECT 33.620 137.870 33.790 138.040 ;
        RECT 33.980 137.870 34.150 138.040 ;
        RECT 34.420 137.870 34.590 138.040 ;
        RECT 35.160 137.820 35.330 137.990 ;
        RECT 35.520 137.820 35.690 137.990 ;
        RECT 37.190 137.870 37.360 138.040 ;
        RECT 37.630 137.870 37.800 138.040 ;
        RECT 38.040 137.870 38.210 138.040 ;
        RECT 38.470 137.870 38.640 138.040 ;
        RECT 38.910 137.870 39.080 138.040 ;
        RECT 39.320 137.870 39.490 138.040 ;
        RECT 41.030 137.870 41.200 138.040 ;
        RECT 41.470 137.870 41.640 138.040 ;
        RECT 41.880 137.870 42.050 138.040 ;
        RECT 42.310 137.870 42.480 138.040 ;
        RECT 42.750 137.870 42.920 138.040 ;
        RECT 43.160 137.870 43.330 138.040 ;
        RECT 44.870 137.870 45.040 138.040 ;
        RECT 45.310 137.870 45.480 138.040 ;
        RECT 45.720 137.870 45.890 138.040 ;
        RECT 46.150 137.870 46.320 138.040 ;
        RECT 46.590 137.870 46.760 138.040 ;
        RECT 47.000 137.870 47.170 138.040 ;
        RECT 48.710 137.870 48.880 138.040 ;
        RECT 49.150 137.870 49.320 138.040 ;
        RECT 49.560 137.870 49.730 138.040 ;
        RECT 49.990 137.870 50.160 138.040 ;
        RECT 50.430 137.870 50.600 138.040 ;
        RECT 50.840 137.870 51.010 138.040 ;
        RECT 52.550 137.870 52.720 138.040 ;
        RECT 52.990 137.870 53.160 138.040 ;
        RECT 53.400 137.870 53.570 138.040 ;
        RECT 53.830 137.870 54.000 138.040 ;
        RECT 54.270 137.870 54.440 138.040 ;
        RECT 54.680 137.870 54.850 138.040 ;
        RECT 56.390 137.870 56.560 138.040 ;
        RECT 56.830 137.870 57.000 138.040 ;
        RECT 57.240 137.870 57.410 138.040 ;
        RECT 57.670 137.870 57.840 138.040 ;
        RECT 58.110 137.870 58.280 138.040 ;
        RECT 58.520 137.870 58.690 138.040 ;
        RECT 60.020 137.870 60.190 138.040 ;
        RECT 60.380 137.870 60.550 138.040 ;
        RECT 60.820 137.870 60.990 138.040 ;
        RECT 63.000 137.820 63.170 137.990 ;
        RECT 63.360 137.820 63.530 137.990 ;
        RECT 65.030 137.870 65.200 138.040 ;
        RECT 65.470 137.870 65.640 138.040 ;
        RECT 65.880 137.870 66.050 138.040 ;
        RECT 66.310 137.870 66.480 138.040 ;
        RECT 66.750 137.870 66.920 138.040 ;
        RECT 67.160 137.870 67.330 138.040 ;
        RECT 68.870 137.870 69.040 138.040 ;
        RECT 69.310 137.870 69.480 138.040 ;
        RECT 69.720 137.870 69.890 138.040 ;
        RECT 70.150 137.870 70.320 138.040 ;
        RECT 70.590 137.870 70.760 138.040 ;
        RECT 71.000 137.870 71.170 138.040 ;
        RECT 72.500 137.870 72.670 138.040 ;
        RECT 72.860 137.870 73.030 138.040 ;
        RECT 73.300 137.870 73.470 138.040 ;
        RECT 75.460 137.820 75.630 137.990 ;
        RECT 75.820 137.820 75.990 137.990 ;
        RECT 76.180 137.820 76.350 137.990 ;
        RECT 76.540 137.820 76.710 137.990 ;
        RECT 77.700 137.820 77.870 137.990 ;
        RECT 78.060 137.820 78.230 137.990 ;
        RECT 78.420 137.820 78.590 137.990 ;
        RECT 78.780 137.820 78.950 137.990 ;
        RECT 79.910 137.870 80.080 138.040 ;
        RECT 80.350 137.870 80.520 138.040 ;
        RECT 80.760 137.870 80.930 138.040 ;
        RECT 81.190 137.870 81.360 138.040 ;
        RECT 81.630 137.870 81.800 138.040 ;
        RECT 82.040 137.870 82.210 138.040 ;
        RECT 83.750 137.870 83.920 138.040 ;
        RECT 84.190 137.870 84.360 138.040 ;
        RECT 84.600 137.870 84.770 138.040 ;
        RECT 85.030 137.870 85.200 138.040 ;
        RECT 85.470 137.870 85.640 138.040 ;
        RECT 85.880 137.870 86.050 138.040 ;
        RECT 87.440 137.820 87.610 137.990 ;
        RECT 87.800 137.820 87.970 137.990 ;
        RECT 88.160 137.820 88.330 137.990 ;
        RECT 88.520 137.820 88.690 137.990 ;
        RECT 88.880 137.820 89.050 137.990 ;
        RECT 89.240 137.820 89.410 137.990 ;
        RECT 89.600 137.820 89.770 137.990 ;
        RECT 89.960 137.820 90.130 137.990 ;
        RECT 90.770 137.820 90.940 137.990 ;
        RECT 91.130 137.820 91.300 137.990 ;
        RECT 91.490 137.820 91.660 137.990 ;
        RECT 91.850 137.820 92.020 137.990 ;
        RECT 92.870 137.870 93.040 138.040 ;
        RECT 93.310 137.870 93.480 138.040 ;
        RECT 93.720 137.870 93.890 138.040 ;
        RECT 94.150 137.870 94.320 138.040 ;
        RECT 94.590 137.870 94.760 138.040 ;
        RECT 95.000 137.870 95.170 138.040 ;
        RECT 96.500 137.870 96.670 138.040 ;
        RECT 96.860 137.870 97.030 138.040 ;
        RECT 97.300 137.870 97.470 138.040 ;
        RECT 98.960 137.820 99.130 137.990 ;
        RECT 99.320 137.820 99.490 137.990 ;
        RECT 99.680 137.820 99.850 137.990 ;
        RECT 100.040 137.820 100.210 137.990 ;
        RECT 100.400 137.820 100.570 137.990 ;
        RECT 100.760 137.820 100.930 137.990 ;
        RECT 101.120 137.820 101.290 137.990 ;
        RECT 101.480 137.820 101.650 137.990 ;
        RECT 102.290 137.820 102.460 137.990 ;
        RECT 102.650 137.820 102.820 137.990 ;
        RECT 103.010 137.820 103.180 137.990 ;
        RECT 103.370 137.820 103.540 137.990 ;
        RECT 104.390 137.870 104.560 138.040 ;
        RECT 104.830 137.870 105.000 138.040 ;
        RECT 105.240 137.870 105.410 138.040 ;
        RECT 105.670 137.870 105.840 138.040 ;
        RECT 106.110 137.870 106.280 138.040 ;
        RECT 106.520 137.870 106.690 138.040 ;
        RECT 108.020 137.870 108.190 138.040 ;
        RECT 108.380 137.870 108.550 138.040 ;
        RECT 108.820 137.870 108.990 138.040 ;
        RECT 110.660 137.820 110.830 137.990 ;
        RECT 111.020 137.820 111.190 137.990 ;
        RECT 113.030 137.870 113.200 138.040 ;
        RECT 113.470 137.870 113.640 138.040 ;
        RECT 113.880 137.870 114.050 138.040 ;
        RECT 114.310 137.870 114.480 138.040 ;
        RECT 114.750 137.870 114.920 138.040 ;
        RECT 115.160 137.870 115.330 138.040 ;
        RECT 116.660 137.870 116.830 138.040 ;
        RECT 117.020 137.870 117.190 138.040 ;
        RECT 117.460 137.870 117.630 138.040 ;
        RECT 118.820 137.820 118.990 137.990 ;
        RECT 119.180 137.820 119.350 137.990 ;
        RECT 121.190 137.870 121.360 138.040 ;
        RECT 121.630 137.870 121.800 138.040 ;
        RECT 122.040 137.870 122.210 138.040 ;
        RECT 122.470 137.870 122.640 138.040 ;
        RECT 122.910 137.870 123.080 138.040 ;
        RECT 123.320 137.870 123.490 138.040 ;
        RECT 125.030 137.870 125.200 138.040 ;
        RECT 125.470 137.870 125.640 138.040 ;
        RECT 125.880 137.870 126.050 138.040 ;
        RECT 126.310 137.870 126.480 138.040 ;
        RECT 126.750 137.870 126.920 138.040 ;
        RECT 127.160 137.870 127.330 138.040 ;
        RECT 128.870 137.870 129.040 138.040 ;
        RECT 129.310 137.870 129.480 138.040 ;
        RECT 129.720 137.870 129.890 138.040 ;
        RECT 130.150 137.870 130.320 138.040 ;
        RECT 130.590 137.870 130.760 138.040 ;
        RECT 131.000 137.870 131.170 138.040 ;
        RECT 132.710 137.870 132.880 138.040 ;
        RECT 133.150 137.870 133.320 138.040 ;
        RECT 133.560 137.870 133.730 138.040 ;
        RECT 133.990 137.870 134.160 138.040 ;
        RECT 134.430 137.870 134.600 138.040 ;
        RECT 134.840 137.870 135.010 138.040 ;
        RECT 136.550 137.870 136.720 138.040 ;
        RECT 136.990 137.870 137.160 138.040 ;
        RECT 137.400 137.870 137.570 138.040 ;
        RECT 137.830 137.870 138.000 138.040 ;
        RECT 138.270 137.870 138.440 138.040 ;
        RECT 138.680 137.870 138.850 138.040 ;
        RECT 140.180 137.870 140.350 138.040 ;
        RECT 140.540 137.870 140.710 138.040 ;
        RECT 140.980 137.870 141.150 138.040 ;
        RECT 6.470 130.580 6.640 130.750 ;
        RECT 6.910 130.580 7.080 130.750 ;
        RECT 7.320 130.580 7.490 130.750 ;
        RECT 7.750 130.580 7.920 130.750 ;
        RECT 8.190 130.580 8.360 130.750 ;
        RECT 8.600 130.580 8.770 130.750 ;
        RECT 10.840 130.630 11.010 130.800 ;
        RECT 11.200 130.630 11.370 130.800 ;
        RECT 13.670 130.580 13.840 130.750 ;
        RECT 14.110 130.580 14.280 130.750 ;
        RECT 14.520 130.580 14.690 130.750 ;
        RECT 14.950 130.580 15.120 130.750 ;
        RECT 15.390 130.580 15.560 130.750 ;
        RECT 15.800 130.580 15.970 130.750 ;
        RECT 17.510 130.580 17.680 130.750 ;
        RECT 17.950 130.580 18.120 130.750 ;
        RECT 18.360 130.580 18.530 130.750 ;
        RECT 18.790 130.580 18.960 130.750 ;
        RECT 19.230 130.580 19.400 130.750 ;
        RECT 19.640 130.580 19.810 130.750 ;
        RECT 21.350 130.580 21.520 130.750 ;
        RECT 21.790 130.580 21.960 130.750 ;
        RECT 22.200 130.580 22.370 130.750 ;
        RECT 22.630 130.580 22.800 130.750 ;
        RECT 23.070 130.580 23.240 130.750 ;
        RECT 23.480 130.580 23.650 130.750 ;
        RECT 25.190 130.580 25.360 130.750 ;
        RECT 25.630 130.580 25.800 130.750 ;
        RECT 26.040 130.580 26.210 130.750 ;
        RECT 26.470 130.580 26.640 130.750 ;
        RECT 26.910 130.580 27.080 130.750 ;
        RECT 27.320 130.580 27.490 130.750 ;
        RECT 28.820 130.580 28.990 130.750 ;
        RECT 29.180 130.580 29.350 130.750 ;
        RECT 29.620 130.580 29.790 130.750 ;
        RECT 31.780 130.630 31.950 130.800 ;
        RECT 32.140 130.630 32.310 130.800 ;
        RECT 32.500 130.630 32.670 130.800 ;
        RECT 32.860 130.630 33.030 130.800 ;
        RECT 34.020 130.630 34.190 130.800 ;
        RECT 34.380 130.630 34.550 130.800 ;
        RECT 34.740 130.630 34.910 130.800 ;
        RECT 35.100 130.630 35.270 130.800 ;
        RECT 36.230 130.580 36.400 130.750 ;
        RECT 36.670 130.580 36.840 130.750 ;
        RECT 37.080 130.580 37.250 130.750 ;
        RECT 37.510 130.580 37.680 130.750 ;
        RECT 37.950 130.580 38.120 130.750 ;
        RECT 38.360 130.580 38.530 130.750 ;
        RECT 40.070 130.580 40.240 130.750 ;
        RECT 40.510 130.580 40.680 130.750 ;
        RECT 40.920 130.580 41.090 130.750 ;
        RECT 41.350 130.580 41.520 130.750 ;
        RECT 41.790 130.580 41.960 130.750 ;
        RECT 42.200 130.580 42.370 130.750 ;
        RECT 43.910 130.580 44.080 130.750 ;
        RECT 44.350 130.580 44.520 130.750 ;
        RECT 44.760 130.580 44.930 130.750 ;
        RECT 45.190 130.580 45.360 130.750 ;
        RECT 45.630 130.580 45.800 130.750 ;
        RECT 46.040 130.580 46.210 130.750 ;
        RECT 47.750 130.580 47.920 130.750 ;
        RECT 48.190 130.580 48.360 130.750 ;
        RECT 48.600 130.580 48.770 130.750 ;
        RECT 49.030 130.580 49.200 130.750 ;
        RECT 49.470 130.580 49.640 130.750 ;
        RECT 49.880 130.580 50.050 130.750 ;
        RECT 51.590 130.580 51.760 130.750 ;
        RECT 52.030 130.580 52.200 130.750 ;
        RECT 52.440 130.580 52.610 130.750 ;
        RECT 52.870 130.580 53.040 130.750 ;
        RECT 53.310 130.580 53.480 130.750 ;
        RECT 53.720 130.580 53.890 130.750 ;
        RECT 55.430 130.580 55.600 130.750 ;
        RECT 55.870 130.580 56.040 130.750 ;
        RECT 56.280 130.580 56.450 130.750 ;
        RECT 56.710 130.580 56.880 130.750 ;
        RECT 57.150 130.580 57.320 130.750 ;
        RECT 57.560 130.580 57.730 130.750 ;
        RECT 59.270 130.580 59.440 130.750 ;
        RECT 59.710 130.580 59.880 130.750 ;
        RECT 60.120 130.580 60.290 130.750 ;
        RECT 60.550 130.580 60.720 130.750 ;
        RECT 60.990 130.580 61.160 130.750 ;
        RECT 61.400 130.580 61.570 130.750 ;
        RECT 63.110 130.580 63.280 130.750 ;
        RECT 63.550 130.580 63.720 130.750 ;
        RECT 63.960 130.580 64.130 130.750 ;
        RECT 64.390 130.580 64.560 130.750 ;
        RECT 64.830 130.580 65.000 130.750 ;
        RECT 65.240 130.580 65.410 130.750 ;
        RECT 66.950 130.580 67.120 130.750 ;
        RECT 67.390 130.580 67.560 130.750 ;
        RECT 67.800 130.580 67.970 130.750 ;
        RECT 68.230 130.580 68.400 130.750 ;
        RECT 68.670 130.580 68.840 130.750 ;
        RECT 69.080 130.580 69.250 130.750 ;
        RECT 70.580 130.580 70.750 130.750 ;
        RECT 70.940 130.580 71.110 130.750 ;
        RECT 71.380 130.580 71.550 130.750 ;
        RECT 73.550 130.630 73.720 130.800 ;
        RECT 73.910 130.630 74.080 130.800 ;
        RECT 74.270 130.630 74.440 130.800 ;
        RECT 74.990 130.630 75.160 130.800 ;
        RECT 75.350 130.630 75.520 130.800 ;
        RECT 75.710 130.630 75.880 130.800 ;
        RECT 76.070 130.630 76.240 130.800 ;
        RECT 77.300 130.580 77.470 130.750 ;
        RECT 77.660 130.580 77.830 130.750 ;
        RECT 78.100 130.580 78.270 130.750 ;
        RECT 78.840 130.630 79.010 130.800 ;
        RECT 79.200 130.630 79.370 130.800 ;
        RECT 79.560 130.630 79.730 130.800 ;
        RECT 79.920 130.630 80.090 130.800 ;
        RECT 80.280 130.630 80.450 130.800 ;
        RECT 82.580 130.580 82.750 130.750 ;
        RECT 82.940 130.580 83.110 130.750 ;
        RECT 83.380 130.580 83.550 130.750 ;
        RECT 85.520 130.630 85.690 130.800 ;
        RECT 85.880 130.630 86.050 130.800 ;
        RECT 86.240 130.630 86.410 130.800 ;
        RECT 86.600 130.630 86.770 130.800 ;
        RECT 86.960 130.630 87.130 130.800 ;
        RECT 87.320 130.630 87.490 130.800 ;
        RECT 87.680 130.630 87.850 130.800 ;
        RECT 88.040 130.630 88.210 130.800 ;
        RECT 88.850 130.630 89.020 130.800 ;
        RECT 89.210 130.630 89.380 130.800 ;
        RECT 89.570 130.630 89.740 130.800 ;
        RECT 89.930 130.630 90.100 130.800 ;
        RECT 90.950 130.580 91.120 130.750 ;
        RECT 91.390 130.580 91.560 130.750 ;
        RECT 91.800 130.580 91.970 130.750 ;
        RECT 92.230 130.580 92.400 130.750 ;
        RECT 92.670 130.580 92.840 130.750 ;
        RECT 93.080 130.580 93.250 130.750 ;
        RECT 94.790 130.580 94.960 130.750 ;
        RECT 95.230 130.580 95.400 130.750 ;
        RECT 95.640 130.580 95.810 130.750 ;
        RECT 96.070 130.580 96.240 130.750 ;
        RECT 96.510 130.580 96.680 130.750 ;
        RECT 96.920 130.580 97.090 130.750 ;
        RECT 98.480 130.630 98.650 130.800 ;
        RECT 98.840 130.630 99.010 130.800 ;
        RECT 99.200 130.630 99.370 130.800 ;
        RECT 99.560 130.630 99.730 130.800 ;
        RECT 99.920 130.630 100.090 130.800 ;
        RECT 100.280 130.630 100.450 130.800 ;
        RECT 100.640 130.630 100.810 130.800 ;
        RECT 101.000 130.630 101.170 130.800 ;
        RECT 101.810 130.630 101.980 130.800 ;
        RECT 102.170 130.630 102.340 130.800 ;
        RECT 102.530 130.630 102.700 130.800 ;
        RECT 102.890 130.630 103.060 130.800 ;
        RECT 103.700 130.580 103.870 130.750 ;
        RECT 104.060 130.580 104.230 130.750 ;
        RECT 104.500 130.580 104.670 130.750 ;
        RECT 105.240 130.630 105.410 130.800 ;
        RECT 105.600 130.630 105.770 130.800 ;
        RECT 105.960 130.630 106.130 130.800 ;
        RECT 107.370 130.630 107.540 130.800 ;
        RECT 107.730 130.630 107.900 130.800 ;
        RECT 108.090 130.630 108.260 130.800 ;
        RECT 108.980 130.580 109.150 130.750 ;
        RECT 109.340 130.580 109.510 130.750 ;
        RECT 109.780 130.580 109.950 130.750 ;
        RECT 111.540 130.630 111.710 130.800 ;
        RECT 111.900 130.630 112.070 130.800 ;
        RECT 113.930 130.630 114.100 130.800 ;
        RECT 116.360 130.630 116.530 130.800 ;
        RECT 116.720 130.630 116.890 130.800 ;
        RECT 117.080 130.630 117.250 130.800 ;
        RECT 118.700 130.630 118.870 130.800 ;
        RECT 119.060 130.630 119.230 130.800 ;
        RECT 119.420 130.630 119.590 130.800 ;
        RECT 121.400 130.630 121.570 130.800 ;
        RECT 121.760 130.630 121.930 130.800 ;
        RECT 122.120 130.630 122.290 130.800 ;
        RECT 123.150 130.630 123.320 130.800 ;
        RECT 123.510 130.630 123.680 130.800 ;
        RECT 123.870 130.630 124.040 130.800 ;
        RECT 124.680 130.630 124.850 130.800 ;
        RECT 125.040 130.630 125.210 130.800 ;
        RECT 125.400 130.630 125.570 130.800 ;
        RECT 126.950 130.580 127.120 130.750 ;
        RECT 127.390 130.580 127.560 130.750 ;
        RECT 127.800 130.580 127.970 130.750 ;
        RECT 128.230 130.580 128.400 130.750 ;
        RECT 128.670 130.580 128.840 130.750 ;
        RECT 129.080 130.580 129.250 130.750 ;
        RECT 130.790 130.580 130.960 130.750 ;
        RECT 131.230 130.580 131.400 130.750 ;
        RECT 131.640 130.580 131.810 130.750 ;
        RECT 132.070 130.580 132.240 130.750 ;
        RECT 132.510 130.580 132.680 130.750 ;
        RECT 132.920 130.580 133.090 130.750 ;
        RECT 134.630 130.580 134.800 130.750 ;
        RECT 135.070 130.580 135.240 130.750 ;
        RECT 135.480 130.580 135.650 130.750 ;
        RECT 135.910 130.580 136.080 130.750 ;
        RECT 136.350 130.580 136.520 130.750 ;
        RECT 136.760 130.580 136.930 130.750 ;
        RECT 138.470 130.580 138.640 130.750 ;
        RECT 138.910 130.580 139.080 130.750 ;
        RECT 139.320 130.580 139.490 130.750 ;
        RECT 139.750 130.580 139.920 130.750 ;
        RECT 140.190 130.580 140.360 130.750 ;
        RECT 140.600 130.580 140.770 130.750 ;
        RECT 5.920 130.150 6.090 130.330 ;
        RECT 6.400 130.150 6.570 130.330 ;
        RECT 6.880 130.150 7.050 130.330 ;
        RECT 7.360 130.150 7.530 130.330 ;
        RECT 7.840 130.150 8.010 130.330 ;
        RECT 8.320 130.150 8.490 130.330 ;
        RECT 8.800 130.150 8.970 130.330 ;
        RECT 9.280 130.150 9.450 130.330 ;
        RECT 9.760 130.150 9.930 130.330 ;
        RECT 10.240 130.150 10.410 130.330 ;
        RECT 10.720 130.150 10.890 130.330 ;
        RECT 11.200 130.150 11.370 130.330 ;
        RECT 11.680 130.150 11.850 130.330 ;
        RECT 12.160 130.150 12.330 130.330 ;
        RECT 12.640 130.150 12.810 130.330 ;
        RECT 13.120 130.150 13.290 130.330 ;
        RECT 13.600 130.150 13.770 130.330 ;
        RECT 14.080 130.150 14.250 130.330 ;
        RECT 14.560 130.150 14.730 130.330 ;
        RECT 15.040 130.150 15.210 130.330 ;
        RECT 15.520 130.150 15.690 130.330 ;
        RECT 16.000 130.150 16.170 130.330 ;
        RECT 16.480 130.150 16.650 130.330 ;
        RECT 16.960 130.150 17.130 130.330 ;
        RECT 17.440 130.150 17.610 130.330 ;
        RECT 17.920 130.150 18.090 130.330 ;
        RECT 18.400 130.150 18.570 130.330 ;
        RECT 18.880 130.150 19.050 130.330 ;
        RECT 19.360 130.150 19.530 130.330 ;
        RECT 19.840 130.150 20.010 130.330 ;
        RECT 20.320 130.150 20.490 130.330 ;
        RECT 20.800 130.150 20.970 130.330 ;
        RECT 21.280 130.150 21.450 130.330 ;
        RECT 21.760 130.150 21.930 130.330 ;
        RECT 22.240 130.150 22.410 130.330 ;
        RECT 22.720 130.150 22.890 130.330 ;
        RECT 23.200 130.150 23.370 130.330 ;
        RECT 23.680 130.150 23.850 130.330 ;
        RECT 24.160 130.150 24.330 130.330 ;
        RECT 24.640 130.150 24.810 130.330 ;
        RECT 25.120 130.150 25.290 130.330 ;
        RECT 25.600 130.150 25.770 130.330 ;
        RECT 26.080 130.150 26.250 130.330 ;
        RECT 26.560 130.150 26.730 130.330 ;
        RECT 27.040 130.150 27.210 130.330 ;
        RECT 27.520 130.150 27.690 130.330 ;
        RECT 28.000 130.150 28.170 130.330 ;
        RECT 28.480 130.150 28.650 130.330 ;
        RECT 28.960 130.150 29.130 130.330 ;
        RECT 29.440 130.150 29.610 130.330 ;
        RECT 29.920 130.150 30.090 130.330 ;
        RECT 30.400 130.150 30.570 130.330 ;
        RECT 30.880 130.150 31.050 130.330 ;
        RECT 31.360 130.320 31.530 130.330 ;
      LAYER li1 ;
        RECT 31.200 130.150 31.680 130.320 ;
      LAYER li1 ;
        RECT 31.840 130.150 32.010 130.330 ;
        RECT 32.320 130.150 32.490 130.330 ;
        RECT 32.800 130.150 32.970 130.330 ;
        RECT 33.280 130.150 33.450 130.330 ;
        RECT 33.760 130.150 33.930 130.330 ;
      LAYER li1 ;
        RECT 34.080 130.320 34.560 130.330 ;
      LAYER li1 ;
        RECT 34.240 130.150 34.410 130.320 ;
        RECT 34.720 130.150 34.890 130.330 ;
        RECT 35.200 130.150 35.370 130.330 ;
        RECT 35.680 130.150 35.850 130.330 ;
        RECT 36.160 130.150 36.330 130.330 ;
        RECT 36.640 130.150 36.810 130.330 ;
        RECT 37.120 130.150 37.290 130.330 ;
        RECT 37.600 130.150 37.770 130.330 ;
        RECT 38.080 130.150 38.250 130.330 ;
        RECT 38.560 130.150 38.730 130.330 ;
        RECT 39.040 130.150 39.210 130.330 ;
        RECT 39.520 130.150 39.690 130.330 ;
        RECT 40.000 130.150 40.170 130.330 ;
        RECT 40.480 130.150 40.650 130.330 ;
        RECT 40.960 130.150 41.130 130.330 ;
        RECT 41.440 130.150 41.610 130.330 ;
        RECT 41.920 130.150 42.090 130.330 ;
        RECT 42.400 130.150 42.570 130.330 ;
        RECT 42.880 130.150 43.050 130.330 ;
        RECT 43.360 130.150 43.530 130.330 ;
      LAYER li1 ;
        RECT 43.680 130.320 44.160 130.330 ;
      LAYER li1 ;
        RECT 43.840 130.150 44.010 130.320 ;
        RECT 44.320 130.150 44.490 130.330 ;
        RECT 44.800 130.150 44.970 130.330 ;
        RECT 45.280 130.150 45.450 130.330 ;
        RECT 45.760 130.150 45.930 130.330 ;
        RECT 46.240 130.150 46.410 130.330 ;
        RECT 46.720 130.150 46.890 130.330 ;
        RECT 47.200 130.150 47.370 130.330 ;
        RECT 47.680 130.150 47.850 130.330 ;
        RECT 48.160 130.150 48.330 130.330 ;
        RECT 48.640 130.150 48.810 130.330 ;
        RECT 49.120 130.150 49.290 130.330 ;
        RECT 49.600 130.150 49.770 130.330 ;
        RECT 50.080 130.150 50.250 130.330 ;
        RECT 50.560 130.150 50.730 130.330 ;
        RECT 51.040 130.150 51.210 130.330 ;
        RECT 51.520 130.150 51.690 130.330 ;
        RECT 52.000 130.150 52.170 130.330 ;
        RECT 52.480 130.150 52.650 130.330 ;
        RECT 52.960 130.150 53.130 130.330 ;
        RECT 53.440 130.150 53.610 130.330 ;
        RECT 53.920 130.150 54.090 130.330 ;
        RECT 54.400 130.150 54.570 130.330 ;
        RECT 54.880 130.150 55.050 130.330 ;
        RECT 55.360 130.150 55.530 130.330 ;
        RECT 55.840 130.150 56.010 130.330 ;
        RECT 56.320 130.150 56.490 130.330 ;
        RECT 56.800 130.150 56.970 130.330 ;
        RECT 57.280 130.150 57.450 130.330 ;
        RECT 57.760 130.150 57.930 130.330 ;
        RECT 58.240 130.150 58.410 130.330 ;
        RECT 58.720 130.150 58.890 130.330 ;
        RECT 59.200 130.150 59.370 130.330 ;
        RECT 59.680 130.150 59.850 130.330 ;
        RECT 60.160 130.150 60.330 130.330 ;
        RECT 60.640 130.150 60.810 130.330 ;
        RECT 61.120 130.150 61.290 130.330 ;
        RECT 61.600 130.150 61.770 130.330 ;
        RECT 62.080 130.150 62.250 130.330 ;
        RECT 62.560 130.150 62.730 130.330 ;
        RECT 63.040 130.150 63.210 130.330 ;
        RECT 63.520 130.150 63.690 130.330 ;
        RECT 64.000 130.150 64.170 130.330 ;
        RECT 64.480 130.150 64.650 130.330 ;
        RECT 64.960 130.150 65.130 130.330 ;
        RECT 65.440 130.150 65.610 130.330 ;
        RECT 65.920 130.150 66.090 130.330 ;
        RECT 66.400 130.150 66.570 130.330 ;
        RECT 66.880 130.150 67.050 130.330 ;
        RECT 67.360 130.150 67.530 130.330 ;
        RECT 67.840 130.150 68.010 130.330 ;
        RECT 68.320 130.150 68.490 130.330 ;
        RECT 68.800 130.150 68.970 130.330 ;
        RECT 69.280 130.150 69.450 130.330 ;
        RECT 69.760 130.150 69.930 130.330 ;
        RECT 70.240 130.150 70.410 130.330 ;
        RECT 70.720 130.150 70.890 130.330 ;
        RECT 71.200 130.150 71.370 130.330 ;
        RECT 71.680 130.150 71.850 130.330 ;
        RECT 72.160 130.150 72.330 130.330 ;
        RECT 72.640 130.150 72.810 130.330 ;
        RECT 73.120 130.320 73.290 130.330 ;
      LAYER li1 ;
        RECT 72.960 130.150 73.440 130.320 ;
      LAYER li1 ;
        RECT 73.600 130.150 73.770 130.330 ;
      LAYER li1 ;
        RECT 73.920 130.320 74.400 130.330 ;
      LAYER li1 ;
        RECT 74.080 130.150 74.250 130.320 ;
        RECT 74.560 130.150 74.730 130.330 ;
        RECT 75.040 130.150 75.210 130.330 ;
        RECT 75.520 130.150 75.690 130.330 ;
        RECT 76.000 130.150 76.170 130.330 ;
        RECT 76.480 130.150 76.650 130.330 ;
        RECT 76.960 130.150 77.130 130.330 ;
        RECT 77.440 130.150 77.610 130.330 ;
        RECT 77.920 130.150 78.090 130.330 ;
        RECT 78.400 130.150 78.570 130.330 ;
        RECT 78.880 130.150 79.050 130.330 ;
        RECT 79.360 130.150 79.530 130.330 ;
        RECT 79.840 130.150 80.010 130.330 ;
        RECT 80.320 130.150 80.490 130.330 ;
        RECT 80.800 130.150 80.970 130.330 ;
        RECT 81.280 130.150 81.450 130.330 ;
        RECT 81.760 130.150 81.930 130.330 ;
        RECT 82.240 130.150 82.410 130.330 ;
        RECT 82.720 130.150 82.890 130.330 ;
        RECT 83.200 130.150 83.370 130.330 ;
        RECT 83.680 130.150 83.850 130.330 ;
        RECT 84.160 130.150 84.330 130.330 ;
        RECT 84.640 130.150 84.810 130.330 ;
        RECT 85.120 130.150 85.290 130.330 ;
        RECT 85.600 130.150 85.770 130.330 ;
        RECT 86.080 130.150 86.250 130.330 ;
        RECT 86.560 130.150 86.730 130.330 ;
        RECT 87.040 130.150 87.210 130.330 ;
        RECT 87.520 130.150 87.690 130.330 ;
        RECT 88.000 130.150 88.170 130.330 ;
        RECT 88.480 130.150 88.650 130.330 ;
        RECT 88.960 130.150 89.130 130.330 ;
        RECT 89.440 130.150 89.610 130.330 ;
        RECT 89.920 130.150 90.090 130.330 ;
        RECT 90.400 130.150 90.570 130.330 ;
        RECT 90.880 130.150 91.050 130.330 ;
        RECT 91.360 130.150 91.530 130.330 ;
        RECT 91.840 130.150 92.010 130.330 ;
        RECT 92.320 130.150 92.490 130.330 ;
        RECT 92.800 130.150 92.970 130.330 ;
        RECT 93.280 130.150 93.450 130.330 ;
        RECT 93.760 130.150 93.930 130.330 ;
        RECT 94.240 130.150 94.410 130.330 ;
        RECT 94.720 130.150 94.890 130.330 ;
        RECT 95.200 130.150 95.370 130.330 ;
        RECT 95.680 130.150 95.850 130.330 ;
        RECT 96.160 130.150 96.330 130.330 ;
        RECT 96.640 130.150 96.810 130.330 ;
        RECT 97.120 130.150 97.290 130.330 ;
        RECT 97.600 130.150 97.770 130.330 ;
        RECT 98.080 130.150 98.250 130.330 ;
        RECT 98.560 130.150 98.730 130.330 ;
        RECT 99.040 130.150 99.210 130.330 ;
        RECT 99.520 130.150 99.690 130.330 ;
        RECT 100.000 130.150 100.170 130.330 ;
        RECT 100.480 130.150 100.650 130.330 ;
        RECT 100.960 130.150 101.130 130.330 ;
        RECT 101.440 130.150 101.610 130.330 ;
        RECT 101.920 130.150 102.090 130.330 ;
        RECT 102.400 130.150 102.570 130.330 ;
        RECT 102.880 130.150 103.050 130.330 ;
        RECT 103.360 130.150 103.530 130.330 ;
        RECT 103.840 130.150 104.010 130.330 ;
        RECT 104.320 130.150 104.490 130.330 ;
        RECT 104.800 130.150 104.970 130.330 ;
        RECT 105.280 130.150 105.450 130.330 ;
        RECT 105.760 130.150 105.930 130.330 ;
        RECT 106.240 130.150 106.410 130.330 ;
        RECT 106.720 130.150 106.890 130.330 ;
        RECT 107.200 130.150 107.370 130.330 ;
        RECT 107.680 130.150 107.850 130.330 ;
        RECT 108.160 130.150 108.330 130.330 ;
        RECT 108.640 130.150 108.810 130.330 ;
        RECT 109.120 130.150 109.290 130.330 ;
        RECT 109.600 130.150 109.770 130.330 ;
        RECT 110.080 130.150 110.250 130.330 ;
      LAYER li1 ;
        RECT 110.400 130.150 110.880 130.330 ;
      LAYER li1 ;
        RECT 111.040 130.150 111.210 130.330 ;
        RECT 111.520 130.150 111.690 130.330 ;
        RECT 112.000 130.150 112.170 130.330 ;
        RECT 112.480 130.150 112.650 130.330 ;
        RECT 112.960 130.150 113.130 130.330 ;
        RECT 113.440 130.150 113.610 130.330 ;
        RECT 113.920 130.150 114.090 130.330 ;
        RECT 114.400 130.150 114.570 130.330 ;
        RECT 114.880 130.150 115.050 130.330 ;
        RECT 115.360 130.150 115.530 130.330 ;
        RECT 115.840 130.150 116.010 130.330 ;
        RECT 116.320 130.150 116.490 130.330 ;
        RECT 116.800 130.150 116.970 130.330 ;
        RECT 117.280 130.150 117.450 130.330 ;
        RECT 117.760 130.150 117.930 130.330 ;
      LAYER li1 ;
        RECT 118.080 130.320 118.560 130.330 ;
      LAYER li1 ;
        RECT 118.240 130.150 118.410 130.320 ;
        RECT 118.720 130.150 118.890 130.330 ;
        RECT 119.200 130.150 119.370 130.330 ;
        RECT 119.680 130.150 119.850 130.330 ;
        RECT 120.160 130.150 120.330 130.330 ;
        RECT 120.640 130.150 120.810 130.330 ;
        RECT 121.120 130.150 121.290 130.330 ;
        RECT 121.600 130.150 121.770 130.330 ;
        RECT 122.080 130.150 122.250 130.330 ;
        RECT 122.560 130.150 122.730 130.330 ;
        RECT 123.040 130.150 123.210 130.330 ;
        RECT 123.520 130.150 123.690 130.330 ;
        RECT 124.000 130.150 124.170 130.330 ;
        RECT 124.480 130.150 124.650 130.330 ;
        RECT 124.960 130.150 125.130 130.330 ;
        RECT 125.440 130.150 125.610 130.330 ;
        RECT 125.920 130.150 126.090 130.330 ;
        RECT 126.400 130.150 126.570 130.330 ;
        RECT 126.880 130.150 127.050 130.330 ;
        RECT 127.360 130.150 127.530 130.330 ;
        RECT 127.840 130.150 128.010 130.330 ;
        RECT 128.320 130.150 128.490 130.330 ;
        RECT 128.800 130.150 128.970 130.330 ;
        RECT 129.280 130.150 129.450 130.330 ;
        RECT 129.760 130.150 129.930 130.330 ;
        RECT 130.240 130.150 130.410 130.330 ;
        RECT 130.720 130.150 130.890 130.330 ;
        RECT 131.200 130.150 131.370 130.330 ;
        RECT 131.680 130.150 131.850 130.330 ;
        RECT 132.160 130.150 132.330 130.330 ;
        RECT 132.640 130.150 132.810 130.330 ;
        RECT 133.120 130.150 133.290 130.330 ;
        RECT 133.600 130.150 133.770 130.330 ;
        RECT 134.080 130.150 134.250 130.330 ;
        RECT 134.560 130.150 134.730 130.330 ;
        RECT 135.040 130.150 135.210 130.330 ;
        RECT 135.520 130.150 135.690 130.330 ;
        RECT 136.000 130.150 136.170 130.330 ;
        RECT 136.480 130.150 136.650 130.330 ;
        RECT 136.960 130.150 137.130 130.330 ;
        RECT 137.440 130.150 137.610 130.330 ;
        RECT 137.920 130.150 138.090 130.330 ;
        RECT 138.400 130.150 138.570 130.330 ;
        RECT 138.880 130.150 139.050 130.330 ;
        RECT 139.360 130.150 139.530 130.330 ;
        RECT 139.840 130.150 140.010 130.330 ;
        RECT 140.320 130.150 140.490 130.330 ;
        RECT 140.800 130.150 140.970 130.330 ;
        RECT 141.280 130.150 141.450 130.330 ;
        RECT 141.760 130.320 141.930 130.330 ;
      LAYER li1 ;
        RECT 141.600 130.150 142.080 130.320 ;
      LAYER li1 ;
        RECT 6.470 129.730 6.640 129.900 ;
        RECT 6.910 129.730 7.080 129.900 ;
        RECT 7.320 129.730 7.490 129.900 ;
        RECT 7.750 129.730 7.920 129.900 ;
        RECT 8.190 129.730 8.360 129.900 ;
        RECT 8.600 129.730 8.770 129.900 ;
        RECT 10.310 129.730 10.480 129.900 ;
        RECT 10.750 129.730 10.920 129.900 ;
        RECT 11.160 129.730 11.330 129.900 ;
        RECT 11.590 129.730 11.760 129.900 ;
        RECT 12.030 129.730 12.200 129.900 ;
        RECT 12.440 129.730 12.610 129.900 ;
        RECT 13.940 129.730 14.110 129.900 ;
        RECT 14.300 129.730 14.470 129.900 ;
        RECT 14.740 129.730 14.910 129.900 ;
        RECT 16.100 129.680 16.270 129.850 ;
        RECT 16.460 129.680 16.630 129.850 ;
        RECT 18.470 129.730 18.640 129.900 ;
        RECT 18.910 129.730 19.080 129.900 ;
        RECT 19.320 129.730 19.490 129.900 ;
        RECT 19.750 129.730 19.920 129.900 ;
        RECT 20.190 129.730 20.360 129.900 ;
        RECT 20.600 129.730 20.770 129.900 ;
        RECT 22.310 129.730 22.480 129.900 ;
        RECT 22.750 129.730 22.920 129.900 ;
        RECT 23.160 129.730 23.330 129.900 ;
        RECT 23.590 129.730 23.760 129.900 ;
        RECT 24.030 129.730 24.200 129.900 ;
        RECT 24.440 129.730 24.610 129.900 ;
        RECT 26.150 129.730 26.320 129.900 ;
        RECT 26.590 129.730 26.760 129.900 ;
        RECT 27.000 129.730 27.170 129.900 ;
        RECT 27.430 129.730 27.600 129.900 ;
        RECT 27.870 129.730 28.040 129.900 ;
        RECT 28.280 129.730 28.450 129.900 ;
        RECT 29.990 129.730 30.160 129.900 ;
        RECT 30.430 129.730 30.600 129.900 ;
        RECT 30.840 129.730 31.010 129.900 ;
        RECT 31.270 129.730 31.440 129.900 ;
        RECT 31.710 129.730 31.880 129.900 ;
        RECT 32.120 129.730 32.290 129.900 ;
        RECT 35.130 129.680 35.300 129.850 ;
        RECT 35.490 129.680 35.660 129.850 ;
        RECT 35.850 129.680 36.020 129.850 ;
        RECT 38.300 129.680 38.470 129.850 ;
        RECT 38.660 129.680 38.830 129.850 ;
        RECT 39.020 129.680 39.190 129.850 ;
        RECT 40.550 129.730 40.720 129.900 ;
        RECT 40.990 129.730 41.160 129.900 ;
        RECT 41.400 129.730 41.570 129.900 ;
        RECT 41.830 129.730 42.000 129.900 ;
        RECT 42.270 129.730 42.440 129.900 ;
        RECT 42.680 129.730 42.850 129.900 ;
        RECT 44.260 129.680 44.430 129.850 ;
        RECT 44.620 129.680 44.790 129.850 ;
        RECT 44.980 129.680 45.150 129.850 ;
        RECT 45.340 129.680 45.510 129.850 ;
        RECT 46.500 129.680 46.670 129.850 ;
        RECT 46.860 129.680 47.030 129.850 ;
        RECT 47.220 129.680 47.390 129.850 ;
        RECT 47.580 129.680 47.750 129.850 ;
        RECT 48.500 129.730 48.670 129.900 ;
        RECT 48.860 129.730 49.030 129.900 ;
        RECT 49.300 129.730 49.470 129.900 ;
        RECT 50.500 129.680 50.670 129.850 ;
        RECT 50.860 129.680 51.030 129.850 ;
        RECT 51.220 129.680 51.390 129.850 ;
        RECT 52.190 129.680 52.360 129.850 ;
        RECT 55.560 129.680 55.730 129.850 ;
        RECT 57.030 129.680 57.200 129.850 ;
        RECT 57.390 129.680 57.560 129.850 ;
        RECT 57.750 129.680 57.920 129.850 ;
        RECT 59.960 129.680 60.130 129.850 ;
        RECT 60.320 129.680 60.490 129.850 ;
        RECT 60.680 129.680 60.850 129.850 ;
        RECT 61.680 129.680 61.850 129.850 ;
        RECT 62.040 129.680 62.210 129.850 ;
        RECT 62.400 129.680 62.570 129.850 ;
        RECT 63.240 129.680 63.410 129.850 ;
        RECT 63.600 129.680 63.770 129.850 ;
        RECT 63.960 129.680 64.130 129.850 ;
        RECT 65.300 129.730 65.470 129.900 ;
        RECT 65.660 129.730 65.830 129.900 ;
        RECT 66.100 129.730 66.270 129.900 ;
        RECT 67.800 129.680 67.970 129.850 ;
        RECT 68.160 129.680 68.330 129.850 ;
        RECT 69.830 129.730 70.000 129.900 ;
        RECT 70.270 129.730 70.440 129.900 ;
        RECT 70.680 129.730 70.850 129.900 ;
        RECT 71.110 129.730 71.280 129.900 ;
        RECT 71.550 129.730 71.720 129.900 ;
        RECT 71.960 129.730 72.130 129.900 ;
        RECT 74.950 129.680 75.120 129.850 ;
        RECT 75.310 129.680 75.480 129.850 ;
        RECT 75.670 129.680 75.840 129.850 ;
        RECT 77.260 129.680 77.430 129.850 ;
        RECT 77.620 129.680 77.790 129.850 ;
        RECT 77.980 129.680 78.150 129.850 ;
        RECT 79.220 129.730 79.390 129.900 ;
        RECT 79.580 129.730 79.750 129.900 ;
        RECT 80.020 129.730 80.190 129.900 ;
        RECT 80.760 129.680 80.930 129.850 ;
        RECT 81.120 129.680 81.290 129.850 ;
        RECT 81.480 129.680 81.650 129.850 ;
        RECT 81.840 129.680 82.010 129.850 ;
        RECT 82.200 129.680 82.370 129.850 ;
        RECT 84.710 129.730 84.880 129.900 ;
        RECT 85.150 129.730 85.320 129.900 ;
        RECT 85.560 129.730 85.730 129.900 ;
        RECT 85.990 129.730 86.160 129.900 ;
        RECT 86.430 129.730 86.600 129.900 ;
        RECT 86.840 129.730 87.010 129.900 ;
        RECT 88.550 129.730 88.720 129.900 ;
        RECT 88.990 129.730 89.160 129.900 ;
        RECT 89.400 129.730 89.570 129.900 ;
        RECT 89.830 129.730 90.000 129.900 ;
        RECT 90.270 129.730 90.440 129.900 ;
        RECT 90.680 129.730 90.850 129.900 ;
        RECT 92.390 129.730 92.560 129.900 ;
        RECT 92.830 129.730 93.000 129.900 ;
        RECT 93.240 129.730 93.410 129.900 ;
        RECT 93.670 129.730 93.840 129.900 ;
        RECT 94.110 129.730 94.280 129.900 ;
        RECT 94.520 129.730 94.690 129.900 ;
        RECT 96.020 129.730 96.190 129.900 ;
        RECT 96.380 129.730 96.550 129.900 ;
        RECT 96.820 129.730 96.990 129.900 ;
        RECT 98.000 129.680 98.170 129.850 ;
        RECT 98.360 129.680 98.530 129.850 ;
        RECT 98.720 129.680 98.890 129.850 ;
        RECT 99.080 129.680 99.250 129.850 ;
        RECT 99.440 129.680 99.610 129.850 ;
        RECT 99.800 129.680 99.970 129.850 ;
        RECT 100.160 129.680 100.330 129.850 ;
        RECT 100.520 129.680 100.690 129.850 ;
        RECT 101.330 129.680 101.500 129.850 ;
        RECT 101.690 129.680 101.860 129.850 ;
        RECT 102.050 129.680 102.220 129.850 ;
        RECT 102.410 129.680 102.580 129.850 ;
        RECT 103.430 129.730 103.600 129.900 ;
        RECT 103.870 129.730 104.040 129.900 ;
        RECT 104.280 129.730 104.450 129.900 ;
        RECT 104.710 129.730 104.880 129.900 ;
        RECT 105.150 129.730 105.320 129.900 ;
        RECT 105.560 129.730 105.730 129.900 ;
        RECT 107.270 129.730 107.440 129.900 ;
        RECT 107.710 129.730 107.880 129.900 ;
        RECT 108.120 129.730 108.290 129.900 ;
        RECT 108.550 129.730 108.720 129.900 ;
        RECT 108.990 129.730 109.160 129.900 ;
        RECT 109.400 129.730 109.570 129.900 ;
        RECT 111.620 129.680 111.790 129.850 ;
        RECT 111.980 129.680 112.150 129.850 ;
        RECT 113.990 129.730 114.160 129.900 ;
        RECT 114.430 129.730 114.600 129.900 ;
        RECT 114.840 129.730 115.010 129.900 ;
        RECT 115.270 129.730 115.440 129.900 ;
        RECT 115.710 129.730 115.880 129.900 ;
        RECT 116.120 129.730 116.290 129.900 ;
        RECT 119.300 129.680 119.470 129.850 ;
        RECT 119.660 129.680 119.830 129.850 ;
        RECT 121.670 129.730 121.840 129.900 ;
        RECT 122.110 129.730 122.280 129.900 ;
        RECT 122.520 129.730 122.690 129.900 ;
        RECT 122.950 129.730 123.120 129.900 ;
        RECT 123.390 129.730 123.560 129.900 ;
        RECT 123.800 129.730 123.970 129.900 ;
        RECT 125.510 129.730 125.680 129.900 ;
        RECT 125.950 129.730 126.120 129.900 ;
        RECT 126.360 129.730 126.530 129.900 ;
        RECT 126.790 129.730 126.960 129.900 ;
        RECT 127.230 129.730 127.400 129.900 ;
        RECT 127.640 129.730 127.810 129.900 ;
        RECT 129.350 129.730 129.520 129.900 ;
        RECT 129.790 129.730 129.960 129.900 ;
        RECT 130.200 129.730 130.370 129.900 ;
        RECT 130.630 129.730 130.800 129.900 ;
        RECT 131.070 129.730 131.240 129.900 ;
        RECT 131.480 129.730 131.650 129.900 ;
        RECT 133.190 129.730 133.360 129.900 ;
        RECT 133.630 129.730 133.800 129.900 ;
        RECT 134.040 129.730 134.210 129.900 ;
        RECT 134.470 129.730 134.640 129.900 ;
        RECT 134.910 129.730 135.080 129.900 ;
        RECT 135.320 129.730 135.490 129.900 ;
        RECT 137.030 129.730 137.200 129.900 ;
        RECT 137.470 129.730 137.640 129.900 ;
        RECT 137.880 129.730 138.050 129.900 ;
        RECT 138.310 129.730 138.480 129.900 ;
        RECT 138.750 129.730 138.920 129.900 ;
        RECT 139.160 129.730 139.330 129.900 ;
        RECT 140.660 129.730 140.830 129.900 ;
        RECT 141.020 129.730 141.190 129.900 ;
        RECT 141.460 129.730 141.630 129.900 ;
        RECT 6.260 122.440 6.430 122.610 ;
        RECT 6.620 122.440 6.790 122.610 ;
        RECT 7.060 122.440 7.230 122.610 ;
        RECT 8.820 122.490 8.990 122.660 ;
        RECT 9.180 122.490 9.350 122.660 ;
        RECT 11.210 122.490 11.380 122.660 ;
        RECT 13.640 122.490 13.810 122.660 ;
        RECT 14.000 122.490 14.170 122.660 ;
        RECT 14.360 122.490 14.530 122.660 ;
        RECT 15.980 122.490 16.150 122.660 ;
        RECT 16.340 122.490 16.510 122.660 ;
        RECT 16.700 122.490 16.870 122.660 ;
        RECT 18.680 122.490 18.850 122.660 ;
        RECT 19.040 122.490 19.210 122.660 ;
        RECT 19.400 122.490 19.570 122.660 ;
        RECT 20.430 122.490 20.600 122.660 ;
        RECT 20.790 122.490 20.960 122.660 ;
        RECT 21.150 122.490 21.320 122.660 ;
        RECT 21.960 122.490 22.130 122.660 ;
        RECT 22.320 122.490 22.490 122.660 ;
        RECT 22.680 122.490 22.850 122.660 ;
        RECT 24.020 122.440 24.190 122.610 ;
        RECT 24.380 122.440 24.550 122.610 ;
        RECT 24.820 122.440 24.990 122.610 ;
        RECT 27.060 122.490 27.230 122.660 ;
        RECT 27.420 122.490 27.590 122.660 ;
        RECT 29.450 122.490 29.620 122.660 ;
        RECT 31.880 122.490 32.050 122.660 ;
        RECT 32.240 122.490 32.410 122.660 ;
        RECT 32.600 122.490 32.770 122.660 ;
        RECT 34.220 122.490 34.390 122.660 ;
        RECT 34.580 122.490 34.750 122.660 ;
        RECT 34.940 122.490 35.110 122.660 ;
        RECT 36.920 122.490 37.090 122.660 ;
        RECT 37.280 122.490 37.450 122.660 ;
        RECT 37.640 122.490 37.810 122.660 ;
        RECT 38.670 122.490 38.840 122.660 ;
        RECT 39.030 122.490 39.200 122.660 ;
        RECT 39.390 122.490 39.560 122.660 ;
        RECT 40.200 122.490 40.370 122.660 ;
        RECT 40.560 122.490 40.730 122.660 ;
        RECT 40.920 122.490 41.090 122.660 ;
        RECT 42.260 122.440 42.430 122.610 ;
        RECT 42.620 122.440 42.790 122.610 ;
        RECT 43.060 122.440 43.230 122.610 ;
        RECT 44.730 122.490 44.900 122.660 ;
        RECT 45.090 122.490 45.260 122.660 ;
        RECT 45.450 122.490 45.620 122.660 ;
        RECT 47.900 122.490 48.070 122.660 ;
        RECT 48.260 122.490 48.430 122.660 ;
        RECT 48.620 122.490 48.790 122.660 ;
        RECT 50.150 122.440 50.320 122.610 ;
        RECT 50.590 122.440 50.760 122.610 ;
        RECT 51.000 122.440 51.170 122.610 ;
        RECT 51.430 122.440 51.600 122.610 ;
        RECT 51.870 122.440 52.040 122.610 ;
        RECT 52.280 122.440 52.450 122.610 ;
        RECT 53.990 122.440 54.160 122.610 ;
        RECT 54.430 122.440 54.600 122.610 ;
        RECT 54.840 122.440 55.010 122.610 ;
        RECT 55.270 122.440 55.440 122.610 ;
        RECT 55.710 122.440 55.880 122.610 ;
        RECT 56.120 122.440 56.290 122.610 ;
        RECT 58.820 122.490 58.990 122.660 ;
        RECT 59.180 122.490 59.350 122.660 ;
        RECT 61.190 122.440 61.360 122.610 ;
        RECT 61.630 122.440 61.800 122.610 ;
        RECT 62.040 122.440 62.210 122.610 ;
        RECT 62.470 122.440 62.640 122.610 ;
        RECT 62.910 122.440 63.080 122.610 ;
        RECT 63.320 122.440 63.490 122.610 ;
        RECT 65.030 122.440 65.200 122.610 ;
        RECT 65.470 122.440 65.640 122.610 ;
        RECT 65.880 122.440 66.050 122.610 ;
        RECT 66.310 122.440 66.480 122.610 ;
        RECT 66.750 122.440 66.920 122.610 ;
        RECT 67.160 122.440 67.330 122.610 ;
        RECT 68.870 122.440 69.040 122.610 ;
        RECT 69.310 122.440 69.480 122.610 ;
        RECT 69.720 122.440 69.890 122.610 ;
        RECT 70.150 122.440 70.320 122.610 ;
        RECT 70.590 122.440 70.760 122.610 ;
        RECT 71.000 122.440 71.170 122.610 ;
        RECT 72.500 122.440 72.670 122.610 ;
        RECT 72.860 122.440 73.030 122.610 ;
        RECT 73.300 122.440 73.470 122.610 ;
        RECT 75.000 122.490 75.170 122.660 ;
        RECT 75.360 122.490 75.530 122.660 ;
        RECT 75.720 122.490 75.890 122.660 ;
        RECT 76.080 122.490 76.250 122.660 ;
        RECT 76.440 122.490 76.610 122.660 ;
        RECT 78.950 122.440 79.120 122.610 ;
        RECT 79.390 122.440 79.560 122.610 ;
        RECT 79.800 122.440 79.970 122.610 ;
        RECT 80.230 122.440 80.400 122.610 ;
        RECT 80.670 122.440 80.840 122.610 ;
        RECT 81.080 122.440 81.250 122.610 ;
        RECT 82.790 122.440 82.960 122.610 ;
        RECT 83.230 122.440 83.400 122.610 ;
        RECT 83.640 122.440 83.810 122.610 ;
        RECT 84.070 122.440 84.240 122.610 ;
        RECT 84.510 122.440 84.680 122.610 ;
        RECT 84.920 122.440 85.090 122.610 ;
        RECT 86.630 122.440 86.800 122.610 ;
        RECT 87.070 122.440 87.240 122.610 ;
        RECT 87.480 122.440 87.650 122.610 ;
        RECT 87.910 122.440 88.080 122.610 ;
        RECT 88.350 122.440 88.520 122.610 ;
        RECT 88.760 122.440 88.930 122.610 ;
        RECT 90.840 122.490 91.010 122.660 ;
        RECT 91.200 122.490 91.370 122.660 ;
        RECT 92.660 122.440 92.830 122.610 ;
        RECT 93.020 122.440 93.190 122.610 ;
        RECT 93.460 122.440 93.630 122.610 ;
        RECT 94.640 122.490 94.810 122.660 ;
        RECT 95.000 122.490 95.170 122.660 ;
        RECT 95.360 122.490 95.530 122.660 ;
        RECT 95.720 122.490 95.890 122.660 ;
        RECT 96.080 122.490 96.250 122.660 ;
        RECT 96.440 122.490 96.610 122.660 ;
        RECT 96.800 122.490 96.970 122.660 ;
        RECT 97.160 122.490 97.330 122.660 ;
        RECT 97.970 122.490 98.140 122.660 ;
        RECT 98.330 122.490 98.500 122.660 ;
        RECT 98.690 122.490 98.860 122.660 ;
        RECT 99.050 122.490 99.220 122.660 ;
        RECT 99.860 122.440 100.030 122.610 ;
        RECT 100.220 122.440 100.390 122.610 ;
        RECT 100.660 122.440 100.830 122.610 ;
        RECT 101.380 122.490 101.550 122.660 ;
        RECT 101.740 122.490 101.910 122.660 ;
        RECT 102.100 122.490 102.270 122.660 ;
        RECT 102.460 122.490 102.630 122.660 ;
        RECT 103.620 122.490 103.790 122.660 ;
        RECT 103.980 122.490 104.150 122.660 ;
        RECT 104.340 122.490 104.510 122.660 ;
        RECT 104.700 122.490 104.870 122.660 ;
        RECT 105.620 122.440 105.790 122.610 ;
        RECT 105.980 122.440 106.150 122.610 ;
        RECT 106.420 122.440 106.590 122.610 ;
        RECT 107.160 122.490 107.330 122.660 ;
        RECT 107.520 122.490 107.690 122.660 ;
        RECT 108.980 122.440 109.150 122.610 ;
        RECT 109.340 122.440 109.510 122.610 ;
        RECT 109.780 122.440 109.950 122.610 ;
        RECT 112.020 122.490 112.190 122.660 ;
        RECT 112.380 122.490 112.550 122.660 ;
        RECT 114.410 122.490 114.580 122.660 ;
        RECT 116.840 122.490 117.010 122.660 ;
        RECT 117.200 122.490 117.370 122.660 ;
        RECT 117.560 122.490 117.730 122.660 ;
        RECT 119.180 122.490 119.350 122.660 ;
        RECT 119.540 122.490 119.710 122.660 ;
        RECT 119.900 122.490 120.070 122.660 ;
        RECT 121.880 122.490 122.050 122.660 ;
        RECT 122.240 122.490 122.410 122.660 ;
        RECT 122.600 122.490 122.770 122.660 ;
        RECT 123.630 122.490 123.800 122.660 ;
        RECT 123.990 122.490 124.160 122.660 ;
        RECT 124.350 122.490 124.520 122.660 ;
        RECT 125.160 122.490 125.330 122.660 ;
        RECT 125.520 122.490 125.690 122.660 ;
        RECT 125.880 122.490 126.050 122.660 ;
        RECT 127.430 122.440 127.600 122.610 ;
        RECT 127.870 122.440 128.040 122.610 ;
        RECT 128.280 122.440 128.450 122.610 ;
        RECT 128.710 122.440 128.880 122.610 ;
        RECT 129.150 122.440 129.320 122.610 ;
        RECT 129.560 122.440 129.730 122.610 ;
        RECT 131.270 122.440 131.440 122.610 ;
        RECT 131.710 122.440 131.880 122.610 ;
        RECT 132.120 122.440 132.290 122.610 ;
        RECT 132.550 122.440 132.720 122.610 ;
        RECT 132.990 122.440 133.160 122.610 ;
        RECT 133.400 122.440 133.570 122.610 ;
        RECT 135.110 122.440 135.280 122.610 ;
        RECT 135.550 122.440 135.720 122.610 ;
        RECT 135.960 122.440 136.130 122.610 ;
        RECT 136.390 122.440 136.560 122.610 ;
        RECT 136.830 122.440 137.000 122.610 ;
        RECT 137.240 122.440 137.410 122.610 ;
        RECT 138.950 122.440 139.120 122.610 ;
        RECT 139.390 122.440 139.560 122.610 ;
        RECT 139.800 122.440 139.970 122.610 ;
        RECT 140.230 122.440 140.400 122.610 ;
        RECT 140.670 122.440 140.840 122.610 ;
        RECT 141.080 122.440 141.250 122.610 ;
        RECT 5.920 122.010 6.090 122.190 ;
        RECT 6.400 122.010 6.570 122.190 ;
        RECT 6.880 122.010 7.050 122.190 ;
        RECT 7.360 122.010 7.530 122.190 ;
        RECT 7.840 122.020 8.010 122.190 ;
      LAYER li1 ;
        RECT 7.680 122.010 8.160 122.020 ;
      LAYER li1 ;
        RECT 8.320 122.010 8.490 122.190 ;
        RECT 8.800 122.010 8.970 122.190 ;
        RECT 9.280 122.010 9.450 122.190 ;
        RECT 9.760 122.010 9.930 122.190 ;
        RECT 10.240 122.010 10.410 122.190 ;
      LAYER li1 ;
        RECT 10.560 122.180 11.040 122.190 ;
      LAYER li1 ;
        RECT 10.720 122.010 10.890 122.180 ;
        RECT 11.200 122.010 11.370 122.190 ;
        RECT 11.680 122.010 11.850 122.190 ;
        RECT 12.160 122.010 12.330 122.190 ;
        RECT 12.640 122.010 12.810 122.190 ;
        RECT 13.120 122.010 13.290 122.190 ;
        RECT 13.600 122.010 13.770 122.190 ;
        RECT 14.080 122.010 14.250 122.190 ;
        RECT 14.560 122.010 14.730 122.190 ;
        RECT 15.040 122.010 15.210 122.190 ;
        RECT 15.520 122.010 15.690 122.190 ;
        RECT 16.000 122.010 16.170 122.190 ;
        RECT 16.480 122.010 16.650 122.190 ;
        RECT 16.960 122.010 17.130 122.190 ;
        RECT 17.440 122.010 17.610 122.190 ;
        RECT 17.920 122.010 18.090 122.190 ;
        RECT 18.400 122.010 18.570 122.190 ;
        RECT 18.880 122.010 19.050 122.190 ;
        RECT 19.360 122.010 19.530 122.190 ;
        RECT 19.840 122.010 20.010 122.190 ;
        RECT 20.320 122.010 20.490 122.190 ;
        RECT 20.800 122.010 20.970 122.190 ;
        RECT 21.280 122.010 21.450 122.190 ;
        RECT 21.760 122.010 21.930 122.190 ;
        RECT 22.240 122.010 22.410 122.190 ;
        RECT 22.720 122.010 22.890 122.190 ;
        RECT 23.200 122.010 23.370 122.190 ;
        RECT 23.680 122.010 23.850 122.190 ;
        RECT 24.160 122.010 24.330 122.190 ;
        RECT 24.640 122.010 24.810 122.190 ;
        RECT 25.120 122.010 25.290 122.190 ;
        RECT 25.600 122.010 25.770 122.190 ;
        RECT 26.080 122.010 26.250 122.190 ;
        RECT 26.560 122.010 26.730 122.190 ;
        RECT 27.040 122.010 27.210 122.190 ;
        RECT 27.520 122.010 27.690 122.190 ;
        RECT 28.000 122.010 28.170 122.190 ;
      LAYER li1 ;
        RECT 28.320 122.020 28.800 122.190 ;
      LAYER li1 ;
        RECT 28.480 122.010 28.650 122.020 ;
        RECT 28.960 122.010 29.130 122.190 ;
        RECT 29.440 122.010 29.610 122.190 ;
        RECT 29.920 122.010 30.090 122.190 ;
        RECT 30.400 122.010 30.570 122.190 ;
        RECT 30.880 122.010 31.050 122.190 ;
        RECT 31.360 122.010 31.530 122.190 ;
        RECT 31.840 122.010 32.010 122.190 ;
        RECT 32.320 122.010 32.490 122.190 ;
        RECT 32.800 122.010 32.970 122.190 ;
        RECT 33.280 122.010 33.450 122.190 ;
        RECT 33.760 122.010 33.930 122.190 ;
        RECT 34.240 122.010 34.410 122.190 ;
        RECT 34.720 122.010 34.890 122.190 ;
        RECT 35.200 122.010 35.370 122.190 ;
        RECT 35.680 122.010 35.850 122.190 ;
        RECT 36.160 122.010 36.330 122.190 ;
        RECT 36.640 122.010 36.810 122.190 ;
        RECT 37.120 122.010 37.290 122.190 ;
        RECT 37.600 122.010 37.770 122.190 ;
        RECT 38.080 122.010 38.250 122.190 ;
        RECT 38.560 122.010 38.730 122.190 ;
        RECT 39.040 122.010 39.210 122.190 ;
        RECT 39.520 122.010 39.690 122.190 ;
        RECT 40.000 122.010 40.170 122.190 ;
        RECT 40.480 122.010 40.650 122.190 ;
        RECT 40.960 122.010 41.130 122.190 ;
        RECT 41.440 122.010 41.610 122.190 ;
        RECT 41.920 122.010 42.090 122.190 ;
        RECT 42.400 122.010 42.570 122.190 ;
        RECT 42.880 122.010 43.050 122.190 ;
      LAYER li1 ;
        RECT 43.200 122.020 43.680 122.190 ;
      LAYER li1 ;
        RECT 43.840 122.020 44.010 122.190 ;
        RECT 43.360 122.010 43.530 122.020 ;
      LAYER li1 ;
        RECT 43.680 122.010 44.160 122.020 ;
      LAYER li1 ;
        RECT 44.320 122.010 44.490 122.190 ;
        RECT 44.800 122.010 44.970 122.190 ;
        RECT 45.280 122.010 45.450 122.190 ;
        RECT 45.760 122.010 45.930 122.190 ;
        RECT 46.240 122.010 46.410 122.190 ;
        RECT 46.720 122.010 46.890 122.190 ;
        RECT 47.200 122.010 47.370 122.190 ;
        RECT 47.680 122.010 47.850 122.190 ;
        RECT 48.160 122.010 48.330 122.190 ;
        RECT 48.640 122.010 48.810 122.190 ;
        RECT 49.120 122.010 49.290 122.190 ;
        RECT 49.600 122.010 49.770 122.190 ;
      LAYER li1 ;
        RECT 49.920 122.020 50.400 122.190 ;
      LAYER li1 ;
        RECT 50.080 122.010 50.250 122.020 ;
        RECT 50.560 122.010 50.730 122.190 ;
        RECT 51.040 122.010 51.210 122.190 ;
        RECT 51.520 122.010 51.690 122.190 ;
        RECT 52.000 122.010 52.170 122.190 ;
        RECT 52.480 122.010 52.650 122.190 ;
        RECT 52.960 122.010 53.130 122.190 ;
        RECT 53.440 122.010 53.610 122.190 ;
        RECT 53.920 122.010 54.090 122.190 ;
        RECT 54.400 122.010 54.570 122.190 ;
        RECT 54.880 122.010 55.050 122.190 ;
        RECT 55.360 122.010 55.530 122.190 ;
        RECT 55.840 122.010 56.010 122.190 ;
        RECT 56.320 122.010 56.490 122.190 ;
        RECT 56.800 122.010 56.970 122.190 ;
        RECT 57.280 122.010 57.450 122.190 ;
        RECT 57.760 122.010 57.930 122.190 ;
        RECT 58.240 122.010 58.410 122.190 ;
        RECT 58.720 122.010 58.890 122.190 ;
        RECT 59.200 122.010 59.370 122.190 ;
        RECT 59.680 122.010 59.850 122.190 ;
        RECT 60.160 122.010 60.330 122.190 ;
        RECT 60.640 122.010 60.810 122.190 ;
        RECT 61.120 122.010 61.290 122.190 ;
        RECT 61.600 122.010 61.770 122.190 ;
        RECT 62.080 122.010 62.250 122.190 ;
        RECT 62.560 122.010 62.730 122.190 ;
        RECT 63.040 122.010 63.210 122.190 ;
        RECT 63.520 122.010 63.690 122.190 ;
        RECT 64.000 122.010 64.170 122.190 ;
        RECT 64.480 122.010 64.650 122.190 ;
        RECT 64.960 122.010 65.130 122.190 ;
        RECT 65.440 122.010 65.610 122.190 ;
        RECT 65.920 122.010 66.090 122.190 ;
        RECT 66.400 122.010 66.570 122.190 ;
        RECT 66.880 122.010 67.050 122.190 ;
      LAYER li1 ;
        RECT 67.200 122.180 67.680 122.190 ;
      LAYER li1 ;
        RECT 67.360 122.010 67.530 122.180 ;
        RECT 67.840 122.010 68.010 122.190 ;
        RECT 68.320 122.010 68.490 122.190 ;
        RECT 68.800 122.010 68.970 122.190 ;
        RECT 69.280 122.010 69.450 122.190 ;
        RECT 69.760 122.010 69.930 122.190 ;
        RECT 70.240 122.010 70.410 122.190 ;
        RECT 70.720 122.010 70.890 122.190 ;
        RECT 71.200 122.010 71.370 122.190 ;
        RECT 71.680 122.010 71.850 122.190 ;
        RECT 72.160 122.010 72.330 122.190 ;
        RECT 72.640 122.010 72.810 122.190 ;
        RECT 73.120 122.010 73.290 122.190 ;
        RECT 73.600 122.010 73.770 122.190 ;
        RECT 74.080 122.010 74.250 122.190 ;
        RECT 74.560 122.010 74.730 122.190 ;
        RECT 75.040 122.010 75.210 122.190 ;
        RECT 75.520 122.010 75.690 122.190 ;
        RECT 76.000 122.010 76.170 122.190 ;
        RECT 76.480 122.010 76.650 122.190 ;
        RECT 76.960 122.010 77.130 122.190 ;
        RECT 77.440 122.010 77.610 122.190 ;
        RECT 77.920 122.010 78.090 122.190 ;
        RECT 78.400 122.010 78.570 122.190 ;
        RECT 78.880 122.010 79.050 122.190 ;
        RECT 79.360 122.010 79.530 122.190 ;
        RECT 79.840 122.010 80.010 122.190 ;
        RECT 80.320 122.010 80.490 122.190 ;
        RECT 80.800 122.010 80.970 122.190 ;
        RECT 81.280 122.010 81.450 122.190 ;
        RECT 81.760 122.010 81.930 122.190 ;
        RECT 82.240 122.010 82.410 122.190 ;
        RECT 82.720 122.010 82.890 122.190 ;
        RECT 83.200 122.010 83.370 122.190 ;
        RECT 83.680 122.010 83.850 122.190 ;
        RECT 84.160 122.010 84.330 122.190 ;
        RECT 84.640 122.010 84.810 122.190 ;
        RECT 85.120 122.010 85.290 122.190 ;
        RECT 85.600 122.010 85.770 122.190 ;
        RECT 86.080 122.010 86.250 122.190 ;
        RECT 86.560 122.010 86.730 122.190 ;
        RECT 87.040 122.010 87.210 122.190 ;
        RECT 87.520 122.010 87.690 122.190 ;
        RECT 88.000 122.010 88.170 122.190 ;
        RECT 88.480 122.010 88.650 122.190 ;
        RECT 88.960 122.010 89.130 122.190 ;
        RECT 89.440 122.010 89.610 122.190 ;
        RECT 89.920 122.010 90.090 122.190 ;
        RECT 90.400 122.010 90.570 122.190 ;
        RECT 90.880 122.010 91.050 122.190 ;
        RECT 91.360 122.010 91.530 122.190 ;
        RECT 91.840 122.010 92.010 122.190 ;
        RECT 92.320 122.010 92.490 122.190 ;
        RECT 92.800 122.010 92.970 122.190 ;
        RECT 93.280 122.010 93.450 122.190 ;
        RECT 93.760 122.010 93.930 122.190 ;
        RECT 94.240 122.010 94.410 122.190 ;
        RECT 94.720 122.010 94.890 122.190 ;
        RECT 95.200 122.010 95.370 122.190 ;
        RECT 95.680 122.010 95.850 122.190 ;
        RECT 96.160 122.010 96.330 122.190 ;
        RECT 96.640 122.010 96.810 122.190 ;
        RECT 97.120 122.010 97.290 122.190 ;
        RECT 97.600 122.010 97.770 122.190 ;
        RECT 98.080 122.010 98.250 122.190 ;
        RECT 98.560 122.010 98.730 122.190 ;
        RECT 99.040 122.010 99.210 122.190 ;
        RECT 99.520 122.010 99.690 122.190 ;
        RECT 100.000 122.010 100.170 122.190 ;
      LAYER li1 ;
        RECT 100.320 122.020 100.800 122.190 ;
      LAYER li1 ;
        RECT 100.480 122.010 100.650 122.020 ;
        RECT 100.960 122.010 101.130 122.190 ;
        RECT 101.440 122.010 101.610 122.190 ;
        RECT 101.920 122.010 102.090 122.190 ;
        RECT 102.400 122.010 102.570 122.190 ;
        RECT 102.880 122.010 103.050 122.190 ;
        RECT 103.360 122.010 103.530 122.190 ;
        RECT 103.840 122.010 104.010 122.190 ;
        RECT 104.320 122.010 104.490 122.190 ;
        RECT 104.800 122.010 104.970 122.190 ;
        RECT 105.280 122.010 105.450 122.190 ;
        RECT 105.760 122.010 105.930 122.190 ;
        RECT 106.240 122.010 106.410 122.190 ;
        RECT 106.720 122.010 106.890 122.190 ;
        RECT 107.200 122.010 107.370 122.190 ;
        RECT 107.680 122.010 107.850 122.190 ;
        RECT 108.160 122.010 108.330 122.190 ;
        RECT 108.640 122.010 108.810 122.190 ;
        RECT 109.120 122.010 109.290 122.190 ;
        RECT 109.600 122.010 109.770 122.190 ;
        RECT 110.080 122.010 110.250 122.190 ;
        RECT 110.560 122.010 110.730 122.190 ;
        RECT 111.040 122.010 111.210 122.190 ;
        RECT 111.520 122.010 111.690 122.190 ;
        RECT 112.000 122.010 112.170 122.190 ;
        RECT 112.480 122.010 112.650 122.190 ;
        RECT 112.960 122.010 113.130 122.190 ;
        RECT 113.440 122.010 113.610 122.190 ;
        RECT 113.920 122.010 114.090 122.190 ;
        RECT 114.400 122.010 114.570 122.190 ;
        RECT 114.880 122.010 115.050 122.190 ;
        RECT 115.360 122.010 115.530 122.190 ;
        RECT 115.840 122.010 116.010 122.190 ;
        RECT 116.320 122.010 116.490 122.190 ;
        RECT 116.800 122.010 116.970 122.190 ;
        RECT 117.280 122.010 117.450 122.190 ;
        RECT 117.760 122.010 117.930 122.190 ;
        RECT 118.240 122.010 118.410 122.190 ;
        RECT 118.720 122.010 118.890 122.190 ;
        RECT 119.200 122.010 119.370 122.190 ;
        RECT 119.680 122.010 119.850 122.190 ;
        RECT 120.160 122.010 120.330 122.190 ;
        RECT 120.640 122.010 120.810 122.190 ;
        RECT 121.120 122.010 121.290 122.190 ;
        RECT 121.600 122.010 121.770 122.190 ;
        RECT 122.080 122.010 122.250 122.190 ;
        RECT 122.560 122.010 122.730 122.190 ;
        RECT 123.040 122.010 123.210 122.190 ;
        RECT 123.520 122.010 123.690 122.190 ;
        RECT 124.000 122.010 124.170 122.190 ;
        RECT 124.480 122.010 124.650 122.190 ;
        RECT 124.960 122.010 125.130 122.190 ;
        RECT 125.440 122.010 125.610 122.190 ;
        RECT 125.920 122.010 126.090 122.190 ;
        RECT 126.400 122.010 126.570 122.190 ;
        RECT 126.880 122.010 127.050 122.190 ;
        RECT 127.360 122.010 127.530 122.190 ;
        RECT 127.840 122.010 128.010 122.190 ;
        RECT 128.320 122.010 128.490 122.190 ;
        RECT 128.800 122.010 128.970 122.190 ;
        RECT 129.280 122.010 129.450 122.190 ;
        RECT 129.760 122.010 129.930 122.190 ;
        RECT 130.240 122.010 130.410 122.190 ;
        RECT 130.720 122.010 130.890 122.190 ;
        RECT 131.200 122.010 131.370 122.190 ;
        RECT 131.680 122.010 131.850 122.190 ;
        RECT 132.160 122.010 132.330 122.190 ;
        RECT 132.640 122.010 132.810 122.190 ;
        RECT 133.120 122.010 133.290 122.190 ;
        RECT 133.600 122.010 133.770 122.190 ;
        RECT 134.080 122.010 134.250 122.190 ;
        RECT 134.560 122.010 134.730 122.190 ;
        RECT 135.040 122.010 135.210 122.190 ;
        RECT 135.520 122.010 135.690 122.190 ;
        RECT 136.000 122.010 136.170 122.190 ;
        RECT 136.480 122.010 136.650 122.190 ;
        RECT 136.960 122.010 137.130 122.190 ;
        RECT 137.440 122.010 137.610 122.190 ;
        RECT 137.920 122.010 138.090 122.190 ;
        RECT 138.400 122.010 138.570 122.190 ;
        RECT 138.880 122.010 139.050 122.190 ;
        RECT 139.360 122.010 139.530 122.190 ;
        RECT 139.840 122.010 140.010 122.190 ;
        RECT 140.320 122.010 140.490 122.190 ;
        RECT 140.800 122.010 140.970 122.190 ;
        RECT 141.280 122.010 141.450 122.190 ;
      LAYER li1 ;
        RECT 141.600 122.180 142.080 122.190 ;
      LAYER li1 ;
        RECT 141.760 122.010 141.930 122.180 ;
        RECT 6.470 121.590 6.640 121.760 ;
        RECT 6.910 121.590 7.080 121.760 ;
        RECT 7.320 121.590 7.490 121.760 ;
        RECT 7.750 121.590 7.920 121.760 ;
        RECT 8.190 121.590 8.360 121.760 ;
        RECT 8.600 121.590 8.770 121.760 ;
        RECT 11.160 121.540 11.330 121.710 ;
        RECT 11.520 121.540 11.690 121.710 ;
        RECT 13.190 121.590 13.360 121.760 ;
        RECT 13.630 121.590 13.800 121.760 ;
        RECT 14.040 121.590 14.210 121.760 ;
        RECT 14.470 121.590 14.640 121.760 ;
        RECT 14.910 121.590 15.080 121.760 ;
        RECT 15.320 121.590 15.490 121.760 ;
        RECT 17.030 121.590 17.200 121.760 ;
        RECT 17.470 121.590 17.640 121.760 ;
        RECT 17.880 121.590 18.050 121.760 ;
        RECT 18.310 121.590 18.480 121.760 ;
        RECT 18.750 121.590 18.920 121.760 ;
        RECT 19.160 121.590 19.330 121.760 ;
        RECT 20.730 121.540 20.900 121.710 ;
        RECT 21.090 121.540 21.260 121.710 ;
        RECT 21.450 121.540 21.620 121.710 ;
        RECT 23.900 121.540 24.070 121.710 ;
        RECT 24.260 121.540 24.430 121.710 ;
        RECT 24.620 121.540 24.790 121.710 ;
        RECT 25.940 121.590 26.110 121.760 ;
        RECT 26.300 121.590 26.470 121.760 ;
        RECT 26.740 121.590 26.910 121.760 ;
        RECT 29.370 121.540 29.540 121.710 ;
        RECT 29.730 121.540 29.900 121.710 ;
        RECT 30.090 121.540 30.260 121.710 ;
        RECT 32.540 121.540 32.710 121.710 ;
        RECT 32.900 121.540 33.070 121.710 ;
        RECT 33.260 121.540 33.430 121.710 ;
        RECT 34.580 121.590 34.750 121.760 ;
        RECT 34.940 121.590 35.110 121.760 ;
        RECT 35.380 121.590 35.550 121.760 ;
        RECT 36.740 121.540 36.910 121.710 ;
        RECT 37.100 121.540 37.270 121.710 ;
        RECT 39.110 121.590 39.280 121.760 ;
        RECT 39.550 121.590 39.720 121.760 ;
        RECT 39.960 121.590 40.130 121.760 ;
        RECT 40.390 121.590 40.560 121.760 ;
        RECT 40.830 121.590 41.000 121.760 ;
        RECT 41.240 121.590 41.410 121.760 ;
        RECT 44.420 121.540 44.590 121.710 ;
        RECT 44.780 121.540 44.950 121.710 ;
        RECT 46.790 121.590 46.960 121.760 ;
        RECT 47.230 121.590 47.400 121.760 ;
        RECT 47.640 121.590 47.810 121.760 ;
        RECT 48.070 121.590 48.240 121.760 ;
        RECT 48.510 121.590 48.680 121.760 ;
        RECT 48.920 121.590 49.090 121.760 ;
        RECT 50.980 121.540 51.150 121.710 ;
        RECT 51.340 121.540 51.510 121.710 ;
        RECT 51.700 121.540 51.870 121.710 ;
        RECT 52.670 121.540 52.840 121.710 ;
        RECT 56.040 121.540 56.210 121.710 ;
        RECT 57.510 121.540 57.680 121.710 ;
        RECT 57.870 121.540 58.040 121.710 ;
        RECT 58.230 121.540 58.400 121.710 ;
        RECT 60.440 121.540 60.610 121.710 ;
        RECT 60.800 121.540 60.970 121.710 ;
        RECT 61.160 121.540 61.330 121.710 ;
        RECT 62.160 121.540 62.330 121.710 ;
        RECT 62.520 121.540 62.690 121.710 ;
        RECT 62.880 121.540 63.050 121.710 ;
        RECT 63.720 121.540 63.890 121.710 ;
        RECT 64.080 121.540 64.250 121.710 ;
        RECT 64.440 121.540 64.610 121.710 ;
        RECT 65.780 121.590 65.950 121.760 ;
        RECT 66.140 121.590 66.310 121.760 ;
        RECT 66.580 121.590 66.750 121.760 ;
        RECT 67.800 121.540 67.970 121.710 ;
        RECT 68.160 121.540 68.330 121.710 ;
        RECT 69.830 121.590 70.000 121.760 ;
        RECT 70.270 121.590 70.440 121.760 ;
        RECT 70.680 121.590 70.850 121.760 ;
        RECT 71.110 121.590 71.280 121.760 ;
        RECT 71.550 121.590 71.720 121.760 ;
        RECT 71.960 121.590 72.130 121.760 ;
        RECT 74.660 121.540 74.830 121.710 ;
        RECT 75.020 121.540 75.190 121.710 ;
        RECT 76.820 121.590 76.990 121.760 ;
        RECT 77.180 121.590 77.350 121.760 ;
        RECT 77.620 121.590 77.790 121.760 ;
        RECT 78.360 121.540 78.530 121.710 ;
        RECT 78.720 121.540 78.890 121.710 ;
        RECT 79.080 121.540 79.250 121.710 ;
        RECT 79.440 121.540 79.610 121.710 ;
        RECT 79.800 121.540 79.970 121.710 ;
        RECT 81.140 121.590 81.310 121.760 ;
        RECT 81.500 121.590 81.670 121.760 ;
        RECT 81.940 121.590 82.110 121.760 ;
        RECT 82.680 121.540 82.850 121.710 ;
        RECT 83.040 121.540 83.210 121.710 ;
        RECT 84.500 121.590 84.670 121.760 ;
        RECT 84.860 121.590 85.030 121.760 ;
        RECT 85.300 121.590 85.470 121.760 ;
        RECT 86.040 121.540 86.210 121.710 ;
        RECT 86.400 121.540 86.570 121.710 ;
        RECT 86.760 121.540 86.930 121.710 ;
        RECT 87.610 121.540 87.780 121.710 ;
        RECT 87.970 121.540 88.140 121.710 ;
        RECT 88.820 121.590 88.990 121.760 ;
        RECT 89.180 121.590 89.350 121.760 ;
        RECT 89.620 121.590 89.790 121.760 ;
        RECT 90.360 121.540 90.530 121.710 ;
        RECT 90.720 121.540 90.890 121.710 ;
        RECT 91.080 121.540 91.250 121.710 ;
        RECT 91.440 121.540 91.610 121.710 ;
        RECT 91.800 121.540 91.970 121.710 ;
        RECT 93.140 121.590 93.310 121.760 ;
        RECT 93.500 121.590 93.670 121.760 ;
        RECT 93.940 121.590 94.110 121.760 ;
        RECT 96.730 121.540 96.900 121.710 ;
        RECT 97.090 121.540 97.260 121.710 ;
        RECT 97.450 121.540 97.620 121.710 ;
        RECT 98.900 121.590 99.070 121.760 ;
        RECT 99.260 121.590 99.430 121.760 ;
        RECT 99.700 121.590 99.870 121.760 ;
        RECT 100.920 121.540 101.090 121.710 ;
        RECT 101.280 121.540 101.450 121.710 ;
        RECT 102.740 121.590 102.910 121.760 ;
        RECT 103.100 121.590 103.270 121.760 ;
        RECT 103.540 121.590 103.710 121.760 ;
        RECT 104.260 121.540 104.430 121.710 ;
        RECT 104.620 121.540 104.790 121.710 ;
        RECT 104.980 121.540 105.150 121.710 ;
        RECT 105.340 121.540 105.510 121.710 ;
        RECT 106.500 121.540 106.670 121.710 ;
        RECT 106.860 121.540 107.030 121.710 ;
        RECT 107.220 121.540 107.390 121.710 ;
        RECT 107.580 121.540 107.750 121.710 ;
        RECT 108.710 121.590 108.880 121.760 ;
        RECT 109.150 121.590 109.320 121.760 ;
        RECT 109.560 121.590 109.730 121.760 ;
        RECT 109.990 121.590 110.160 121.760 ;
        RECT 110.430 121.590 110.600 121.760 ;
        RECT 110.840 121.590 111.010 121.760 ;
        RECT 112.550 121.590 112.720 121.760 ;
        RECT 112.990 121.590 113.160 121.760 ;
        RECT 113.400 121.590 113.570 121.760 ;
        RECT 113.830 121.590 114.000 121.760 ;
        RECT 114.270 121.590 114.440 121.760 ;
        RECT 114.680 121.590 114.850 121.760 ;
        RECT 116.390 121.590 116.560 121.760 ;
        RECT 116.830 121.590 117.000 121.760 ;
        RECT 117.240 121.590 117.410 121.760 ;
        RECT 117.670 121.590 117.840 121.760 ;
        RECT 118.110 121.590 118.280 121.760 ;
        RECT 118.520 121.590 118.690 121.760 ;
        RECT 120.230 121.590 120.400 121.760 ;
        RECT 120.670 121.590 120.840 121.760 ;
        RECT 121.080 121.590 121.250 121.760 ;
        RECT 121.510 121.590 121.680 121.760 ;
        RECT 121.950 121.590 122.120 121.760 ;
        RECT 122.360 121.590 122.530 121.760 ;
        RECT 124.070 121.590 124.240 121.760 ;
        RECT 124.510 121.590 124.680 121.760 ;
        RECT 124.920 121.590 125.090 121.760 ;
        RECT 125.350 121.590 125.520 121.760 ;
        RECT 125.790 121.590 125.960 121.760 ;
        RECT 126.200 121.590 126.370 121.760 ;
        RECT 127.910 121.590 128.080 121.760 ;
        RECT 128.350 121.590 128.520 121.760 ;
        RECT 128.760 121.590 128.930 121.760 ;
        RECT 129.190 121.590 129.360 121.760 ;
        RECT 129.630 121.590 129.800 121.760 ;
        RECT 130.040 121.590 130.210 121.760 ;
        RECT 131.750 121.590 131.920 121.760 ;
        RECT 132.190 121.590 132.360 121.760 ;
        RECT 132.600 121.590 132.770 121.760 ;
        RECT 133.030 121.590 133.200 121.760 ;
        RECT 133.470 121.590 133.640 121.760 ;
        RECT 133.880 121.590 134.050 121.760 ;
        RECT 135.590 121.590 135.760 121.760 ;
        RECT 136.030 121.590 136.200 121.760 ;
        RECT 136.440 121.590 136.610 121.760 ;
        RECT 136.870 121.590 137.040 121.760 ;
        RECT 137.310 121.590 137.480 121.760 ;
        RECT 137.720 121.590 137.890 121.760 ;
        RECT 139.220 121.590 139.390 121.760 ;
        RECT 139.580 121.590 139.750 121.760 ;
        RECT 140.020 121.590 140.190 121.760 ;
        RECT 6.470 114.300 6.640 114.470 ;
        RECT 6.910 114.300 7.080 114.470 ;
        RECT 7.320 114.300 7.490 114.470 ;
        RECT 7.750 114.300 7.920 114.470 ;
        RECT 8.190 114.300 8.360 114.470 ;
        RECT 8.600 114.300 8.770 114.470 ;
        RECT 10.310 114.300 10.480 114.470 ;
        RECT 10.750 114.300 10.920 114.470 ;
        RECT 11.160 114.300 11.330 114.470 ;
        RECT 11.590 114.300 11.760 114.470 ;
        RECT 12.030 114.300 12.200 114.470 ;
        RECT 12.440 114.300 12.610 114.470 ;
        RECT 14.660 114.350 14.830 114.520 ;
        RECT 15.020 114.350 15.190 114.520 ;
        RECT 17.030 114.300 17.200 114.470 ;
        RECT 17.470 114.300 17.640 114.470 ;
        RECT 17.880 114.300 18.050 114.470 ;
        RECT 18.310 114.300 18.480 114.470 ;
        RECT 18.750 114.300 18.920 114.470 ;
        RECT 19.160 114.300 19.330 114.470 ;
        RECT 20.870 114.300 21.040 114.470 ;
        RECT 21.310 114.300 21.480 114.470 ;
        RECT 21.720 114.300 21.890 114.470 ;
        RECT 22.150 114.300 22.320 114.470 ;
        RECT 22.590 114.300 22.760 114.470 ;
        RECT 23.000 114.300 23.170 114.470 ;
        RECT 25.080 114.350 25.250 114.520 ;
        RECT 25.440 114.350 25.610 114.520 ;
        RECT 27.110 114.300 27.280 114.470 ;
        RECT 27.550 114.300 27.720 114.470 ;
        RECT 27.960 114.300 28.130 114.470 ;
        RECT 28.390 114.300 28.560 114.470 ;
        RECT 28.830 114.300 29.000 114.470 ;
        RECT 29.240 114.300 29.410 114.470 ;
        RECT 30.950 114.300 31.120 114.470 ;
        RECT 31.390 114.300 31.560 114.470 ;
        RECT 31.800 114.300 31.970 114.470 ;
        RECT 32.230 114.300 32.400 114.470 ;
        RECT 32.670 114.300 32.840 114.470 ;
        RECT 33.080 114.300 33.250 114.470 ;
        RECT 34.790 114.300 34.960 114.470 ;
        RECT 35.230 114.300 35.400 114.470 ;
        RECT 35.640 114.300 35.810 114.470 ;
        RECT 36.070 114.300 36.240 114.470 ;
        RECT 36.510 114.300 36.680 114.470 ;
        RECT 36.920 114.300 37.090 114.470 ;
        RECT 38.630 114.300 38.800 114.470 ;
        RECT 39.070 114.300 39.240 114.470 ;
        RECT 39.480 114.300 39.650 114.470 ;
        RECT 39.910 114.300 40.080 114.470 ;
        RECT 40.350 114.300 40.520 114.470 ;
        RECT 40.760 114.300 40.930 114.470 ;
        RECT 42.820 114.350 42.990 114.520 ;
        RECT 43.180 114.350 43.350 114.520 ;
        RECT 43.540 114.350 43.710 114.520 ;
        RECT 43.900 114.350 44.070 114.520 ;
        RECT 45.060 114.350 45.230 114.520 ;
        RECT 45.420 114.350 45.590 114.520 ;
        RECT 45.780 114.350 45.950 114.520 ;
        RECT 46.140 114.350 46.310 114.520 ;
        RECT 47.060 114.300 47.230 114.470 ;
        RECT 47.420 114.300 47.590 114.470 ;
        RECT 47.860 114.300 48.030 114.470 ;
        RECT 48.600 114.350 48.770 114.520 ;
        RECT 48.960 114.350 49.130 114.520 ;
        RECT 49.320 114.350 49.490 114.520 ;
        RECT 50.160 114.350 50.330 114.520 ;
        RECT 50.520 114.350 50.690 114.520 ;
        RECT 50.880 114.350 51.050 114.520 ;
        RECT 51.800 114.350 51.970 114.520 ;
        RECT 52.160 114.350 52.330 114.520 ;
        RECT 52.520 114.350 52.690 114.520 ;
        RECT 53.780 114.300 53.950 114.470 ;
        RECT 54.140 114.300 54.310 114.470 ;
        RECT 54.580 114.300 54.750 114.470 ;
        RECT 56.900 114.350 57.070 114.520 ;
        RECT 57.260 114.350 57.430 114.520 ;
        RECT 59.060 114.300 59.230 114.470 ;
        RECT 59.420 114.300 59.590 114.470 ;
        RECT 59.860 114.300 60.030 114.470 ;
        RECT 61.220 114.350 61.390 114.520 ;
        RECT 61.580 114.350 61.750 114.520 ;
        RECT 63.590 114.300 63.760 114.470 ;
        RECT 64.030 114.300 64.200 114.470 ;
        RECT 64.440 114.300 64.610 114.470 ;
        RECT 64.870 114.300 65.040 114.470 ;
        RECT 65.310 114.300 65.480 114.470 ;
        RECT 65.720 114.300 65.890 114.470 ;
        RECT 67.460 114.350 67.630 114.520 ;
        RECT 67.820 114.350 67.990 114.520 ;
        RECT 69.620 114.300 69.790 114.470 ;
        RECT 69.980 114.300 70.150 114.470 ;
        RECT 70.420 114.300 70.590 114.470 ;
        RECT 71.700 114.350 71.870 114.520 ;
        RECT 72.060 114.350 72.230 114.520 ;
        RECT 74.090 114.350 74.260 114.520 ;
        RECT 76.520 114.350 76.690 114.520 ;
        RECT 76.880 114.350 77.050 114.520 ;
        RECT 77.240 114.350 77.410 114.520 ;
        RECT 78.860 114.350 79.030 114.520 ;
        RECT 79.220 114.350 79.390 114.520 ;
        RECT 79.580 114.350 79.750 114.520 ;
        RECT 81.560 114.350 81.730 114.520 ;
        RECT 81.920 114.350 82.090 114.520 ;
        RECT 82.280 114.350 82.450 114.520 ;
        RECT 83.310 114.350 83.480 114.520 ;
        RECT 83.670 114.350 83.840 114.520 ;
        RECT 84.030 114.350 84.200 114.520 ;
        RECT 84.840 114.350 85.010 114.520 ;
        RECT 85.200 114.350 85.370 114.520 ;
        RECT 85.560 114.350 85.730 114.520 ;
        RECT 86.900 114.300 87.070 114.470 ;
        RECT 87.260 114.300 87.430 114.470 ;
        RECT 87.700 114.300 87.870 114.470 ;
        RECT 89.540 114.350 89.710 114.520 ;
        RECT 89.900 114.350 90.070 114.520 ;
        RECT 91.700 114.300 91.870 114.470 ;
        RECT 92.060 114.300 92.230 114.470 ;
        RECT 92.500 114.300 92.670 114.470 ;
        RECT 93.680 114.350 93.850 114.520 ;
        RECT 94.040 114.350 94.210 114.520 ;
        RECT 94.400 114.350 94.570 114.520 ;
        RECT 94.760 114.350 94.930 114.520 ;
        RECT 95.120 114.350 95.290 114.520 ;
        RECT 95.480 114.350 95.650 114.520 ;
        RECT 95.840 114.350 96.010 114.520 ;
        RECT 96.200 114.350 96.370 114.520 ;
        RECT 97.010 114.350 97.180 114.520 ;
        RECT 97.370 114.350 97.540 114.520 ;
        RECT 97.730 114.350 97.900 114.520 ;
        RECT 98.090 114.350 98.260 114.520 ;
        RECT 98.900 114.300 99.070 114.470 ;
        RECT 99.260 114.300 99.430 114.470 ;
        RECT 99.700 114.300 99.870 114.470 ;
        RECT 101.060 114.350 101.230 114.520 ;
        RECT 101.420 114.350 101.590 114.520 ;
        RECT 103.220 114.300 103.390 114.470 ;
        RECT 103.580 114.300 103.750 114.470 ;
        RECT 104.020 114.300 104.190 114.470 ;
        RECT 104.760 114.350 104.930 114.520 ;
        RECT 105.120 114.350 105.290 114.520 ;
        RECT 105.480 114.350 105.650 114.520 ;
        RECT 106.320 114.350 106.490 114.520 ;
        RECT 106.680 114.350 106.850 114.520 ;
        RECT 107.040 114.350 107.210 114.520 ;
        RECT 107.960 114.350 108.130 114.520 ;
        RECT 108.320 114.350 108.490 114.520 ;
        RECT 108.680 114.350 108.850 114.520 ;
        RECT 109.940 114.300 110.110 114.470 ;
        RECT 110.300 114.300 110.470 114.470 ;
        RECT 110.740 114.300 110.910 114.470 ;
        RECT 112.100 114.350 112.270 114.520 ;
        RECT 112.460 114.350 112.630 114.520 ;
        RECT 114.260 114.300 114.430 114.470 ;
        RECT 114.620 114.300 114.790 114.470 ;
        RECT 115.060 114.300 115.230 114.470 ;
        RECT 117.860 114.350 118.030 114.520 ;
        RECT 118.220 114.350 118.390 114.520 ;
        RECT 120.020 114.300 120.190 114.470 ;
        RECT 120.380 114.300 120.550 114.470 ;
        RECT 120.820 114.300 120.990 114.470 ;
        RECT 121.560 114.350 121.730 114.520 ;
        RECT 121.920 114.350 122.090 114.520 ;
        RECT 123.590 114.300 123.760 114.470 ;
        RECT 124.030 114.300 124.200 114.470 ;
        RECT 124.440 114.300 124.610 114.470 ;
        RECT 124.870 114.300 125.040 114.470 ;
        RECT 125.310 114.300 125.480 114.470 ;
        RECT 125.720 114.300 125.890 114.470 ;
        RECT 127.430 114.300 127.600 114.470 ;
        RECT 127.870 114.300 128.040 114.470 ;
        RECT 128.280 114.300 128.450 114.470 ;
        RECT 128.710 114.300 128.880 114.470 ;
        RECT 129.150 114.300 129.320 114.470 ;
        RECT 129.560 114.300 129.730 114.470 ;
        RECT 131.270 114.300 131.440 114.470 ;
        RECT 131.710 114.300 131.880 114.470 ;
        RECT 132.120 114.300 132.290 114.470 ;
        RECT 132.550 114.300 132.720 114.470 ;
        RECT 132.990 114.300 133.160 114.470 ;
        RECT 133.400 114.300 133.570 114.470 ;
        RECT 135.110 114.300 135.280 114.470 ;
        RECT 135.550 114.300 135.720 114.470 ;
        RECT 135.960 114.300 136.130 114.470 ;
        RECT 136.390 114.300 136.560 114.470 ;
        RECT 136.830 114.300 137.000 114.470 ;
        RECT 137.240 114.300 137.410 114.470 ;
        RECT 138.950 114.300 139.120 114.470 ;
        RECT 139.390 114.300 139.560 114.470 ;
        RECT 139.800 114.300 139.970 114.470 ;
        RECT 140.230 114.300 140.400 114.470 ;
        RECT 140.670 114.300 140.840 114.470 ;
        RECT 141.080 114.300 141.250 114.470 ;
        RECT 5.920 113.870 6.090 114.050 ;
        RECT 6.400 113.870 6.570 114.050 ;
        RECT 6.880 113.870 7.050 114.050 ;
        RECT 7.360 113.870 7.530 114.050 ;
        RECT 7.840 113.870 8.010 114.050 ;
        RECT 8.320 113.870 8.490 114.050 ;
        RECT 8.800 113.870 8.970 114.050 ;
        RECT 9.280 113.870 9.450 114.050 ;
        RECT 9.760 113.870 9.930 114.050 ;
        RECT 10.240 113.870 10.410 114.050 ;
        RECT 10.720 113.870 10.890 114.050 ;
        RECT 11.200 113.870 11.370 114.050 ;
        RECT 11.680 113.870 11.850 114.050 ;
        RECT 12.160 113.870 12.330 114.050 ;
        RECT 12.640 113.870 12.810 114.050 ;
        RECT 13.120 113.870 13.290 114.050 ;
        RECT 13.600 114.040 13.770 114.050 ;
      LAYER li1 ;
        RECT 13.440 113.870 13.920 114.040 ;
      LAYER li1 ;
        RECT 14.080 113.870 14.250 114.050 ;
        RECT 14.560 113.870 14.730 114.050 ;
        RECT 15.040 113.870 15.210 114.050 ;
        RECT 15.520 113.870 15.690 114.050 ;
        RECT 16.000 113.870 16.170 114.050 ;
        RECT 16.480 113.870 16.650 114.050 ;
        RECT 16.960 113.870 17.130 114.050 ;
        RECT 17.440 113.870 17.610 114.050 ;
        RECT 17.920 113.870 18.090 114.050 ;
        RECT 18.400 113.870 18.570 114.050 ;
        RECT 18.880 113.870 19.050 114.050 ;
        RECT 19.360 113.870 19.530 114.050 ;
        RECT 19.840 113.870 20.010 114.050 ;
        RECT 20.320 113.870 20.490 114.050 ;
        RECT 20.800 113.870 20.970 114.050 ;
        RECT 21.280 113.870 21.450 114.050 ;
        RECT 21.760 113.870 21.930 114.050 ;
        RECT 22.240 113.870 22.410 114.050 ;
        RECT 22.720 113.870 22.890 114.050 ;
        RECT 23.200 113.870 23.370 114.050 ;
        RECT 23.680 113.870 23.850 114.050 ;
      LAYER li1 ;
        RECT 24.000 114.040 24.480 114.050 ;
      LAYER li1 ;
        RECT 24.160 113.870 24.330 114.040 ;
        RECT 24.640 113.870 24.810 114.050 ;
        RECT 25.120 113.870 25.290 114.050 ;
        RECT 25.600 113.870 25.770 114.050 ;
        RECT 26.080 113.870 26.250 114.050 ;
        RECT 26.560 113.870 26.730 114.050 ;
        RECT 27.040 113.870 27.210 114.050 ;
        RECT 27.520 113.870 27.690 114.050 ;
        RECT 28.000 113.870 28.170 114.050 ;
        RECT 28.480 113.870 28.650 114.050 ;
        RECT 28.960 113.870 29.130 114.050 ;
        RECT 29.440 113.870 29.610 114.050 ;
        RECT 29.920 113.870 30.090 114.050 ;
        RECT 30.400 113.870 30.570 114.050 ;
        RECT 30.880 113.870 31.050 114.050 ;
        RECT 31.360 113.870 31.530 114.050 ;
        RECT 31.840 113.870 32.010 114.050 ;
        RECT 32.320 113.870 32.490 114.050 ;
        RECT 32.800 113.870 32.970 114.050 ;
        RECT 33.280 113.870 33.450 114.050 ;
        RECT 33.760 113.870 33.930 114.050 ;
        RECT 34.240 113.870 34.410 114.050 ;
        RECT 34.720 113.870 34.890 114.050 ;
        RECT 35.200 113.870 35.370 114.050 ;
        RECT 35.680 113.870 35.850 114.050 ;
        RECT 36.160 113.870 36.330 114.050 ;
        RECT 36.640 113.870 36.810 114.050 ;
      LAYER li1 ;
        RECT 36.960 114.040 37.440 114.050 ;
      LAYER li1 ;
        RECT 37.120 113.870 37.290 114.040 ;
        RECT 37.600 113.870 37.770 114.050 ;
        RECT 38.080 113.870 38.250 114.050 ;
        RECT 38.560 113.870 38.730 114.050 ;
        RECT 39.040 113.870 39.210 114.050 ;
        RECT 39.520 113.870 39.690 114.050 ;
        RECT 40.000 113.870 40.170 114.050 ;
        RECT 40.480 113.870 40.650 114.050 ;
        RECT 40.960 113.870 41.130 114.050 ;
        RECT 41.440 113.870 41.610 114.050 ;
        RECT 41.920 113.870 42.090 114.050 ;
        RECT 42.400 113.870 42.570 114.050 ;
        RECT 42.880 113.870 43.050 114.050 ;
        RECT 43.360 113.870 43.530 114.050 ;
        RECT 43.840 113.870 44.010 114.050 ;
        RECT 44.320 113.870 44.490 114.050 ;
        RECT 44.800 113.870 44.970 114.050 ;
        RECT 45.280 113.870 45.450 114.050 ;
        RECT 45.760 113.870 45.930 114.050 ;
        RECT 46.240 113.870 46.410 114.050 ;
        RECT 46.720 113.870 46.890 114.050 ;
        RECT 47.200 113.870 47.370 114.050 ;
        RECT 47.680 113.870 47.850 114.050 ;
        RECT 48.160 113.870 48.330 114.050 ;
        RECT 48.640 113.870 48.810 114.050 ;
        RECT 49.120 113.870 49.290 114.050 ;
        RECT 49.600 113.870 49.770 114.050 ;
        RECT 50.080 113.870 50.250 114.050 ;
        RECT 50.560 113.870 50.730 114.050 ;
        RECT 51.040 113.870 51.210 114.050 ;
        RECT 51.520 113.870 51.690 114.050 ;
        RECT 52.000 113.870 52.170 114.050 ;
        RECT 52.480 113.870 52.650 114.050 ;
        RECT 52.960 113.870 53.130 114.050 ;
        RECT 53.440 113.870 53.610 114.050 ;
        RECT 53.920 113.870 54.090 114.050 ;
        RECT 54.400 113.870 54.570 114.050 ;
        RECT 54.880 113.870 55.050 114.050 ;
        RECT 55.360 113.870 55.530 114.050 ;
        RECT 55.840 113.870 56.010 114.050 ;
        RECT 56.320 113.870 56.490 114.050 ;
        RECT 56.800 113.870 56.970 114.050 ;
        RECT 57.280 113.870 57.450 114.050 ;
        RECT 57.760 113.870 57.930 114.050 ;
        RECT 58.240 113.870 58.410 114.050 ;
        RECT 58.720 113.870 58.890 114.050 ;
        RECT 59.200 113.870 59.370 114.050 ;
        RECT 59.680 113.870 59.850 114.050 ;
        RECT 60.160 113.870 60.330 114.050 ;
        RECT 60.640 113.870 60.810 114.050 ;
        RECT 61.120 113.870 61.290 114.050 ;
        RECT 61.600 113.870 61.770 114.050 ;
        RECT 62.080 113.870 62.250 114.050 ;
        RECT 62.560 113.870 62.730 114.050 ;
        RECT 63.040 113.870 63.210 114.050 ;
        RECT 63.520 113.870 63.690 114.050 ;
        RECT 64.000 113.870 64.170 114.050 ;
        RECT 64.480 113.870 64.650 114.050 ;
        RECT 64.960 113.870 65.130 114.050 ;
        RECT 65.440 113.870 65.610 114.050 ;
        RECT 65.920 113.870 66.090 114.050 ;
        RECT 66.400 113.870 66.570 114.050 ;
        RECT 66.880 113.870 67.050 114.050 ;
        RECT 67.360 113.870 67.530 114.050 ;
        RECT 67.840 113.870 68.010 114.050 ;
        RECT 68.320 113.870 68.490 114.050 ;
        RECT 68.800 113.870 68.970 114.050 ;
        RECT 69.280 113.870 69.450 114.050 ;
        RECT 69.760 113.870 69.930 114.050 ;
        RECT 70.240 113.870 70.410 114.050 ;
        RECT 70.720 113.870 70.890 114.050 ;
        RECT 71.200 113.870 71.370 114.050 ;
      LAYER li1 ;
        RECT 71.520 114.040 72.000 114.050 ;
      LAYER li1 ;
        RECT 71.680 113.870 71.850 114.040 ;
        RECT 72.160 113.870 72.330 114.050 ;
        RECT 72.640 113.870 72.810 114.050 ;
        RECT 73.120 113.870 73.290 114.050 ;
        RECT 73.600 113.870 73.770 114.050 ;
        RECT 74.080 113.870 74.250 114.050 ;
        RECT 74.560 113.870 74.730 114.050 ;
        RECT 75.040 113.870 75.210 114.050 ;
        RECT 75.520 113.870 75.690 114.050 ;
        RECT 76.000 113.870 76.170 114.050 ;
        RECT 76.480 113.870 76.650 114.050 ;
        RECT 76.960 113.870 77.130 114.050 ;
        RECT 77.440 113.870 77.610 114.050 ;
        RECT 77.920 113.870 78.090 114.050 ;
        RECT 78.400 113.870 78.570 114.050 ;
        RECT 78.880 113.870 79.050 114.050 ;
        RECT 79.360 113.870 79.530 114.050 ;
        RECT 79.840 113.870 80.010 114.050 ;
        RECT 80.320 113.870 80.490 114.050 ;
        RECT 80.800 113.870 80.970 114.050 ;
        RECT 81.280 113.870 81.450 114.050 ;
        RECT 81.760 113.870 81.930 114.050 ;
        RECT 82.240 113.870 82.410 114.050 ;
        RECT 82.720 113.870 82.890 114.050 ;
        RECT 83.200 113.870 83.370 114.050 ;
        RECT 83.680 113.870 83.850 114.050 ;
        RECT 84.160 113.870 84.330 114.050 ;
        RECT 84.640 113.870 84.810 114.050 ;
        RECT 85.120 113.870 85.290 114.050 ;
        RECT 85.600 113.870 85.770 114.050 ;
        RECT 86.080 113.870 86.250 114.050 ;
        RECT 86.560 113.870 86.730 114.050 ;
        RECT 87.040 113.870 87.210 114.050 ;
        RECT 87.520 113.870 87.690 114.050 ;
        RECT 88.000 113.870 88.170 114.050 ;
        RECT 88.480 114.040 88.650 114.050 ;
      LAYER li1 ;
        RECT 88.320 113.870 88.800 114.040 ;
      LAYER li1 ;
        RECT 88.960 113.870 89.130 114.050 ;
        RECT 89.440 113.870 89.610 114.050 ;
        RECT 89.920 113.870 90.090 114.050 ;
        RECT 90.400 113.870 90.570 114.050 ;
        RECT 90.880 113.870 91.050 114.050 ;
        RECT 91.360 113.870 91.530 114.050 ;
        RECT 91.840 113.870 92.010 114.050 ;
        RECT 92.320 113.870 92.490 114.050 ;
        RECT 92.800 113.870 92.970 114.050 ;
        RECT 93.280 113.870 93.450 114.050 ;
        RECT 93.760 113.870 93.930 114.050 ;
        RECT 94.240 113.870 94.410 114.050 ;
        RECT 94.720 113.870 94.890 114.050 ;
        RECT 95.200 113.870 95.370 114.050 ;
        RECT 95.680 113.870 95.850 114.050 ;
        RECT 96.160 113.870 96.330 114.050 ;
        RECT 96.640 113.870 96.810 114.050 ;
        RECT 97.120 113.870 97.290 114.050 ;
        RECT 97.600 113.870 97.770 114.050 ;
        RECT 98.080 113.870 98.250 114.050 ;
        RECT 98.560 113.870 98.730 114.050 ;
        RECT 99.040 113.870 99.210 114.050 ;
        RECT 99.520 113.870 99.690 114.050 ;
        RECT 100.000 113.870 100.170 114.050 ;
        RECT 100.480 113.870 100.650 114.050 ;
        RECT 100.960 113.870 101.130 114.050 ;
        RECT 101.440 113.870 101.610 114.050 ;
        RECT 101.920 113.870 102.090 114.050 ;
        RECT 102.400 113.870 102.570 114.050 ;
        RECT 102.880 113.870 103.050 114.050 ;
        RECT 103.360 113.870 103.530 114.050 ;
        RECT 103.840 113.870 104.010 114.050 ;
        RECT 104.320 113.870 104.490 114.050 ;
        RECT 104.800 113.870 104.970 114.050 ;
        RECT 105.280 113.870 105.450 114.050 ;
        RECT 105.760 113.870 105.930 114.050 ;
        RECT 106.240 113.870 106.410 114.050 ;
        RECT 106.720 113.870 106.890 114.050 ;
        RECT 107.200 113.870 107.370 114.050 ;
        RECT 107.680 113.870 107.850 114.050 ;
        RECT 108.160 113.870 108.330 114.050 ;
        RECT 108.640 113.870 108.810 114.050 ;
        RECT 109.120 113.870 109.290 114.050 ;
        RECT 109.600 113.870 109.770 114.050 ;
        RECT 110.080 113.870 110.250 114.050 ;
        RECT 110.560 113.870 110.730 114.050 ;
        RECT 111.040 113.870 111.210 114.050 ;
        RECT 111.520 113.870 111.690 114.050 ;
        RECT 112.000 113.870 112.170 114.050 ;
        RECT 112.480 113.870 112.650 114.050 ;
        RECT 112.960 113.870 113.130 114.050 ;
        RECT 113.440 113.870 113.610 114.050 ;
        RECT 113.920 113.870 114.090 114.050 ;
        RECT 114.400 113.870 114.570 114.050 ;
        RECT 114.880 113.870 115.050 114.050 ;
        RECT 115.360 113.870 115.530 114.050 ;
        RECT 115.840 113.870 116.010 114.050 ;
        RECT 116.320 113.870 116.490 114.050 ;
        RECT 116.800 114.040 116.970 114.050 ;
      LAYER li1 ;
        RECT 116.640 113.870 117.120 114.040 ;
      LAYER li1 ;
        RECT 117.280 113.870 117.450 114.050 ;
        RECT 117.760 113.870 117.930 114.050 ;
        RECT 118.240 113.870 118.410 114.050 ;
        RECT 118.720 113.870 118.890 114.050 ;
        RECT 119.200 113.870 119.370 114.050 ;
        RECT 119.680 113.870 119.850 114.050 ;
        RECT 120.160 113.870 120.330 114.050 ;
        RECT 120.640 113.870 120.810 114.050 ;
        RECT 121.120 113.870 121.290 114.050 ;
        RECT 121.600 113.870 121.770 114.050 ;
        RECT 122.080 113.870 122.250 114.050 ;
        RECT 122.560 113.870 122.730 114.050 ;
        RECT 123.040 113.870 123.210 114.050 ;
        RECT 123.520 113.870 123.690 114.050 ;
        RECT 124.000 113.870 124.170 114.050 ;
        RECT 124.480 113.870 124.650 114.050 ;
        RECT 124.960 113.870 125.130 114.050 ;
        RECT 125.440 113.870 125.610 114.050 ;
        RECT 125.920 113.870 126.090 114.050 ;
        RECT 126.400 113.870 126.570 114.050 ;
        RECT 126.880 113.870 127.050 114.050 ;
        RECT 127.360 113.870 127.530 114.050 ;
        RECT 127.840 113.870 128.010 114.050 ;
        RECT 128.320 113.870 128.490 114.050 ;
        RECT 128.800 113.870 128.970 114.050 ;
        RECT 129.280 113.870 129.450 114.050 ;
        RECT 129.760 113.870 129.930 114.050 ;
        RECT 130.240 113.870 130.410 114.050 ;
        RECT 130.720 113.870 130.890 114.050 ;
        RECT 131.200 113.870 131.370 114.050 ;
        RECT 131.680 113.870 131.850 114.050 ;
        RECT 132.160 113.870 132.330 114.050 ;
        RECT 132.640 113.870 132.810 114.050 ;
        RECT 133.120 113.870 133.290 114.050 ;
        RECT 133.600 113.870 133.770 114.050 ;
        RECT 134.080 113.870 134.250 114.050 ;
        RECT 134.560 113.870 134.730 114.050 ;
        RECT 135.040 113.870 135.210 114.050 ;
        RECT 135.520 113.870 135.690 114.050 ;
        RECT 136.000 113.870 136.170 114.050 ;
        RECT 136.480 113.870 136.650 114.050 ;
        RECT 136.960 113.870 137.130 114.050 ;
        RECT 137.440 113.870 137.610 114.050 ;
        RECT 137.920 113.870 138.090 114.050 ;
        RECT 138.400 113.870 138.570 114.050 ;
        RECT 138.880 113.870 139.050 114.050 ;
        RECT 139.360 113.870 139.530 114.050 ;
        RECT 139.840 113.870 140.010 114.050 ;
        RECT 140.320 113.870 140.490 114.050 ;
        RECT 140.800 113.870 140.970 114.050 ;
        RECT 141.280 113.870 141.450 114.050 ;
        RECT 141.760 113.870 141.930 114.050 ;
        RECT 6.420 113.400 6.590 113.570 ;
        RECT 6.780 113.400 6.950 113.570 ;
        RECT 8.810 113.400 8.980 113.570 ;
        RECT 11.240 113.400 11.410 113.570 ;
        RECT 11.600 113.400 11.770 113.570 ;
        RECT 11.960 113.400 12.130 113.570 ;
        RECT 13.580 113.400 13.750 113.570 ;
        RECT 13.940 113.400 14.110 113.570 ;
        RECT 14.300 113.400 14.470 113.570 ;
        RECT 16.280 113.400 16.450 113.570 ;
        RECT 16.640 113.400 16.810 113.570 ;
        RECT 17.000 113.400 17.170 113.570 ;
        RECT 18.030 113.400 18.200 113.570 ;
        RECT 18.390 113.400 18.560 113.570 ;
        RECT 18.750 113.400 18.920 113.570 ;
        RECT 19.560 113.400 19.730 113.570 ;
        RECT 19.920 113.400 20.090 113.570 ;
        RECT 20.280 113.400 20.450 113.570 ;
        RECT 21.620 113.450 21.790 113.620 ;
        RECT 21.980 113.450 22.150 113.620 ;
        RECT 22.420 113.450 22.590 113.620 ;
        RECT 24.580 113.400 24.750 113.570 ;
        RECT 24.940 113.400 25.110 113.570 ;
        RECT 25.300 113.400 25.470 113.570 ;
        RECT 25.660 113.400 25.830 113.570 ;
        RECT 26.820 113.400 26.990 113.570 ;
        RECT 27.180 113.400 27.350 113.570 ;
        RECT 27.540 113.400 27.710 113.570 ;
        RECT 27.900 113.400 28.070 113.570 ;
        RECT 29.030 113.450 29.200 113.620 ;
        RECT 29.470 113.450 29.640 113.620 ;
        RECT 29.880 113.450 30.050 113.620 ;
        RECT 30.310 113.450 30.480 113.620 ;
        RECT 30.750 113.450 30.920 113.620 ;
        RECT 31.160 113.450 31.330 113.620 ;
        RECT 32.870 113.450 33.040 113.620 ;
        RECT 33.310 113.450 33.480 113.620 ;
        RECT 33.720 113.450 33.890 113.620 ;
        RECT 34.150 113.450 34.320 113.620 ;
        RECT 34.590 113.450 34.760 113.620 ;
        RECT 35.000 113.450 35.170 113.620 ;
        RECT 38.180 113.400 38.350 113.570 ;
        RECT 38.540 113.400 38.710 113.570 ;
        RECT 40.340 113.450 40.510 113.620 ;
        RECT 40.700 113.450 40.870 113.620 ;
        RECT 41.140 113.450 41.310 113.620 ;
        RECT 41.880 113.400 42.050 113.570 ;
        RECT 42.240 113.400 42.410 113.570 ;
        RECT 42.600 113.400 42.770 113.570 ;
        RECT 43.440 113.400 43.610 113.570 ;
        RECT 43.800 113.400 43.970 113.570 ;
        RECT 44.160 113.400 44.330 113.570 ;
        RECT 45.080 113.400 45.250 113.570 ;
        RECT 45.440 113.400 45.610 113.570 ;
        RECT 45.800 113.400 45.970 113.570 ;
        RECT 47.060 113.450 47.230 113.620 ;
        RECT 47.420 113.450 47.590 113.620 ;
        RECT 47.860 113.450 48.030 113.620 ;
        RECT 48.600 113.400 48.770 113.570 ;
        RECT 48.960 113.400 49.130 113.570 ;
        RECT 49.320 113.400 49.490 113.570 ;
        RECT 50.160 113.400 50.330 113.570 ;
        RECT 50.520 113.400 50.690 113.570 ;
        RECT 50.880 113.400 51.050 113.570 ;
        RECT 51.800 113.400 51.970 113.570 ;
        RECT 52.160 113.400 52.330 113.570 ;
        RECT 52.520 113.400 52.690 113.570 ;
        RECT 53.780 113.450 53.950 113.620 ;
        RECT 54.140 113.450 54.310 113.620 ;
        RECT 54.580 113.450 54.750 113.620 ;
        RECT 55.320 113.400 55.490 113.570 ;
        RECT 55.680 113.400 55.850 113.570 ;
        RECT 56.040 113.400 56.210 113.570 ;
        RECT 56.880 113.400 57.050 113.570 ;
        RECT 57.240 113.400 57.410 113.570 ;
        RECT 57.600 113.400 57.770 113.570 ;
        RECT 58.520 113.400 58.690 113.570 ;
        RECT 58.880 113.400 59.050 113.570 ;
        RECT 59.240 113.400 59.410 113.570 ;
        RECT 60.500 113.450 60.670 113.620 ;
        RECT 60.860 113.450 61.030 113.620 ;
        RECT 61.300 113.450 61.470 113.620 ;
        RECT 63.000 113.400 63.170 113.570 ;
        RECT 63.360 113.400 63.530 113.570 ;
        RECT 63.720 113.400 63.890 113.570 ;
        RECT 64.560 113.400 64.730 113.570 ;
        RECT 64.920 113.400 65.090 113.570 ;
        RECT 65.280 113.400 65.450 113.570 ;
        RECT 66.200 113.400 66.370 113.570 ;
        RECT 66.560 113.400 66.730 113.570 ;
        RECT 66.920 113.400 67.090 113.570 ;
        RECT 68.390 113.450 68.560 113.620 ;
        RECT 68.830 113.450 69.000 113.620 ;
        RECT 69.240 113.450 69.410 113.620 ;
        RECT 69.670 113.450 69.840 113.620 ;
        RECT 70.110 113.450 70.280 113.620 ;
        RECT 70.520 113.450 70.690 113.620 ;
        RECT 72.740 113.400 72.910 113.570 ;
        RECT 73.100 113.400 73.270 113.570 ;
        RECT 74.900 113.450 75.070 113.620 ;
        RECT 75.260 113.450 75.430 113.620 ;
        RECT 75.700 113.450 75.870 113.620 ;
        RECT 77.400 113.400 77.570 113.570 ;
        RECT 77.760 113.400 77.930 113.570 ;
        RECT 78.120 113.400 78.290 113.570 ;
        RECT 79.530 113.400 79.700 113.570 ;
        RECT 79.890 113.400 80.060 113.570 ;
        RECT 80.250 113.400 80.420 113.570 ;
        RECT 81.140 113.450 81.310 113.620 ;
        RECT 81.500 113.450 81.670 113.620 ;
        RECT 81.940 113.450 82.110 113.620 ;
        RECT 83.120 113.400 83.290 113.570 ;
        RECT 83.480 113.400 83.650 113.570 ;
        RECT 83.840 113.400 84.010 113.570 ;
        RECT 84.200 113.400 84.370 113.570 ;
        RECT 84.560 113.400 84.730 113.570 ;
        RECT 84.920 113.400 85.090 113.570 ;
        RECT 85.280 113.400 85.450 113.570 ;
        RECT 85.640 113.400 85.810 113.570 ;
        RECT 86.450 113.400 86.620 113.570 ;
        RECT 86.810 113.400 86.980 113.570 ;
        RECT 87.170 113.400 87.340 113.570 ;
        RECT 87.530 113.400 87.700 113.570 ;
        RECT 88.340 113.450 88.510 113.620 ;
        RECT 88.700 113.450 88.870 113.620 ;
        RECT 89.140 113.450 89.310 113.620 ;
        RECT 90.310 113.400 90.480 113.570 ;
        RECT 90.670 113.400 90.840 113.570 ;
        RECT 91.030 113.400 91.200 113.570 ;
        RECT 92.620 113.400 92.790 113.570 ;
        RECT 92.980 113.400 93.150 113.570 ;
        RECT 93.340 113.400 93.510 113.570 ;
        RECT 94.580 113.450 94.750 113.620 ;
        RECT 94.940 113.450 95.110 113.620 ;
        RECT 95.380 113.450 95.550 113.620 ;
        RECT 96.120 113.400 96.290 113.570 ;
        RECT 96.480 113.400 96.650 113.570 ;
        RECT 96.840 113.400 97.010 113.570 ;
        RECT 97.680 113.400 97.850 113.570 ;
        RECT 98.040 113.400 98.210 113.570 ;
        RECT 98.400 113.400 98.570 113.570 ;
        RECT 99.320 113.400 99.490 113.570 ;
        RECT 99.680 113.400 99.850 113.570 ;
        RECT 100.040 113.400 100.210 113.570 ;
        RECT 101.300 113.450 101.470 113.620 ;
        RECT 101.660 113.450 101.830 113.620 ;
        RECT 102.100 113.450 102.270 113.620 ;
        RECT 102.840 113.400 103.010 113.570 ;
        RECT 103.200 113.400 103.370 113.570 ;
        RECT 103.560 113.400 103.730 113.570 ;
        RECT 104.400 113.400 104.570 113.570 ;
        RECT 104.760 113.400 104.930 113.570 ;
        RECT 105.120 113.400 105.290 113.570 ;
        RECT 106.040 113.400 106.210 113.570 ;
        RECT 106.400 113.400 106.570 113.570 ;
        RECT 106.760 113.400 106.930 113.570 ;
        RECT 108.020 113.450 108.190 113.620 ;
        RECT 108.380 113.450 108.550 113.620 ;
        RECT 108.820 113.450 108.990 113.620 ;
        RECT 110.100 113.400 110.270 113.570 ;
        RECT 110.460 113.400 110.630 113.570 ;
        RECT 112.490 113.400 112.660 113.570 ;
        RECT 114.920 113.400 115.090 113.570 ;
        RECT 115.280 113.400 115.450 113.570 ;
        RECT 115.640 113.400 115.810 113.570 ;
        RECT 117.260 113.400 117.430 113.570 ;
        RECT 117.620 113.400 117.790 113.570 ;
        RECT 117.980 113.400 118.150 113.570 ;
        RECT 119.960 113.400 120.130 113.570 ;
        RECT 120.320 113.400 120.490 113.570 ;
        RECT 120.680 113.400 120.850 113.570 ;
        RECT 121.710 113.400 121.880 113.570 ;
        RECT 122.070 113.400 122.240 113.570 ;
        RECT 122.430 113.400 122.600 113.570 ;
        RECT 123.240 113.400 123.410 113.570 ;
        RECT 123.600 113.400 123.770 113.570 ;
        RECT 123.960 113.400 124.130 113.570 ;
        RECT 125.510 113.450 125.680 113.620 ;
        RECT 125.950 113.450 126.120 113.620 ;
        RECT 126.360 113.450 126.530 113.620 ;
        RECT 126.790 113.450 126.960 113.620 ;
        RECT 127.230 113.450 127.400 113.620 ;
        RECT 127.640 113.450 127.810 113.620 ;
        RECT 129.350 113.450 129.520 113.620 ;
        RECT 129.790 113.450 129.960 113.620 ;
        RECT 130.200 113.450 130.370 113.620 ;
        RECT 130.630 113.450 130.800 113.620 ;
        RECT 131.070 113.450 131.240 113.620 ;
        RECT 131.480 113.450 131.650 113.620 ;
        RECT 133.190 113.450 133.360 113.620 ;
        RECT 133.630 113.450 133.800 113.620 ;
        RECT 134.040 113.450 134.210 113.620 ;
        RECT 134.470 113.450 134.640 113.620 ;
        RECT 134.910 113.450 135.080 113.620 ;
        RECT 135.320 113.450 135.490 113.620 ;
        RECT 137.030 113.450 137.200 113.620 ;
        RECT 137.470 113.450 137.640 113.620 ;
        RECT 137.880 113.450 138.050 113.620 ;
        RECT 138.310 113.450 138.480 113.620 ;
        RECT 138.750 113.450 138.920 113.620 ;
        RECT 139.160 113.450 139.330 113.620 ;
        RECT 140.660 113.450 140.830 113.620 ;
        RECT 141.020 113.450 141.190 113.620 ;
        RECT 141.460 113.450 141.630 113.620 ;
        RECT 6.470 106.160 6.640 106.330 ;
        RECT 6.910 106.160 7.080 106.330 ;
        RECT 7.320 106.160 7.490 106.330 ;
        RECT 7.750 106.160 7.920 106.330 ;
        RECT 8.190 106.160 8.360 106.330 ;
        RECT 8.600 106.160 8.770 106.330 ;
        RECT 10.310 106.160 10.480 106.330 ;
        RECT 10.750 106.160 10.920 106.330 ;
        RECT 11.160 106.160 11.330 106.330 ;
        RECT 11.590 106.160 11.760 106.330 ;
        RECT 12.030 106.160 12.200 106.330 ;
        RECT 12.440 106.160 12.610 106.330 ;
        RECT 14.150 106.160 14.320 106.330 ;
        RECT 14.590 106.160 14.760 106.330 ;
        RECT 15.000 106.160 15.170 106.330 ;
        RECT 15.430 106.160 15.600 106.330 ;
        RECT 15.870 106.160 16.040 106.330 ;
        RECT 16.280 106.160 16.450 106.330 ;
        RECT 17.990 106.160 18.160 106.330 ;
        RECT 18.430 106.160 18.600 106.330 ;
        RECT 18.840 106.160 19.010 106.330 ;
        RECT 19.270 106.160 19.440 106.330 ;
        RECT 19.710 106.160 19.880 106.330 ;
        RECT 20.120 106.160 20.290 106.330 ;
        RECT 21.620 106.160 21.790 106.330 ;
        RECT 21.980 106.160 22.150 106.330 ;
        RECT 22.420 106.160 22.590 106.330 ;
        RECT 23.140 106.210 23.310 106.380 ;
        RECT 23.500 106.210 23.670 106.380 ;
        RECT 23.860 106.210 24.030 106.380 ;
        RECT 24.220 106.210 24.390 106.380 ;
        RECT 25.380 106.210 25.550 106.380 ;
        RECT 25.740 106.210 25.910 106.380 ;
        RECT 26.100 106.210 26.270 106.380 ;
        RECT 26.460 106.210 26.630 106.380 ;
        RECT 27.380 106.160 27.550 106.330 ;
        RECT 27.740 106.160 27.910 106.330 ;
        RECT 28.180 106.160 28.350 106.330 ;
        RECT 29.460 106.210 29.630 106.380 ;
        RECT 29.820 106.210 29.990 106.380 ;
        RECT 31.850 106.210 32.020 106.380 ;
        RECT 34.280 106.210 34.450 106.380 ;
        RECT 34.640 106.210 34.810 106.380 ;
        RECT 35.000 106.210 35.170 106.380 ;
        RECT 36.620 106.210 36.790 106.380 ;
        RECT 36.980 106.210 37.150 106.380 ;
        RECT 37.340 106.210 37.510 106.380 ;
        RECT 39.320 106.210 39.490 106.380 ;
        RECT 39.680 106.210 39.850 106.380 ;
        RECT 40.040 106.210 40.210 106.380 ;
        RECT 41.070 106.210 41.240 106.380 ;
        RECT 41.430 106.210 41.600 106.380 ;
        RECT 41.790 106.210 41.960 106.380 ;
        RECT 42.600 106.210 42.770 106.380 ;
        RECT 42.960 106.210 43.130 106.380 ;
        RECT 43.320 106.210 43.490 106.380 ;
        RECT 44.660 106.160 44.830 106.330 ;
        RECT 45.020 106.160 45.190 106.330 ;
        RECT 45.460 106.160 45.630 106.330 ;
        RECT 46.200 106.210 46.370 106.380 ;
        RECT 46.560 106.210 46.730 106.380 ;
        RECT 48.020 106.160 48.190 106.330 ;
        RECT 48.380 106.160 48.550 106.330 ;
        RECT 48.820 106.160 48.990 106.330 ;
        RECT 50.100 106.210 50.270 106.380 ;
        RECT 50.460 106.210 50.630 106.380 ;
        RECT 52.490 106.210 52.660 106.380 ;
        RECT 54.920 106.210 55.090 106.380 ;
        RECT 55.280 106.210 55.450 106.380 ;
        RECT 55.640 106.210 55.810 106.380 ;
        RECT 57.260 106.210 57.430 106.380 ;
        RECT 57.620 106.210 57.790 106.380 ;
        RECT 57.980 106.210 58.150 106.380 ;
        RECT 59.960 106.210 60.130 106.380 ;
        RECT 60.320 106.210 60.490 106.380 ;
        RECT 60.680 106.210 60.850 106.380 ;
        RECT 61.710 106.210 61.880 106.380 ;
        RECT 62.070 106.210 62.240 106.380 ;
        RECT 62.430 106.210 62.600 106.380 ;
        RECT 63.240 106.210 63.410 106.380 ;
        RECT 63.600 106.210 63.770 106.380 ;
        RECT 63.960 106.210 64.130 106.380 ;
        RECT 65.300 106.160 65.470 106.330 ;
        RECT 65.660 106.160 65.830 106.330 ;
        RECT 66.100 106.160 66.270 106.330 ;
        RECT 66.840 106.210 67.010 106.380 ;
        RECT 67.200 106.210 67.370 106.380 ;
        RECT 67.560 106.210 67.730 106.380 ;
        RECT 68.400 106.210 68.570 106.380 ;
        RECT 68.760 106.210 68.930 106.380 ;
        RECT 69.120 106.210 69.290 106.380 ;
        RECT 70.040 106.210 70.210 106.380 ;
        RECT 70.400 106.210 70.570 106.380 ;
        RECT 70.760 106.210 70.930 106.380 ;
        RECT 72.020 106.160 72.190 106.330 ;
        RECT 72.380 106.160 72.550 106.330 ;
        RECT 72.820 106.160 72.990 106.330 ;
        RECT 74.040 106.210 74.210 106.380 ;
        RECT 74.400 106.210 74.570 106.380 ;
        RECT 74.760 106.210 74.930 106.380 ;
        RECT 75.120 106.210 75.290 106.380 ;
        RECT 75.480 106.210 75.650 106.380 ;
        RECT 76.820 106.160 76.990 106.330 ;
        RECT 77.180 106.160 77.350 106.330 ;
        RECT 77.620 106.160 77.790 106.330 ;
        RECT 78.340 106.210 78.510 106.380 ;
        RECT 78.700 106.210 78.870 106.380 ;
        RECT 79.060 106.210 79.230 106.380 ;
        RECT 79.420 106.210 79.590 106.380 ;
        RECT 80.580 106.210 80.750 106.380 ;
        RECT 80.940 106.210 81.110 106.380 ;
        RECT 81.300 106.210 81.470 106.380 ;
        RECT 81.660 106.210 81.830 106.380 ;
        RECT 82.580 106.160 82.750 106.330 ;
        RECT 82.940 106.160 83.110 106.330 ;
        RECT 83.380 106.160 83.550 106.330 ;
        RECT 84.560 106.210 84.730 106.380 ;
        RECT 84.920 106.210 85.090 106.380 ;
        RECT 85.280 106.210 85.450 106.380 ;
        RECT 85.640 106.210 85.810 106.380 ;
        RECT 86.000 106.210 86.170 106.380 ;
        RECT 86.360 106.210 86.530 106.380 ;
        RECT 86.720 106.210 86.890 106.380 ;
        RECT 87.080 106.210 87.250 106.380 ;
        RECT 87.890 106.210 88.060 106.380 ;
        RECT 88.250 106.210 88.420 106.380 ;
        RECT 88.610 106.210 88.780 106.380 ;
        RECT 88.970 106.210 89.140 106.380 ;
        RECT 89.780 106.160 89.950 106.330 ;
        RECT 90.140 106.160 90.310 106.330 ;
        RECT 90.580 106.160 90.750 106.330 ;
        RECT 92.280 106.210 92.450 106.380 ;
        RECT 92.640 106.210 92.810 106.380 ;
        RECT 93.000 106.210 93.170 106.380 ;
        RECT 93.840 106.210 94.010 106.380 ;
        RECT 94.200 106.210 94.370 106.380 ;
        RECT 94.560 106.210 94.730 106.380 ;
        RECT 95.480 106.210 95.650 106.380 ;
        RECT 95.840 106.210 96.010 106.380 ;
        RECT 96.200 106.210 96.370 106.380 ;
        RECT 97.460 106.160 97.630 106.330 ;
        RECT 97.820 106.160 97.990 106.330 ;
        RECT 98.260 106.160 98.430 106.330 ;
        RECT 99.000 106.210 99.170 106.380 ;
        RECT 99.360 106.210 99.530 106.380 ;
        RECT 99.720 106.210 99.890 106.380 ;
        RECT 100.560 106.210 100.730 106.380 ;
        RECT 100.920 106.210 101.090 106.380 ;
        RECT 101.280 106.210 101.450 106.380 ;
        RECT 102.200 106.210 102.370 106.380 ;
        RECT 102.560 106.210 102.730 106.380 ;
        RECT 102.920 106.210 103.090 106.380 ;
        RECT 104.180 106.160 104.350 106.330 ;
        RECT 104.540 106.160 104.710 106.330 ;
        RECT 104.980 106.160 105.150 106.330 ;
        RECT 105.720 106.210 105.890 106.380 ;
        RECT 106.080 106.210 106.250 106.380 ;
        RECT 106.440 106.210 106.610 106.380 ;
        RECT 107.280 106.210 107.450 106.380 ;
        RECT 107.640 106.210 107.810 106.380 ;
        RECT 108.000 106.210 108.170 106.380 ;
        RECT 108.920 106.210 109.090 106.380 ;
        RECT 109.280 106.210 109.450 106.380 ;
        RECT 109.640 106.210 109.810 106.380 ;
        RECT 110.900 106.160 111.070 106.330 ;
        RECT 111.260 106.160 111.430 106.330 ;
        RECT 111.700 106.160 111.870 106.330 ;
        RECT 113.060 106.210 113.230 106.380 ;
        RECT 113.420 106.210 113.590 106.380 ;
        RECT 115.220 106.160 115.390 106.330 ;
        RECT 115.580 106.160 115.750 106.330 ;
        RECT 116.020 106.160 116.190 106.330 ;
        RECT 117.860 106.210 118.030 106.380 ;
        RECT 118.220 106.210 118.390 106.380 ;
        RECT 120.020 106.160 120.190 106.330 ;
        RECT 120.380 106.160 120.550 106.330 ;
        RECT 120.820 106.160 120.990 106.330 ;
        RECT 121.560 106.210 121.730 106.380 ;
        RECT 121.920 106.210 122.090 106.380 ;
        RECT 122.280 106.210 122.450 106.380 ;
        RECT 123.120 106.210 123.290 106.380 ;
        RECT 123.480 106.210 123.650 106.380 ;
        RECT 123.840 106.210 124.010 106.380 ;
        RECT 124.760 106.210 124.930 106.380 ;
        RECT 125.120 106.210 125.290 106.380 ;
        RECT 125.480 106.210 125.650 106.380 ;
        RECT 126.950 106.160 127.120 106.330 ;
        RECT 127.390 106.160 127.560 106.330 ;
        RECT 127.800 106.160 127.970 106.330 ;
        RECT 128.230 106.160 128.400 106.330 ;
        RECT 128.670 106.160 128.840 106.330 ;
        RECT 129.080 106.160 129.250 106.330 ;
        RECT 130.790 106.160 130.960 106.330 ;
        RECT 131.230 106.160 131.400 106.330 ;
        RECT 131.640 106.160 131.810 106.330 ;
        RECT 132.070 106.160 132.240 106.330 ;
        RECT 132.510 106.160 132.680 106.330 ;
        RECT 132.920 106.160 133.090 106.330 ;
        RECT 134.630 106.160 134.800 106.330 ;
        RECT 135.070 106.160 135.240 106.330 ;
        RECT 135.480 106.160 135.650 106.330 ;
        RECT 135.910 106.160 136.080 106.330 ;
        RECT 136.350 106.160 136.520 106.330 ;
        RECT 136.760 106.160 136.930 106.330 ;
        RECT 138.470 106.160 138.640 106.330 ;
        RECT 138.910 106.160 139.080 106.330 ;
        RECT 139.320 106.160 139.490 106.330 ;
        RECT 139.750 106.160 139.920 106.330 ;
        RECT 140.190 106.160 140.360 106.330 ;
        RECT 140.600 106.160 140.770 106.330 ;
        RECT 5.920 105.730 6.090 105.910 ;
        RECT 6.400 105.730 6.570 105.910 ;
        RECT 6.880 105.730 7.050 105.910 ;
        RECT 7.360 105.730 7.530 105.910 ;
        RECT 7.840 105.730 8.010 105.910 ;
        RECT 8.320 105.730 8.490 105.910 ;
        RECT 8.800 105.730 8.970 105.910 ;
        RECT 9.280 105.730 9.450 105.910 ;
        RECT 9.760 105.730 9.930 105.910 ;
        RECT 10.240 105.730 10.410 105.910 ;
        RECT 10.720 105.730 10.890 105.910 ;
        RECT 11.200 105.730 11.370 105.910 ;
        RECT 11.680 105.730 11.850 105.910 ;
        RECT 12.160 105.730 12.330 105.910 ;
        RECT 12.640 105.730 12.810 105.910 ;
        RECT 13.120 105.730 13.290 105.910 ;
        RECT 13.600 105.730 13.770 105.910 ;
        RECT 14.080 105.730 14.250 105.910 ;
        RECT 14.560 105.730 14.730 105.910 ;
        RECT 15.040 105.730 15.210 105.910 ;
        RECT 15.520 105.730 15.690 105.910 ;
        RECT 16.000 105.730 16.170 105.910 ;
        RECT 16.480 105.730 16.650 105.910 ;
        RECT 16.960 105.730 17.130 105.910 ;
        RECT 17.440 105.730 17.610 105.910 ;
        RECT 17.920 105.730 18.090 105.910 ;
        RECT 18.400 105.730 18.570 105.910 ;
        RECT 18.880 105.730 19.050 105.910 ;
        RECT 19.360 105.730 19.530 105.910 ;
        RECT 19.840 105.730 20.010 105.910 ;
        RECT 20.320 105.730 20.490 105.910 ;
        RECT 20.800 105.730 20.970 105.910 ;
        RECT 21.280 105.730 21.450 105.910 ;
        RECT 21.760 105.730 21.930 105.910 ;
        RECT 22.240 105.730 22.410 105.910 ;
        RECT 22.720 105.730 22.890 105.910 ;
        RECT 23.200 105.730 23.370 105.910 ;
        RECT 23.680 105.730 23.850 105.910 ;
        RECT 24.160 105.730 24.330 105.910 ;
        RECT 24.640 105.730 24.810 105.910 ;
        RECT 25.120 105.730 25.290 105.910 ;
        RECT 25.600 105.730 25.770 105.910 ;
        RECT 26.080 105.730 26.250 105.910 ;
        RECT 26.560 105.730 26.730 105.910 ;
        RECT 27.040 105.730 27.210 105.910 ;
        RECT 27.520 105.730 27.690 105.910 ;
        RECT 28.000 105.730 28.170 105.910 ;
        RECT 28.480 105.730 28.650 105.910 ;
        RECT 28.960 105.730 29.130 105.910 ;
        RECT 29.440 105.730 29.610 105.910 ;
        RECT 29.920 105.730 30.090 105.910 ;
        RECT 30.400 105.730 30.570 105.910 ;
        RECT 30.880 105.730 31.050 105.910 ;
        RECT 31.360 105.730 31.530 105.910 ;
        RECT 31.840 105.730 32.010 105.910 ;
        RECT 32.320 105.730 32.490 105.910 ;
        RECT 32.800 105.730 32.970 105.910 ;
        RECT 33.280 105.730 33.450 105.910 ;
        RECT 33.760 105.730 33.930 105.910 ;
        RECT 34.240 105.730 34.410 105.910 ;
        RECT 34.720 105.730 34.890 105.910 ;
        RECT 35.200 105.730 35.370 105.910 ;
        RECT 35.680 105.730 35.850 105.910 ;
        RECT 36.160 105.730 36.330 105.910 ;
        RECT 36.640 105.730 36.810 105.910 ;
        RECT 37.120 105.730 37.290 105.910 ;
        RECT 37.600 105.730 37.770 105.910 ;
        RECT 38.080 105.730 38.250 105.910 ;
        RECT 38.560 105.730 38.730 105.910 ;
        RECT 39.040 105.730 39.210 105.910 ;
        RECT 39.520 105.730 39.690 105.910 ;
        RECT 40.000 105.730 40.170 105.910 ;
      LAYER li1 ;
        RECT 40.320 105.900 40.800 105.910 ;
      LAYER li1 ;
        RECT 40.480 105.730 40.650 105.900 ;
        RECT 40.960 105.730 41.130 105.910 ;
        RECT 41.440 105.730 41.610 105.910 ;
        RECT 41.920 105.730 42.090 105.910 ;
        RECT 42.400 105.730 42.570 105.910 ;
        RECT 42.880 105.730 43.050 105.910 ;
        RECT 43.360 105.730 43.530 105.910 ;
        RECT 43.840 105.730 44.010 105.910 ;
        RECT 44.320 105.730 44.490 105.910 ;
        RECT 44.800 105.730 44.970 105.910 ;
        RECT 45.280 105.730 45.450 105.910 ;
        RECT 45.760 105.730 45.930 105.910 ;
        RECT 46.240 105.730 46.410 105.910 ;
        RECT 46.720 105.730 46.890 105.910 ;
        RECT 47.200 105.730 47.370 105.910 ;
        RECT 47.680 105.730 47.850 105.910 ;
        RECT 48.160 105.730 48.330 105.910 ;
        RECT 48.640 105.730 48.810 105.910 ;
        RECT 49.120 105.730 49.290 105.910 ;
        RECT 49.600 105.730 49.770 105.910 ;
        RECT 50.080 105.730 50.250 105.910 ;
        RECT 50.560 105.730 50.730 105.910 ;
        RECT 51.040 105.730 51.210 105.910 ;
        RECT 51.520 105.730 51.690 105.910 ;
        RECT 52.000 105.730 52.170 105.910 ;
        RECT 52.480 105.730 52.650 105.910 ;
        RECT 52.960 105.730 53.130 105.910 ;
        RECT 53.440 105.730 53.610 105.910 ;
        RECT 53.920 105.730 54.090 105.910 ;
        RECT 54.400 105.730 54.570 105.910 ;
        RECT 54.880 105.730 55.050 105.910 ;
        RECT 55.360 105.730 55.530 105.910 ;
        RECT 55.840 105.730 56.010 105.910 ;
        RECT 56.320 105.730 56.490 105.910 ;
        RECT 56.800 105.730 56.970 105.910 ;
        RECT 57.280 105.730 57.450 105.910 ;
        RECT 57.760 105.730 57.930 105.910 ;
        RECT 58.240 105.730 58.410 105.910 ;
        RECT 58.720 105.730 58.890 105.910 ;
        RECT 59.200 105.730 59.370 105.910 ;
        RECT 59.680 105.730 59.850 105.910 ;
        RECT 60.160 105.730 60.330 105.910 ;
        RECT 60.640 105.730 60.810 105.910 ;
      LAYER li1 ;
        RECT 60.960 105.900 61.440 105.910 ;
      LAYER li1 ;
        RECT 61.120 105.730 61.290 105.900 ;
        RECT 61.600 105.730 61.770 105.910 ;
        RECT 62.080 105.730 62.250 105.910 ;
        RECT 62.560 105.730 62.730 105.910 ;
        RECT 63.040 105.730 63.210 105.910 ;
        RECT 63.520 105.730 63.690 105.910 ;
        RECT 64.000 105.730 64.170 105.910 ;
        RECT 64.480 105.730 64.650 105.910 ;
        RECT 64.960 105.730 65.130 105.910 ;
        RECT 65.440 105.730 65.610 105.910 ;
        RECT 65.920 105.730 66.090 105.910 ;
        RECT 66.400 105.730 66.570 105.910 ;
        RECT 66.880 105.730 67.050 105.910 ;
        RECT 67.360 105.730 67.530 105.910 ;
        RECT 67.840 105.730 68.010 105.910 ;
        RECT 68.320 105.730 68.490 105.910 ;
        RECT 68.800 105.730 68.970 105.910 ;
        RECT 69.280 105.730 69.450 105.910 ;
        RECT 69.760 105.730 69.930 105.910 ;
        RECT 70.240 105.730 70.410 105.910 ;
        RECT 70.720 105.730 70.890 105.910 ;
        RECT 71.200 105.730 71.370 105.910 ;
        RECT 71.680 105.730 71.850 105.910 ;
        RECT 72.160 105.730 72.330 105.910 ;
        RECT 72.640 105.730 72.810 105.910 ;
        RECT 73.120 105.730 73.290 105.910 ;
        RECT 73.600 105.900 73.770 105.910 ;
      LAYER li1 ;
        RECT 73.440 105.730 73.920 105.900 ;
      LAYER li1 ;
        RECT 74.080 105.730 74.250 105.910 ;
        RECT 74.560 105.730 74.730 105.910 ;
        RECT 75.040 105.730 75.210 105.910 ;
        RECT 75.520 105.730 75.690 105.910 ;
        RECT 76.000 105.730 76.170 105.910 ;
        RECT 76.480 105.730 76.650 105.910 ;
        RECT 76.960 105.730 77.130 105.910 ;
        RECT 77.440 105.730 77.610 105.910 ;
        RECT 77.920 105.730 78.090 105.910 ;
        RECT 78.400 105.730 78.570 105.910 ;
        RECT 78.880 105.730 79.050 105.910 ;
        RECT 79.360 105.730 79.530 105.910 ;
        RECT 79.840 105.730 80.010 105.910 ;
        RECT 80.320 105.730 80.490 105.910 ;
        RECT 80.800 105.730 80.970 105.910 ;
        RECT 81.280 105.730 81.450 105.910 ;
        RECT 81.760 105.730 81.930 105.910 ;
        RECT 82.240 105.730 82.410 105.910 ;
        RECT 82.720 105.730 82.890 105.910 ;
        RECT 83.200 105.730 83.370 105.910 ;
        RECT 83.680 105.730 83.850 105.910 ;
        RECT 84.160 105.730 84.330 105.910 ;
        RECT 84.640 105.730 84.810 105.910 ;
        RECT 85.120 105.730 85.290 105.910 ;
        RECT 85.600 105.730 85.770 105.910 ;
        RECT 86.080 105.730 86.250 105.910 ;
        RECT 86.560 105.730 86.730 105.910 ;
        RECT 87.040 105.730 87.210 105.910 ;
        RECT 87.520 105.730 87.690 105.910 ;
        RECT 88.000 105.730 88.170 105.910 ;
        RECT 88.480 105.730 88.650 105.910 ;
        RECT 88.960 105.730 89.130 105.910 ;
        RECT 89.440 105.730 89.610 105.910 ;
        RECT 89.920 105.730 90.090 105.910 ;
        RECT 90.400 105.730 90.570 105.910 ;
        RECT 90.880 105.730 91.050 105.910 ;
        RECT 91.360 105.730 91.530 105.910 ;
        RECT 91.840 105.730 92.010 105.910 ;
        RECT 92.320 105.730 92.490 105.910 ;
        RECT 92.800 105.730 92.970 105.910 ;
        RECT 93.280 105.730 93.450 105.910 ;
        RECT 93.760 105.730 93.930 105.910 ;
        RECT 94.240 105.730 94.410 105.910 ;
        RECT 94.720 105.730 94.890 105.910 ;
        RECT 95.200 105.730 95.370 105.910 ;
        RECT 95.680 105.730 95.850 105.910 ;
        RECT 96.160 105.730 96.330 105.910 ;
        RECT 96.640 105.730 96.810 105.910 ;
        RECT 97.120 105.730 97.290 105.910 ;
        RECT 97.600 105.730 97.770 105.910 ;
        RECT 98.080 105.730 98.250 105.910 ;
        RECT 98.560 105.730 98.730 105.910 ;
        RECT 99.040 105.730 99.210 105.910 ;
        RECT 99.520 105.730 99.690 105.910 ;
        RECT 100.000 105.730 100.170 105.910 ;
        RECT 100.480 105.730 100.650 105.910 ;
        RECT 100.960 105.730 101.130 105.910 ;
        RECT 101.440 105.730 101.610 105.910 ;
        RECT 101.920 105.730 102.090 105.910 ;
        RECT 102.400 105.730 102.570 105.910 ;
        RECT 102.880 105.730 103.050 105.910 ;
        RECT 103.360 105.730 103.530 105.910 ;
        RECT 103.840 105.730 104.010 105.910 ;
        RECT 104.320 105.730 104.490 105.910 ;
        RECT 104.800 105.730 104.970 105.910 ;
        RECT 105.280 105.730 105.450 105.910 ;
        RECT 105.760 105.730 105.930 105.910 ;
        RECT 106.240 105.730 106.410 105.910 ;
        RECT 106.720 105.730 106.890 105.910 ;
        RECT 107.200 105.730 107.370 105.910 ;
        RECT 107.680 105.730 107.850 105.910 ;
        RECT 108.160 105.730 108.330 105.910 ;
        RECT 108.640 105.730 108.810 105.910 ;
        RECT 109.120 105.730 109.290 105.910 ;
        RECT 109.600 105.730 109.770 105.910 ;
        RECT 110.080 105.730 110.250 105.910 ;
        RECT 110.560 105.730 110.730 105.910 ;
        RECT 111.040 105.730 111.210 105.910 ;
        RECT 111.520 105.730 111.690 105.910 ;
        RECT 112.000 105.730 112.170 105.910 ;
        RECT 112.480 105.730 112.650 105.910 ;
        RECT 112.960 105.730 113.130 105.910 ;
        RECT 113.440 105.730 113.610 105.910 ;
        RECT 113.920 105.730 114.090 105.910 ;
        RECT 114.400 105.730 114.570 105.910 ;
        RECT 114.880 105.730 115.050 105.910 ;
        RECT 115.360 105.730 115.530 105.910 ;
        RECT 115.840 105.730 116.010 105.910 ;
        RECT 116.320 105.730 116.490 105.910 ;
        RECT 116.800 105.900 116.970 105.910 ;
      LAYER li1 ;
        RECT 116.640 105.730 117.120 105.900 ;
      LAYER li1 ;
        RECT 117.280 105.730 117.450 105.910 ;
        RECT 117.760 105.730 117.930 105.910 ;
        RECT 118.240 105.730 118.410 105.910 ;
        RECT 118.720 105.730 118.890 105.910 ;
        RECT 119.200 105.730 119.370 105.910 ;
        RECT 119.680 105.730 119.850 105.910 ;
        RECT 120.160 105.730 120.330 105.910 ;
        RECT 120.640 105.730 120.810 105.910 ;
      LAYER li1 ;
        RECT 120.960 105.900 121.440 105.910 ;
      LAYER li1 ;
        RECT 121.120 105.730 121.290 105.900 ;
        RECT 121.600 105.730 121.770 105.910 ;
        RECT 122.080 105.730 122.250 105.910 ;
        RECT 122.560 105.730 122.730 105.910 ;
        RECT 123.040 105.730 123.210 105.910 ;
        RECT 123.520 105.730 123.690 105.910 ;
        RECT 124.000 105.730 124.170 105.910 ;
        RECT 124.480 105.730 124.650 105.910 ;
        RECT 124.960 105.730 125.130 105.910 ;
        RECT 125.440 105.730 125.610 105.910 ;
        RECT 125.920 105.730 126.090 105.910 ;
        RECT 126.400 105.730 126.570 105.910 ;
        RECT 126.880 105.730 127.050 105.910 ;
        RECT 127.360 105.730 127.530 105.910 ;
        RECT 127.840 105.730 128.010 105.910 ;
        RECT 128.320 105.730 128.490 105.910 ;
        RECT 128.800 105.730 128.970 105.910 ;
        RECT 129.280 105.730 129.450 105.910 ;
        RECT 129.760 105.730 129.930 105.910 ;
        RECT 130.240 105.730 130.410 105.910 ;
        RECT 130.720 105.730 130.890 105.910 ;
        RECT 131.200 105.730 131.370 105.910 ;
        RECT 131.680 105.730 131.850 105.910 ;
        RECT 132.160 105.730 132.330 105.910 ;
        RECT 132.640 105.730 132.810 105.910 ;
        RECT 133.120 105.730 133.290 105.910 ;
        RECT 133.600 105.730 133.770 105.910 ;
        RECT 134.080 105.730 134.250 105.910 ;
        RECT 134.560 105.730 134.730 105.910 ;
        RECT 135.040 105.730 135.210 105.910 ;
        RECT 135.520 105.730 135.690 105.910 ;
        RECT 136.000 105.730 136.170 105.910 ;
        RECT 136.480 105.730 136.650 105.910 ;
        RECT 136.960 105.730 137.130 105.910 ;
        RECT 137.440 105.730 137.610 105.910 ;
        RECT 137.920 105.730 138.090 105.910 ;
        RECT 138.400 105.730 138.570 105.910 ;
        RECT 138.880 105.730 139.050 105.910 ;
        RECT 139.360 105.730 139.530 105.910 ;
        RECT 139.840 105.730 140.010 105.910 ;
        RECT 140.320 105.730 140.490 105.910 ;
        RECT 140.800 105.730 140.970 105.910 ;
        RECT 141.280 105.730 141.450 105.910 ;
        RECT 141.760 105.900 141.930 105.910 ;
      LAYER li1 ;
        RECT 141.600 105.730 142.080 105.900 ;
      LAYER li1 ;
        RECT 6.470 105.310 6.640 105.480 ;
        RECT 6.910 105.310 7.080 105.480 ;
        RECT 7.320 105.310 7.490 105.480 ;
        RECT 7.750 105.310 7.920 105.480 ;
        RECT 8.190 105.310 8.360 105.480 ;
        RECT 8.600 105.310 8.770 105.480 ;
        RECT 10.260 105.260 10.430 105.430 ;
        RECT 10.620 105.260 10.790 105.430 ;
        RECT 12.650 105.260 12.820 105.430 ;
        RECT 15.080 105.260 15.250 105.430 ;
        RECT 15.440 105.260 15.610 105.430 ;
        RECT 15.800 105.260 15.970 105.430 ;
        RECT 17.420 105.260 17.590 105.430 ;
        RECT 17.780 105.260 17.950 105.430 ;
        RECT 18.140 105.260 18.310 105.430 ;
        RECT 20.120 105.260 20.290 105.430 ;
        RECT 20.480 105.260 20.650 105.430 ;
        RECT 20.840 105.260 21.010 105.430 ;
        RECT 21.870 105.260 22.040 105.430 ;
        RECT 22.230 105.260 22.400 105.430 ;
        RECT 22.590 105.260 22.760 105.430 ;
        RECT 23.400 105.260 23.570 105.430 ;
        RECT 23.760 105.260 23.930 105.430 ;
        RECT 24.120 105.260 24.290 105.430 ;
        RECT 25.460 105.310 25.630 105.480 ;
        RECT 25.820 105.310 25.990 105.480 ;
        RECT 26.260 105.310 26.430 105.480 ;
        RECT 27.000 105.260 27.170 105.430 ;
        RECT 27.360 105.260 27.530 105.430 ;
        RECT 28.820 105.310 28.990 105.480 ;
        RECT 29.180 105.310 29.350 105.480 ;
        RECT 29.620 105.310 29.790 105.480 ;
        RECT 31.770 105.260 31.940 105.430 ;
        RECT 32.130 105.260 32.300 105.430 ;
        RECT 32.490 105.260 32.660 105.430 ;
        RECT 34.940 105.260 35.110 105.430 ;
        RECT 35.300 105.260 35.470 105.430 ;
        RECT 35.660 105.260 35.830 105.430 ;
        RECT 37.190 105.310 37.360 105.480 ;
        RECT 37.630 105.310 37.800 105.480 ;
        RECT 38.040 105.310 38.210 105.480 ;
        RECT 38.470 105.310 38.640 105.480 ;
        RECT 38.910 105.310 39.080 105.480 ;
        RECT 39.320 105.310 39.490 105.480 ;
        RECT 40.920 105.260 41.090 105.430 ;
        RECT 41.280 105.260 41.450 105.430 ;
        RECT 41.640 105.260 41.810 105.430 ;
        RECT 42.480 105.260 42.650 105.430 ;
        RECT 42.840 105.260 43.010 105.430 ;
        RECT 43.200 105.260 43.370 105.430 ;
        RECT 44.120 105.260 44.290 105.430 ;
        RECT 44.480 105.260 44.650 105.430 ;
        RECT 44.840 105.260 45.010 105.430 ;
        RECT 46.100 105.310 46.270 105.480 ;
        RECT 46.460 105.310 46.630 105.480 ;
        RECT 46.900 105.310 47.070 105.480 ;
        RECT 47.640 105.260 47.810 105.430 ;
        RECT 48.000 105.260 48.170 105.430 ;
        RECT 48.360 105.260 48.530 105.430 ;
        RECT 49.200 105.260 49.370 105.430 ;
        RECT 49.560 105.260 49.730 105.430 ;
        RECT 49.920 105.260 50.090 105.430 ;
        RECT 50.840 105.260 51.010 105.430 ;
        RECT 51.200 105.260 51.370 105.430 ;
        RECT 51.560 105.260 51.730 105.430 ;
        RECT 52.820 105.310 52.990 105.480 ;
        RECT 53.180 105.310 53.350 105.480 ;
        RECT 53.620 105.310 53.790 105.480 ;
        RECT 54.360 105.260 54.530 105.430 ;
        RECT 54.720 105.260 54.890 105.430 ;
        RECT 55.080 105.260 55.250 105.430 ;
        RECT 55.920 105.260 56.090 105.430 ;
        RECT 56.280 105.260 56.450 105.430 ;
        RECT 56.640 105.260 56.810 105.430 ;
        RECT 57.560 105.260 57.730 105.430 ;
        RECT 57.920 105.260 58.090 105.430 ;
        RECT 58.280 105.260 58.450 105.430 ;
        RECT 59.540 105.310 59.710 105.480 ;
        RECT 59.900 105.310 60.070 105.480 ;
        RECT 60.340 105.310 60.510 105.480 ;
        RECT 61.560 105.260 61.730 105.430 ;
        RECT 61.920 105.260 62.090 105.430 ;
        RECT 63.380 105.310 63.550 105.480 ;
        RECT 63.740 105.310 63.910 105.480 ;
        RECT 64.180 105.310 64.350 105.480 ;
        RECT 65.460 105.260 65.630 105.430 ;
        RECT 65.820 105.260 65.990 105.430 ;
        RECT 67.850 105.260 68.020 105.430 ;
        RECT 70.280 105.260 70.450 105.430 ;
        RECT 70.640 105.260 70.810 105.430 ;
        RECT 71.000 105.260 71.170 105.430 ;
        RECT 72.620 105.260 72.790 105.430 ;
        RECT 72.980 105.260 73.150 105.430 ;
        RECT 73.340 105.260 73.510 105.430 ;
        RECT 75.320 105.260 75.490 105.430 ;
        RECT 75.680 105.260 75.850 105.430 ;
        RECT 76.040 105.260 76.210 105.430 ;
        RECT 77.070 105.260 77.240 105.430 ;
        RECT 77.430 105.260 77.600 105.430 ;
        RECT 77.790 105.260 77.960 105.430 ;
        RECT 78.600 105.260 78.770 105.430 ;
        RECT 78.960 105.260 79.130 105.430 ;
        RECT 79.320 105.260 79.490 105.430 ;
        RECT 80.660 105.310 80.830 105.480 ;
        RECT 81.020 105.310 81.190 105.480 ;
        RECT 81.460 105.310 81.630 105.480 ;
        RECT 82.200 105.260 82.370 105.430 ;
        RECT 82.560 105.260 82.730 105.430 ;
        RECT 82.920 105.260 83.090 105.430 ;
        RECT 83.760 105.260 83.930 105.430 ;
        RECT 84.120 105.260 84.290 105.430 ;
        RECT 84.480 105.260 84.650 105.430 ;
        RECT 85.400 105.260 85.570 105.430 ;
        RECT 85.760 105.260 85.930 105.430 ;
        RECT 86.120 105.260 86.290 105.430 ;
        RECT 87.380 105.310 87.550 105.480 ;
        RECT 87.740 105.310 87.910 105.480 ;
        RECT 88.180 105.310 88.350 105.480 ;
        RECT 88.920 105.260 89.090 105.430 ;
        RECT 89.280 105.260 89.450 105.430 ;
        RECT 89.640 105.260 89.810 105.430 ;
        RECT 90.480 105.260 90.650 105.430 ;
        RECT 90.840 105.260 91.010 105.430 ;
        RECT 91.200 105.260 91.370 105.430 ;
        RECT 92.120 105.260 92.290 105.430 ;
        RECT 92.480 105.260 92.650 105.430 ;
        RECT 92.840 105.260 93.010 105.430 ;
        RECT 94.310 105.310 94.480 105.480 ;
        RECT 94.750 105.310 94.920 105.480 ;
        RECT 95.160 105.310 95.330 105.480 ;
        RECT 95.590 105.310 95.760 105.480 ;
        RECT 96.030 105.310 96.200 105.480 ;
        RECT 96.440 105.310 96.610 105.480 ;
        RECT 98.960 105.260 99.130 105.430 ;
        RECT 99.320 105.260 99.490 105.430 ;
        RECT 99.680 105.260 99.850 105.430 ;
        RECT 100.040 105.260 100.210 105.430 ;
        RECT 100.400 105.260 100.570 105.430 ;
        RECT 100.760 105.260 100.930 105.430 ;
        RECT 101.120 105.260 101.290 105.430 ;
        RECT 101.480 105.260 101.650 105.430 ;
        RECT 102.290 105.260 102.460 105.430 ;
        RECT 102.650 105.260 102.820 105.430 ;
        RECT 103.010 105.260 103.180 105.430 ;
        RECT 103.370 105.260 103.540 105.430 ;
        RECT 104.180 105.310 104.350 105.480 ;
        RECT 104.540 105.310 104.710 105.480 ;
        RECT 104.980 105.310 105.150 105.480 ;
        RECT 105.720 105.260 105.890 105.430 ;
        RECT 106.080 105.260 106.250 105.430 ;
        RECT 106.440 105.260 106.610 105.430 ;
        RECT 107.280 105.260 107.450 105.430 ;
        RECT 107.640 105.260 107.810 105.430 ;
        RECT 108.000 105.260 108.170 105.430 ;
        RECT 108.920 105.260 109.090 105.430 ;
        RECT 109.280 105.260 109.450 105.430 ;
        RECT 109.640 105.260 109.810 105.430 ;
        RECT 110.900 105.310 111.070 105.480 ;
        RECT 111.260 105.310 111.430 105.480 ;
        RECT 111.700 105.310 111.870 105.480 ;
        RECT 112.440 105.260 112.610 105.430 ;
        RECT 112.800 105.260 112.970 105.430 ;
        RECT 113.160 105.260 113.330 105.430 ;
        RECT 114.000 105.260 114.170 105.430 ;
        RECT 114.360 105.260 114.530 105.430 ;
        RECT 114.720 105.260 114.890 105.430 ;
        RECT 115.640 105.260 115.810 105.430 ;
        RECT 116.000 105.260 116.170 105.430 ;
        RECT 116.360 105.260 116.530 105.430 ;
        RECT 117.830 105.310 118.000 105.480 ;
        RECT 118.270 105.310 118.440 105.480 ;
        RECT 118.680 105.310 118.850 105.480 ;
        RECT 119.110 105.310 119.280 105.480 ;
        RECT 119.550 105.310 119.720 105.480 ;
        RECT 119.960 105.310 120.130 105.480 ;
        RECT 121.560 105.260 121.730 105.430 ;
        RECT 121.920 105.260 122.090 105.430 ;
        RECT 122.280 105.260 122.450 105.430 ;
        RECT 123.120 105.260 123.290 105.430 ;
        RECT 123.480 105.260 123.650 105.430 ;
        RECT 123.840 105.260 124.010 105.430 ;
        RECT 124.760 105.260 124.930 105.430 ;
        RECT 125.120 105.260 125.290 105.430 ;
        RECT 125.480 105.260 125.650 105.430 ;
        RECT 126.950 105.310 127.120 105.480 ;
        RECT 127.390 105.310 127.560 105.480 ;
        RECT 127.800 105.310 127.970 105.480 ;
        RECT 128.230 105.310 128.400 105.480 ;
        RECT 128.670 105.310 128.840 105.480 ;
        RECT 129.080 105.310 129.250 105.480 ;
        RECT 130.790 105.310 130.960 105.480 ;
        RECT 131.230 105.310 131.400 105.480 ;
        RECT 131.640 105.310 131.810 105.480 ;
        RECT 132.070 105.310 132.240 105.480 ;
        RECT 132.510 105.310 132.680 105.480 ;
        RECT 132.920 105.310 133.090 105.480 ;
        RECT 135.000 105.260 135.170 105.430 ;
        RECT 135.360 105.260 135.530 105.430 ;
        RECT 137.030 105.310 137.200 105.480 ;
        RECT 137.470 105.310 137.640 105.480 ;
        RECT 137.880 105.310 138.050 105.480 ;
        RECT 138.310 105.310 138.480 105.480 ;
        RECT 138.750 105.310 138.920 105.480 ;
        RECT 139.160 105.310 139.330 105.480 ;
        RECT 140.660 105.310 140.830 105.480 ;
        RECT 141.020 105.310 141.190 105.480 ;
        RECT 141.460 105.310 141.630 105.480 ;
        RECT 6.470 98.020 6.640 98.190 ;
        RECT 6.910 98.020 7.080 98.190 ;
        RECT 7.320 98.020 7.490 98.190 ;
        RECT 7.750 98.020 7.920 98.190 ;
        RECT 8.190 98.020 8.360 98.190 ;
        RECT 8.600 98.020 8.770 98.190 ;
        RECT 10.310 98.020 10.480 98.190 ;
        RECT 10.750 98.020 10.920 98.190 ;
        RECT 11.160 98.020 11.330 98.190 ;
        RECT 11.590 98.020 11.760 98.190 ;
        RECT 12.030 98.020 12.200 98.190 ;
        RECT 12.440 98.020 12.610 98.190 ;
        RECT 13.940 98.020 14.110 98.190 ;
        RECT 14.300 98.020 14.470 98.190 ;
        RECT 14.740 98.020 14.910 98.190 ;
        RECT 17.060 98.070 17.230 98.240 ;
        RECT 17.420 98.070 17.590 98.240 ;
        RECT 19.220 98.020 19.390 98.190 ;
        RECT 19.580 98.020 19.750 98.190 ;
        RECT 20.020 98.020 20.190 98.190 ;
        RECT 22.200 98.070 22.370 98.240 ;
        RECT 22.560 98.070 22.730 98.240 ;
        RECT 24.230 98.020 24.400 98.190 ;
        RECT 24.670 98.020 24.840 98.190 ;
        RECT 25.080 98.020 25.250 98.190 ;
        RECT 25.510 98.020 25.680 98.190 ;
        RECT 25.950 98.020 26.120 98.190 ;
        RECT 26.360 98.020 26.530 98.190 ;
        RECT 28.920 98.070 29.090 98.240 ;
        RECT 29.280 98.070 29.450 98.240 ;
        RECT 30.740 98.020 30.910 98.190 ;
        RECT 31.100 98.020 31.270 98.190 ;
        RECT 31.540 98.020 31.710 98.190 ;
        RECT 32.900 98.070 33.070 98.240 ;
        RECT 33.260 98.070 33.430 98.240 ;
        RECT 35.060 98.020 35.230 98.190 ;
        RECT 35.420 98.020 35.590 98.190 ;
        RECT 35.860 98.020 36.030 98.190 ;
        RECT 37.220 98.070 37.390 98.240 ;
        RECT 37.580 98.070 37.750 98.240 ;
        RECT 39.380 98.020 39.550 98.190 ;
        RECT 39.740 98.020 39.910 98.190 ;
        RECT 40.180 98.020 40.350 98.190 ;
        RECT 40.920 98.070 41.090 98.240 ;
        RECT 41.280 98.070 41.450 98.240 ;
        RECT 41.640 98.070 41.810 98.240 ;
        RECT 42.480 98.070 42.650 98.240 ;
        RECT 42.840 98.070 43.010 98.240 ;
        RECT 43.200 98.070 43.370 98.240 ;
        RECT 44.120 98.070 44.290 98.240 ;
        RECT 44.480 98.070 44.650 98.240 ;
        RECT 44.840 98.070 45.010 98.240 ;
        RECT 46.100 98.020 46.270 98.190 ;
        RECT 46.460 98.020 46.630 98.190 ;
        RECT 46.900 98.020 47.070 98.190 ;
        RECT 47.640 98.070 47.810 98.240 ;
        RECT 48.000 98.070 48.170 98.240 ;
        RECT 48.360 98.070 48.530 98.240 ;
        RECT 49.200 98.070 49.370 98.240 ;
        RECT 49.560 98.070 49.730 98.240 ;
        RECT 49.920 98.070 50.090 98.240 ;
        RECT 50.840 98.070 51.010 98.240 ;
        RECT 51.200 98.070 51.370 98.240 ;
        RECT 51.560 98.070 51.730 98.240 ;
        RECT 52.820 98.020 52.990 98.190 ;
        RECT 53.180 98.020 53.350 98.190 ;
        RECT 53.620 98.020 53.790 98.190 ;
        RECT 54.360 98.070 54.530 98.240 ;
        RECT 54.720 98.070 54.890 98.240 ;
        RECT 55.080 98.070 55.250 98.240 ;
        RECT 55.920 98.070 56.090 98.240 ;
        RECT 56.280 98.070 56.450 98.240 ;
        RECT 56.640 98.070 56.810 98.240 ;
        RECT 57.560 98.070 57.730 98.240 ;
        RECT 57.920 98.070 58.090 98.240 ;
        RECT 58.280 98.070 58.450 98.240 ;
        RECT 59.540 98.020 59.710 98.190 ;
        RECT 59.900 98.020 60.070 98.190 ;
        RECT 60.340 98.020 60.510 98.190 ;
        RECT 61.060 98.070 61.230 98.240 ;
        RECT 61.420 98.070 61.590 98.240 ;
        RECT 61.780 98.070 61.950 98.240 ;
        RECT 62.140 98.070 62.310 98.240 ;
        RECT 63.300 98.070 63.470 98.240 ;
        RECT 63.660 98.070 63.830 98.240 ;
        RECT 64.020 98.070 64.190 98.240 ;
        RECT 64.380 98.070 64.550 98.240 ;
        RECT 65.300 98.020 65.470 98.190 ;
        RECT 65.660 98.020 65.830 98.190 ;
        RECT 66.100 98.020 66.270 98.190 ;
        RECT 67.460 98.070 67.630 98.240 ;
        RECT 67.820 98.070 67.990 98.240 ;
        RECT 69.620 98.020 69.790 98.190 ;
        RECT 69.980 98.020 70.150 98.190 ;
        RECT 70.420 98.020 70.590 98.190 ;
        RECT 72.600 98.070 72.770 98.240 ;
        RECT 72.960 98.070 73.130 98.240 ;
        RECT 73.320 98.070 73.490 98.240 ;
        RECT 73.680 98.070 73.850 98.240 ;
        RECT 74.040 98.070 74.210 98.240 ;
        RECT 76.340 98.020 76.510 98.190 ;
        RECT 76.700 98.020 76.870 98.190 ;
        RECT 77.140 98.020 77.310 98.190 ;
        RECT 77.880 98.070 78.050 98.240 ;
        RECT 78.240 98.070 78.410 98.240 ;
        RECT 78.600 98.070 78.770 98.240 ;
        RECT 79.440 98.070 79.610 98.240 ;
        RECT 79.800 98.070 79.970 98.240 ;
        RECT 80.160 98.070 80.330 98.240 ;
        RECT 81.080 98.070 81.250 98.240 ;
        RECT 81.440 98.070 81.610 98.240 ;
        RECT 81.800 98.070 81.970 98.240 ;
        RECT 83.060 98.020 83.230 98.190 ;
        RECT 83.420 98.020 83.590 98.190 ;
        RECT 83.860 98.020 84.030 98.190 ;
        RECT 84.600 98.070 84.770 98.240 ;
        RECT 84.960 98.070 85.130 98.240 ;
        RECT 85.320 98.070 85.490 98.240 ;
        RECT 86.160 98.070 86.330 98.240 ;
        RECT 86.520 98.070 86.690 98.240 ;
        RECT 86.880 98.070 87.050 98.240 ;
        RECT 87.800 98.070 87.970 98.240 ;
        RECT 88.160 98.070 88.330 98.240 ;
        RECT 88.520 98.070 88.690 98.240 ;
        RECT 89.990 98.020 90.160 98.190 ;
        RECT 90.430 98.020 90.600 98.190 ;
        RECT 90.840 98.020 91.010 98.190 ;
        RECT 91.270 98.020 91.440 98.190 ;
        RECT 91.710 98.020 91.880 98.190 ;
        RECT 92.120 98.020 92.290 98.190 ;
        RECT 93.240 98.070 93.410 98.240 ;
        RECT 93.600 98.070 93.770 98.240 ;
        RECT 93.960 98.070 94.130 98.240 ;
        RECT 94.800 98.070 94.970 98.240 ;
        RECT 95.160 98.070 95.330 98.240 ;
        RECT 95.520 98.070 95.690 98.240 ;
        RECT 96.440 98.070 96.610 98.240 ;
        RECT 96.800 98.070 96.970 98.240 ;
        RECT 97.160 98.070 97.330 98.240 ;
        RECT 98.420 98.020 98.590 98.190 ;
        RECT 98.780 98.020 98.950 98.190 ;
        RECT 99.220 98.020 99.390 98.190 ;
        RECT 100.400 98.070 100.570 98.240 ;
        RECT 100.760 98.070 100.930 98.240 ;
        RECT 101.120 98.070 101.290 98.240 ;
        RECT 101.480 98.070 101.650 98.240 ;
        RECT 101.840 98.070 102.010 98.240 ;
        RECT 102.200 98.070 102.370 98.240 ;
        RECT 102.560 98.070 102.730 98.240 ;
        RECT 102.920 98.070 103.090 98.240 ;
        RECT 103.730 98.070 103.900 98.240 ;
        RECT 104.090 98.070 104.260 98.240 ;
        RECT 104.450 98.070 104.620 98.240 ;
        RECT 104.810 98.070 104.980 98.240 ;
        RECT 105.620 98.020 105.790 98.190 ;
        RECT 105.980 98.020 106.150 98.190 ;
        RECT 106.420 98.020 106.590 98.190 ;
        RECT 107.780 98.070 107.950 98.240 ;
        RECT 108.140 98.070 108.310 98.240 ;
        RECT 109.940 98.020 110.110 98.190 ;
        RECT 110.300 98.020 110.470 98.190 ;
        RECT 110.740 98.020 110.910 98.190 ;
        RECT 111.940 98.070 112.110 98.240 ;
        RECT 112.300 98.070 112.470 98.240 ;
        RECT 112.660 98.070 112.830 98.240 ;
        RECT 113.630 98.070 113.800 98.240 ;
        RECT 117.000 98.070 117.170 98.240 ;
        RECT 118.470 98.070 118.640 98.240 ;
        RECT 118.830 98.070 119.000 98.240 ;
        RECT 119.190 98.070 119.360 98.240 ;
        RECT 121.400 98.070 121.570 98.240 ;
        RECT 121.760 98.070 121.930 98.240 ;
        RECT 122.120 98.070 122.290 98.240 ;
        RECT 123.120 98.070 123.290 98.240 ;
        RECT 123.480 98.070 123.650 98.240 ;
        RECT 123.840 98.070 124.010 98.240 ;
        RECT 124.680 98.070 124.850 98.240 ;
        RECT 125.040 98.070 125.210 98.240 ;
        RECT 125.400 98.070 125.570 98.240 ;
        RECT 126.740 98.020 126.910 98.190 ;
        RECT 127.100 98.020 127.270 98.190 ;
        RECT 127.540 98.020 127.710 98.190 ;
        RECT 128.280 98.070 128.450 98.240 ;
        RECT 128.640 98.070 128.810 98.240 ;
        RECT 129.000 98.070 129.170 98.240 ;
        RECT 129.840 98.070 130.010 98.240 ;
        RECT 130.200 98.070 130.370 98.240 ;
        RECT 130.560 98.070 130.730 98.240 ;
        RECT 131.480 98.070 131.650 98.240 ;
        RECT 131.840 98.070 132.010 98.240 ;
        RECT 132.200 98.070 132.370 98.240 ;
        RECT 133.670 98.020 133.840 98.190 ;
        RECT 134.110 98.020 134.280 98.190 ;
        RECT 134.520 98.020 134.690 98.190 ;
        RECT 134.950 98.020 135.120 98.190 ;
        RECT 135.390 98.020 135.560 98.190 ;
        RECT 135.800 98.020 135.970 98.190 ;
        RECT 137.510 98.020 137.680 98.190 ;
        RECT 137.950 98.020 138.120 98.190 ;
        RECT 138.360 98.020 138.530 98.190 ;
        RECT 138.790 98.020 138.960 98.190 ;
        RECT 139.230 98.020 139.400 98.190 ;
        RECT 139.640 98.020 139.810 98.190 ;
        RECT 5.920 97.590 6.090 97.770 ;
        RECT 6.400 97.590 6.570 97.770 ;
        RECT 6.880 97.590 7.050 97.770 ;
        RECT 7.360 97.590 7.530 97.770 ;
        RECT 7.840 97.590 8.010 97.770 ;
        RECT 8.320 97.590 8.490 97.770 ;
        RECT 8.800 97.590 8.970 97.770 ;
        RECT 9.280 97.590 9.450 97.770 ;
        RECT 9.760 97.590 9.930 97.770 ;
        RECT 10.240 97.590 10.410 97.770 ;
        RECT 10.720 97.590 10.890 97.770 ;
        RECT 11.200 97.590 11.370 97.770 ;
        RECT 11.680 97.590 11.850 97.770 ;
        RECT 12.160 97.590 12.330 97.770 ;
        RECT 12.640 97.590 12.810 97.770 ;
        RECT 13.120 97.590 13.290 97.770 ;
        RECT 13.600 97.590 13.770 97.770 ;
        RECT 14.080 97.590 14.250 97.770 ;
        RECT 14.560 97.590 14.730 97.770 ;
        RECT 15.040 97.590 15.210 97.770 ;
        RECT 15.520 97.590 15.690 97.770 ;
        RECT 16.000 97.590 16.170 97.770 ;
        RECT 16.480 97.590 16.650 97.770 ;
        RECT 16.960 97.590 17.130 97.770 ;
        RECT 17.440 97.590 17.610 97.770 ;
        RECT 17.920 97.590 18.090 97.770 ;
        RECT 18.400 97.590 18.570 97.770 ;
        RECT 18.880 97.590 19.050 97.770 ;
        RECT 19.360 97.590 19.530 97.770 ;
        RECT 19.840 97.590 20.010 97.770 ;
        RECT 20.320 97.590 20.490 97.770 ;
        RECT 20.800 97.590 20.970 97.770 ;
        RECT 21.280 97.590 21.450 97.770 ;
        RECT 21.760 97.760 21.930 97.770 ;
      LAYER li1 ;
        RECT 21.600 97.590 22.080 97.760 ;
      LAYER li1 ;
        RECT 22.240 97.590 22.410 97.770 ;
        RECT 22.720 97.590 22.890 97.770 ;
        RECT 23.200 97.590 23.370 97.770 ;
        RECT 23.680 97.590 23.850 97.770 ;
        RECT 24.160 97.590 24.330 97.770 ;
        RECT 24.640 97.590 24.810 97.770 ;
        RECT 25.120 97.590 25.290 97.770 ;
        RECT 25.600 97.590 25.770 97.770 ;
        RECT 26.080 97.590 26.250 97.770 ;
        RECT 26.560 97.590 26.730 97.770 ;
        RECT 27.040 97.590 27.210 97.770 ;
        RECT 27.520 97.590 27.690 97.770 ;
        RECT 28.000 97.590 28.170 97.770 ;
        RECT 28.480 97.760 28.650 97.770 ;
      LAYER li1 ;
        RECT 28.320 97.590 28.800 97.760 ;
      LAYER li1 ;
        RECT 28.960 97.590 29.130 97.770 ;
        RECT 29.440 97.590 29.610 97.770 ;
        RECT 29.920 97.590 30.090 97.770 ;
        RECT 30.400 97.590 30.570 97.770 ;
        RECT 30.880 97.590 31.050 97.770 ;
        RECT 31.360 97.590 31.530 97.770 ;
        RECT 31.840 97.590 32.010 97.770 ;
        RECT 32.320 97.590 32.490 97.770 ;
      LAYER li1 ;
        RECT 32.640 97.760 33.120 97.770 ;
      LAYER li1 ;
        RECT 32.800 97.590 32.970 97.760 ;
        RECT 33.280 97.590 33.450 97.770 ;
        RECT 33.760 97.590 33.930 97.770 ;
        RECT 34.240 97.590 34.410 97.770 ;
        RECT 34.720 97.590 34.890 97.770 ;
        RECT 35.200 97.590 35.370 97.770 ;
        RECT 35.680 97.590 35.850 97.770 ;
        RECT 36.160 97.590 36.330 97.770 ;
        RECT 36.640 97.590 36.810 97.770 ;
        RECT 37.120 97.590 37.290 97.770 ;
        RECT 37.600 97.590 37.770 97.770 ;
        RECT 38.080 97.590 38.250 97.770 ;
        RECT 38.560 97.590 38.730 97.770 ;
        RECT 39.040 97.590 39.210 97.770 ;
        RECT 39.520 97.590 39.690 97.770 ;
        RECT 40.000 97.590 40.170 97.770 ;
        RECT 40.480 97.590 40.650 97.770 ;
        RECT 40.960 97.590 41.130 97.770 ;
        RECT 41.440 97.590 41.610 97.770 ;
        RECT 41.920 97.590 42.090 97.770 ;
        RECT 42.400 97.590 42.570 97.770 ;
        RECT 42.880 97.590 43.050 97.770 ;
        RECT 43.360 97.590 43.530 97.770 ;
        RECT 43.840 97.590 44.010 97.770 ;
        RECT 44.320 97.590 44.490 97.770 ;
        RECT 44.800 97.590 44.970 97.770 ;
        RECT 45.280 97.590 45.450 97.770 ;
        RECT 45.760 97.590 45.930 97.770 ;
        RECT 46.240 97.590 46.410 97.770 ;
        RECT 46.720 97.590 46.890 97.770 ;
        RECT 47.200 97.590 47.370 97.770 ;
        RECT 47.680 97.590 47.850 97.770 ;
        RECT 48.160 97.590 48.330 97.770 ;
        RECT 48.640 97.590 48.810 97.770 ;
        RECT 49.120 97.590 49.290 97.770 ;
        RECT 49.600 97.590 49.770 97.770 ;
        RECT 50.080 97.590 50.250 97.770 ;
        RECT 50.560 97.590 50.730 97.770 ;
        RECT 51.040 97.590 51.210 97.770 ;
        RECT 51.520 97.590 51.690 97.770 ;
        RECT 52.000 97.590 52.170 97.770 ;
        RECT 52.480 97.590 52.650 97.770 ;
        RECT 52.960 97.590 53.130 97.770 ;
        RECT 53.440 97.590 53.610 97.770 ;
        RECT 53.920 97.590 54.090 97.770 ;
        RECT 54.400 97.590 54.570 97.770 ;
        RECT 54.880 97.590 55.050 97.770 ;
        RECT 55.360 97.590 55.530 97.770 ;
        RECT 55.840 97.590 56.010 97.770 ;
        RECT 56.320 97.590 56.490 97.770 ;
        RECT 56.800 97.590 56.970 97.770 ;
        RECT 57.280 97.590 57.450 97.770 ;
        RECT 57.760 97.590 57.930 97.770 ;
        RECT 58.240 97.590 58.410 97.770 ;
        RECT 58.720 97.590 58.890 97.770 ;
        RECT 59.200 97.590 59.370 97.770 ;
        RECT 59.680 97.590 59.850 97.770 ;
        RECT 60.160 97.590 60.330 97.770 ;
        RECT 60.640 97.590 60.810 97.770 ;
        RECT 61.120 97.590 61.290 97.770 ;
        RECT 61.600 97.590 61.770 97.770 ;
        RECT 62.080 97.590 62.250 97.770 ;
        RECT 62.560 97.590 62.730 97.770 ;
        RECT 63.040 97.590 63.210 97.770 ;
        RECT 63.520 97.590 63.690 97.770 ;
        RECT 64.000 97.590 64.170 97.770 ;
        RECT 64.480 97.590 64.650 97.770 ;
        RECT 64.960 97.590 65.130 97.770 ;
        RECT 65.440 97.590 65.610 97.770 ;
        RECT 65.920 97.590 66.090 97.770 ;
        RECT 66.400 97.590 66.570 97.770 ;
        RECT 66.880 97.590 67.050 97.770 ;
        RECT 67.360 97.590 67.530 97.770 ;
        RECT 67.840 97.590 68.010 97.770 ;
        RECT 68.320 97.590 68.490 97.770 ;
        RECT 68.800 97.590 68.970 97.770 ;
        RECT 69.280 97.590 69.450 97.770 ;
        RECT 69.760 97.590 69.930 97.770 ;
        RECT 70.240 97.590 70.410 97.770 ;
        RECT 70.720 97.590 70.890 97.770 ;
        RECT 71.200 97.590 71.370 97.770 ;
        RECT 71.680 97.590 71.850 97.770 ;
        RECT 72.160 97.760 72.330 97.770 ;
      LAYER li1 ;
        RECT 72.000 97.590 72.480 97.760 ;
      LAYER li1 ;
        RECT 72.640 97.590 72.810 97.770 ;
        RECT 73.120 97.590 73.290 97.770 ;
        RECT 73.600 97.590 73.770 97.770 ;
      LAYER li1 ;
        RECT 73.920 97.760 74.400 97.770 ;
      LAYER li1 ;
        RECT 74.080 97.590 74.250 97.760 ;
        RECT 74.560 97.590 74.730 97.770 ;
        RECT 75.040 97.590 75.210 97.770 ;
        RECT 75.520 97.590 75.690 97.770 ;
        RECT 76.000 97.590 76.170 97.770 ;
        RECT 76.480 97.590 76.650 97.770 ;
        RECT 76.960 97.590 77.130 97.770 ;
        RECT 77.440 97.590 77.610 97.770 ;
        RECT 77.920 97.590 78.090 97.770 ;
        RECT 78.400 97.590 78.570 97.770 ;
        RECT 78.880 97.590 79.050 97.770 ;
        RECT 79.360 97.590 79.530 97.770 ;
        RECT 79.840 97.590 80.010 97.770 ;
        RECT 80.320 97.590 80.490 97.770 ;
        RECT 80.800 97.590 80.970 97.770 ;
        RECT 81.280 97.590 81.450 97.770 ;
        RECT 81.760 97.590 81.930 97.770 ;
        RECT 82.240 97.590 82.410 97.770 ;
        RECT 82.720 97.590 82.890 97.770 ;
        RECT 83.200 97.590 83.370 97.770 ;
        RECT 83.680 97.590 83.850 97.770 ;
        RECT 84.160 97.590 84.330 97.770 ;
        RECT 84.640 97.590 84.810 97.770 ;
        RECT 85.120 97.590 85.290 97.770 ;
        RECT 85.600 97.590 85.770 97.770 ;
        RECT 86.080 97.590 86.250 97.770 ;
        RECT 86.560 97.590 86.730 97.770 ;
        RECT 87.040 97.590 87.210 97.770 ;
        RECT 87.520 97.590 87.690 97.770 ;
        RECT 88.000 97.590 88.170 97.770 ;
        RECT 88.480 97.590 88.650 97.770 ;
        RECT 88.960 97.590 89.130 97.770 ;
        RECT 89.440 97.590 89.610 97.770 ;
        RECT 89.920 97.590 90.090 97.770 ;
        RECT 90.400 97.590 90.570 97.770 ;
        RECT 90.880 97.590 91.050 97.770 ;
        RECT 91.360 97.590 91.530 97.770 ;
        RECT 91.840 97.590 92.010 97.770 ;
        RECT 92.320 97.590 92.490 97.770 ;
        RECT 92.800 97.590 92.970 97.770 ;
        RECT 93.280 97.590 93.450 97.770 ;
        RECT 93.760 97.590 93.930 97.770 ;
        RECT 94.240 97.590 94.410 97.770 ;
        RECT 94.720 97.590 94.890 97.770 ;
        RECT 95.200 97.590 95.370 97.770 ;
        RECT 95.680 97.590 95.850 97.770 ;
        RECT 96.160 97.590 96.330 97.770 ;
        RECT 96.640 97.590 96.810 97.770 ;
        RECT 97.120 97.590 97.290 97.770 ;
        RECT 97.600 97.590 97.770 97.770 ;
        RECT 98.080 97.590 98.250 97.770 ;
      LAYER li1 ;
        RECT 98.400 97.760 98.880 97.770 ;
      LAYER li1 ;
        RECT 98.560 97.590 98.730 97.760 ;
        RECT 99.040 97.590 99.210 97.770 ;
        RECT 99.520 97.590 99.690 97.770 ;
        RECT 100.000 97.590 100.170 97.770 ;
        RECT 100.480 97.590 100.650 97.770 ;
        RECT 100.960 97.590 101.130 97.770 ;
        RECT 101.440 97.590 101.610 97.770 ;
        RECT 101.920 97.590 102.090 97.770 ;
        RECT 102.400 97.590 102.570 97.770 ;
        RECT 102.880 97.590 103.050 97.770 ;
        RECT 103.360 97.590 103.530 97.770 ;
        RECT 103.840 97.590 104.010 97.770 ;
        RECT 104.320 97.590 104.490 97.770 ;
        RECT 104.800 97.590 104.970 97.770 ;
        RECT 105.280 97.590 105.450 97.770 ;
        RECT 105.760 97.590 105.930 97.770 ;
        RECT 106.240 97.590 106.410 97.770 ;
        RECT 106.720 97.590 106.890 97.770 ;
        RECT 107.200 97.590 107.370 97.770 ;
        RECT 107.680 97.590 107.850 97.770 ;
        RECT 108.160 97.590 108.330 97.770 ;
        RECT 108.640 97.590 108.810 97.770 ;
        RECT 109.120 97.590 109.290 97.770 ;
        RECT 109.600 97.590 109.770 97.770 ;
        RECT 110.080 97.590 110.250 97.770 ;
        RECT 110.560 97.590 110.730 97.770 ;
        RECT 111.040 97.590 111.210 97.770 ;
        RECT 111.520 97.590 111.690 97.770 ;
        RECT 112.000 97.590 112.170 97.770 ;
        RECT 112.480 97.590 112.650 97.770 ;
        RECT 112.960 97.590 113.130 97.770 ;
        RECT 113.440 97.590 113.610 97.770 ;
        RECT 113.920 97.590 114.090 97.770 ;
        RECT 114.400 97.590 114.570 97.770 ;
        RECT 114.880 97.590 115.050 97.770 ;
        RECT 115.360 97.590 115.530 97.770 ;
        RECT 115.840 97.590 116.010 97.770 ;
        RECT 116.320 97.590 116.490 97.770 ;
        RECT 116.800 97.590 116.970 97.770 ;
        RECT 117.280 97.590 117.450 97.770 ;
        RECT 117.760 97.590 117.930 97.770 ;
        RECT 118.240 97.590 118.410 97.770 ;
        RECT 118.720 97.590 118.890 97.770 ;
        RECT 119.200 97.590 119.370 97.770 ;
        RECT 119.680 97.590 119.850 97.770 ;
        RECT 120.160 97.590 120.330 97.770 ;
        RECT 120.640 97.590 120.810 97.770 ;
      LAYER li1 ;
        RECT 120.960 97.760 121.440 97.770 ;
      LAYER li1 ;
        RECT 121.120 97.590 121.290 97.760 ;
        RECT 121.600 97.590 121.770 97.770 ;
        RECT 122.080 97.590 122.250 97.770 ;
        RECT 122.560 97.590 122.730 97.770 ;
        RECT 123.040 97.590 123.210 97.770 ;
        RECT 123.520 97.590 123.690 97.770 ;
        RECT 124.000 97.590 124.170 97.770 ;
        RECT 124.480 97.590 124.650 97.770 ;
        RECT 124.960 97.590 125.130 97.770 ;
        RECT 125.440 97.590 125.610 97.770 ;
        RECT 125.920 97.590 126.090 97.770 ;
        RECT 126.400 97.590 126.570 97.770 ;
        RECT 126.880 97.590 127.050 97.770 ;
        RECT 127.360 97.590 127.530 97.770 ;
        RECT 127.840 97.590 128.010 97.770 ;
        RECT 128.320 97.590 128.490 97.770 ;
        RECT 128.800 97.590 128.970 97.770 ;
        RECT 129.280 97.590 129.450 97.770 ;
        RECT 129.760 97.590 129.930 97.770 ;
        RECT 130.240 97.590 130.410 97.770 ;
        RECT 130.720 97.590 130.890 97.770 ;
        RECT 131.200 97.590 131.370 97.770 ;
        RECT 131.680 97.590 131.850 97.770 ;
        RECT 132.160 97.590 132.330 97.770 ;
        RECT 132.640 97.590 132.810 97.770 ;
        RECT 133.120 97.590 133.290 97.770 ;
        RECT 133.600 97.590 133.770 97.770 ;
        RECT 134.080 97.590 134.250 97.770 ;
        RECT 134.560 97.590 134.730 97.770 ;
        RECT 135.040 97.590 135.210 97.770 ;
        RECT 135.520 97.590 135.690 97.770 ;
        RECT 136.000 97.590 136.170 97.770 ;
        RECT 136.480 97.590 136.650 97.770 ;
        RECT 136.960 97.590 137.130 97.770 ;
        RECT 137.440 97.590 137.610 97.770 ;
        RECT 137.920 97.590 138.090 97.770 ;
        RECT 138.400 97.590 138.570 97.770 ;
        RECT 138.880 97.590 139.050 97.770 ;
        RECT 139.360 97.590 139.530 97.770 ;
        RECT 139.840 97.590 140.010 97.770 ;
        RECT 140.320 97.590 140.490 97.770 ;
        RECT 140.800 97.590 140.970 97.770 ;
        RECT 141.280 97.590 141.450 97.770 ;
        RECT 141.760 97.760 141.930 97.770 ;
      LAYER li1 ;
        RECT 141.600 97.590 142.080 97.760 ;
      LAYER li1 ;
        RECT 6.420 97.120 6.590 97.290 ;
        RECT 6.780 97.120 6.950 97.290 ;
        RECT 8.810 97.120 8.980 97.290 ;
        RECT 11.240 97.120 11.410 97.290 ;
        RECT 11.600 97.120 11.770 97.290 ;
        RECT 11.960 97.120 12.130 97.290 ;
        RECT 13.580 97.120 13.750 97.290 ;
        RECT 13.940 97.120 14.110 97.290 ;
        RECT 14.300 97.120 14.470 97.290 ;
        RECT 16.280 97.120 16.450 97.290 ;
        RECT 16.640 97.120 16.810 97.290 ;
        RECT 17.000 97.120 17.170 97.290 ;
        RECT 18.030 97.120 18.200 97.290 ;
        RECT 18.390 97.120 18.560 97.290 ;
        RECT 18.750 97.120 18.920 97.290 ;
        RECT 19.560 97.120 19.730 97.290 ;
        RECT 19.920 97.120 20.090 97.290 ;
        RECT 20.280 97.120 20.450 97.290 ;
        RECT 21.830 97.170 22.000 97.340 ;
        RECT 22.270 97.170 22.440 97.340 ;
        RECT 22.680 97.170 22.850 97.340 ;
        RECT 23.110 97.170 23.280 97.340 ;
        RECT 23.550 97.170 23.720 97.340 ;
        RECT 23.960 97.170 24.130 97.340 ;
        RECT 25.060 97.120 25.230 97.290 ;
        RECT 25.420 97.120 25.590 97.290 ;
        RECT 25.780 97.120 25.950 97.290 ;
        RECT 26.140 97.120 26.310 97.290 ;
        RECT 27.300 97.120 27.470 97.290 ;
        RECT 27.660 97.120 27.830 97.290 ;
        RECT 28.020 97.120 28.190 97.290 ;
        RECT 28.380 97.120 28.550 97.290 ;
        RECT 29.510 97.170 29.680 97.340 ;
        RECT 29.950 97.170 30.120 97.340 ;
        RECT 30.360 97.170 30.530 97.340 ;
        RECT 30.790 97.170 30.960 97.340 ;
        RECT 31.230 97.170 31.400 97.340 ;
        RECT 31.640 97.170 31.810 97.340 ;
        RECT 33.860 97.120 34.030 97.290 ;
        RECT 34.220 97.120 34.390 97.290 ;
        RECT 36.020 97.170 36.190 97.340 ;
        RECT 36.380 97.170 36.550 97.340 ;
        RECT 36.820 97.170 36.990 97.340 ;
        RECT 38.180 97.120 38.350 97.290 ;
        RECT 38.540 97.120 38.710 97.290 ;
        RECT 40.340 97.170 40.510 97.340 ;
        RECT 40.700 97.170 40.870 97.340 ;
        RECT 41.140 97.170 41.310 97.340 ;
        RECT 41.880 97.120 42.050 97.290 ;
        RECT 42.240 97.120 42.410 97.290 ;
        RECT 42.600 97.120 42.770 97.290 ;
        RECT 43.440 97.120 43.610 97.290 ;
        RECT 43.800 97.120 43.970 97.290 ;
        RECT 44.160 97.120 44.330 97.290 ;
        RECT 45.080 97.120 45.250 97.290 ;
        RECT 45.440 97.120 45.610 97.290 ;
        RECT 45.800 97.120 45.970 97.290 ;
        RECT 47.060 97.170 47.230 97.340 ;
        RECT 47.420 97.170 47.590 97.340 ;
        RECT 47.860 97.170 48.030 97.340 ;
        RECT 48.600 97.120 48.770 97.290 ;
        RECT 48.960 97.120 49.130 97.290 ;
        RECT 49.320 97.120 49.490 97.290 ;
        RECT 50.160 97.120 50.330 97.290 ;
        RECT 50.520 97.120 50.690 97.290 ;
        RECT 50.880 97.120 51.050 97.290 ;
        RECT 51.800 97.120 51.970 97.290 ;
        RECT 52.160 97.120 52.330 97.290 ;
        RECT 52.520 97.120 52.690 97.290 ;
        RECT 53.780 97.170 53.950 97.340 ;
        RECT 54.140 97.170 54.310 97.340 ;
        RECT 54.580 97.170 54.750 97.340 ;
        RECT 55.320 97.120 55.490 97.290 ;
        RECT 55.680 97.120 55.850 97.290 ;
        RECT 56.040 97.120 56.210 97.290 ;
        RECT 56.880 97.120 57.050 97.290 ;
        RECT 57.240 97.120 57.410 97.290 ;
        RECT 57.600 97.120 57.770 97.290 ;
        RECT 58.520 97.120 58.690 97.290 ;
        RECT 58.880 97.120 59.050 97.290 ;
        RECT 59.240 97.120 59.410 97.290 ;
        RECT 60.500 97.170 60.670 97.340 ;
        RECT 60.860 97.170 61.030 97.340 ;
        RECT 61.300 97.170 61.470 97.340 ;
        RECT 62.660 97.120 62.830 97.290 ;
        RECT 63.020 97.120 63.190 97.290 ;
        RECT 64.820 97.170 64.990 97.340 ;
        RECT 65.180 97.170 65.350 97.340 ;
        RECT 65.620 97.170 65.790 97.340 ;
        RECT 66.360 97.120 66.530 97.290 ;
        RECT 66.720 97.120 66.890 97.290 ;
        RECT 68.180 97.170 68.350 97.340 ;
        RECT 68.540 97.170 68.710 97.340 ;
        RECT 68.980 97.170 69.150 97.340 ;
        RECT 70.340 97.120 70.510 97.290 ;
        RECT 70.700 97.120 70.870 97.290 ;
        RECT 72.500 97.170 72.670 97.340 ;
        RECT 72.860 97.170 73.030 97.340 ;
        RECT 73.300 97.170 73.470 97.340 ;
        RECT 74.520 97.120 74.690 97.290 ;
        RECT 74.880 97.120 75.050 97.290 ;
        RECT 75.240 97.120 75.410 97.290 ;
        RECT 76.650 97.120 76.820 97.290 ;
        RECT 77.010 97.120 77.180 97.290 ;
        RECT 77.370 97.120 77.540 97.290 ;
        RECT 78.260 97.170 78.430 97.340 ;
        RECT 78.620 97.170 78.790 97.340 ;
        RECT 79.060 97.170 79.230 97.340 ;
        RECT 79.800 97.120 79.970 97.290 ;
        RECT 80.160 97.120 80.330 97.290 ;
        RECT 80.520 97.120 80.690 97.290 ;
        RECT 81.360 97.120 81.530 97.290 ;
        RECT 81.720 97.120 81.890 97.290 ;
        RECT 82.080 97.120 82.250 97.290 ;
        RECT 83.000 97.120 83.170 97.290 ;
        RECT 83.360 97.120 83.530 97.290 ;
        RECT 83.720 97.120 83.890 97.290 ;
        RECT 84.980 97.170 85.150 97.340 ;
        RECT 85.340 97.170 85.510 97.340 ;
        RECT 85.780 97.170 85.950 97.340 ;
        RECT 86.520 97.120 86.690 97.290 ;
        RECT 86.880 97.120 87.050 97.290 ;
        RECT 87.240 97.120 87.410 97.290 ;
        RECT 88.080 97.120 88.250 97.290 ;
        RECT 88.440 97.120 88.610 97.290 ;
        RECT 88.800 97.120 88.970 97.290 ;
        RECT 89.720 97.120 89.890 97.290 ;
        RECT 90.080 97.120 90.250 97.290 ;
        RECT 90.440 97.120 90.610 97.290 ;
        RECT 91.700 97.170 91.870 97.340 ;
        RECT 92.060 97.170 92.230 97.340 ;
        RECT 92.500 97.170 92.670 97.340 ;
        RECT 93.240 97.120 93.410 97.290 ;
        RECT 93.600 97.120 93.770 97.290 ;
        RECT 93.960 97.120 94.130 97.290 ;
        RECT 94.320 97.120 94.490 97.290 ;
        RECT 94.680 97.120 94.850 97.290 ;
        RECT 96.980 97.170 97.150 97.340 ;
        RECT 97.340 97.170 97.510 97.340 ;
        RECT 97.780 97.170 97.950 97.340 ;
        RECT 99.000 97.120 99.170 97.290 ;
        RECT 99.360 97.120 99.530 97.290 ;
        RECT 99.720 97.120 99.890 97.290 ;
        RECT 100.560 97.120 100.730 97.290 ;
        RECT 100.920 97.120 101.090 97.290 ;
        RECT 101.280 97.120 101.450 97.290 ;
        RECT 102.200 97.120 102.370 97.290 ;
        RECT 102.560 97.120 102.730 97.290 ;
        RECT 102.920 97.120 103.090 97.290 ;
        RECT 104.180 97.170 104.350 97.340 ;
        RECT 104.540 97.170 104.710 97.340 ;
        RECT 104.980 97.170 105.150 97.340 ;
        RECT 105.720 97.120 105.890 97.290 ;
        RECT 106.080 97.120 106.250 97.290 ;
        RECT 106.440 97.120 106.610 97.290 ;
        RECT 107.280 97.120 107.450 97.290 ;
        RECT 107.640 97.120 107.810 97.290 ;
        RECT 108.000 97.120 108.170 97.290 ;
        RECT 108.920 97.120 109.090 97.290 ;
        RECT 109.280 97.120 109.450 97.290 ;
        RECT 109.640 97.120 109.810 97.290 ;
        RECT 110.900 97.170 111.070 97.340 ;
        RECT 111.260 97.170 111.430 97.340 ;
        RECT 111.700 97.170 111.870 97.340 ;
        RECT 112.440 97.120 112.610 97.290 ;
        RECT 112.800 97.120 112.970 97.290 ;
        RECT 113.160 97.120 113.330 97.290 ;
        RECT 113.520 97.120 113.690 97.290 ;
        RECT 113.880 97.120 114.050 97.290 ;
        RECT 115.220 97.170 115.390 97.340 ;
        RECT 115.580 97.170 115.750 97.340 ;
        RECT 116.020 97.170 116.190 97.340 ;
        RECT 117.380 97.120 117.550 97.290 ;
        RECT 117.740 97.120 117.910 97.290 ;
        RECT 119.540 97.170 119.710 97.340 ;
        RECT 119.900 97.170 120.070 97.340 ;
        RECT 120.340 97.170 120.510 97.340 ;
        RECT 121.560 97.120 121.730 97.290 ;
        RECT 121.920 97.120 122.090 97.290 ;
        RECT 122.280 97.120 122.450 97.290 ;
        RECT 123.120 97.120 123.290 97.290 ;
        RECT 123.480 97.120 123.650 97.290 ;
        RECT 123.840 97.120 124.010 97.290 ;
        RECT 124.760 97.120 124.930 97.290 ;
        RECT 125.120 97.120 125.290 97.290 ;
        RECT 125.480 97.120 125.650 97.290 ;
        RECT 126.740 97.170 126.910 97.340 ;
        RECT 127.100 97.170 127.270 97.340 ;
        RECT 127.540 97.170 127.710 97.340 ;
        RECT 128.900 97.120 129.070 97.290 ;
        RECT 129.260 97.120 129.430 97.290 ;
        RECT 131.270 97.170 131.440 97.340 ;
        RECT 131.710 97.170 131.880 97.340 ;
        RECT 132.120 97.170 132.290 97.340 ;
        RECT 132.550 97.170 132.720 97.340 ;
        RECT 132.990 97.170 133.160 97.340 ;
        RECT 133.400 97.170 133.570 97.340 ;
        RECT 135.110 97.170 135.280 97.340 ;
        RECT 135.550 97.170 135.720 97.340 ;
        RECT 135.960 97.170 136.130 97.340 ;
        RECT 136.390 97.170 136.560 97.340 ;
        RECT 136.830 97.170 137.000 97.340 ;
        RECT 137.240 97.170 137.410 97.340 ;
        RECT 138.950 97.170 139.120 97.340 ;
        RECT 139.390 97.170 139.560 97.340 ;
        RECT 139.800 97.170 139.970 97.340 ;
        RECT 140.230 97.170 140.400 97.340 ;
        RECT 140.670 97.170 140.840 97.340 ;
        RECT 141.080 97.170 141.250 97.340 ;
        RECT 6.470 89.880 6.640 90.050 ;
        RECT 6.910 89.880 7.080 90.050 ;
        RECT 7.320 89.880 7.490 90.050 ;
        RECT 7.750 89.880 7.920 90.050 ;
        RECT 8.190 89.880 8.360 90.050 ;
        RECT 8.600 89.880 8.770 90.050 ;
        RECT 10.100 89.880 10.270 90.050 ;
        RECT 10.460 89.880 10.630 90.050 ;
        RECT 10.900 89.880 11.070 90.050 ;
        RECT 13.700 89.930 13.870 90.100 ;
        RECT 14.060 89.930 14.230 90.100 ;
        RECT 16.070 89.880 16.240 90.050 ;
        RECT 16.510 89.880 16.680 90.050 ;
        RECT 16.920 89.880 17.090 90.050 ;
        RECT 17.350 89.880 17.520 90.050 ;
        RECT 17.790 89.880 17.960 90.050 ;
        RECT 18.200 89.880 18.370 90.050 ;
        RECT 19.910 89.880 20.080 90.050 ;
        RECT 20.350 89.880 20.520 90.050 ;
        RECT 20.760 89.880 20.930 90.050 ;
        RECT 21.190 89.880 21.360 90.050 ;
        RECT 21.630 89.880 21.800 90.050 ;
        RECT 22.040 89.880 22.210 90.050 ;
        RECT 24.120 89.930 24.290 90.100 ;
        RECT 24.480 89.930 24.650 90.100 ;
        RECT 25.940 89.880 26.110 90.050 ;
        RECT 26.300 89.880 26.470 90.050 ;
        RECT 26.740 89.880 26.910 90.050 ;
        RECT 27.460 89.930 27.630 90.100 ;
        RECT 27.820 89.930 27.990 90.100 ;
        RECT 28.180 89.930 28.350 90.100 ;
        RECT 28.540 89.930 28.710 90.100 ;
        RECT 29.700 89.930 29.870 90.100 ;
        RECT 30.060 89.930 30.230 90.100 ;
        RECT 30.420 89.930 30.590 90.100 ;
        RECT 30.780 89.930 30.950 90.100 ;
        RECT 31.700 89.880 31.870 90.050 ;
        RECT 32.060 89.880 32.230 90.050 ;
        RECT 32.500 89.880 32.670 90.050 ;
        RECT 33.860 89.930 34.030 90.100 ;
        RECT 34.220 89.930 34.390 90.100 ;
        RECT 36.020 89.880 36.190 90.050 ;
        RECT 36.380 89.880 36.550 90.050 ;
        RECT 36.820 89.880 36.990 90.050 ;
        RECT 38.020 89.930 38.190 90.100 ;
        RECT 38.380 89.930 38.550 90.100 ;
        RECT 38.740 89.930 38.910 90.100 ;
        RECT 39.710 89.930 39.880 90.100 ;
        RECT 43.080 89.930 43.250 90.100 ;
        RECT 44.550 89.930 44.720 90.100 ;
        RECT 44.910 89.930 45.080 90.100 ;
        RECT 45.270 89.930 45.440 90.100 ;
        RECT 47.480 89.930 47.650 90.100 ;
        RECT 47.840 89.930 48.010 90.100 ;
        RECT 48.200 89.930 48.370 90.100 ;
        RECT 49.200 89.930 49.370 90.100 ;
        RECT 49.560 89.930 49.730 90.100 ;
        RECT 49.920 89.930 50.090 90.100 ;
        RECT 50.760 89.930 50.930 90.100 ;
        RECT 51.120 89.930 51.290 90.100 ;
        RECT 51.480 89.930 51.650 90.100 ;
        RECT 53.030 89.880 53.200 90.050 ;
        RECT 53.470 89.880 53.640 90.050 ;
        RECT 53.880 89.880 54.050 90.050 ;
        RECT 54.310 89.880 54.480 90.050 ;
        RECT 54.750 89.880 54.920 90.050 ;
        RECT 55.160 89.880 55.330 90.050 ;
        RECT 57.300 89.930 57.470 90.100 ;
        RECT 57.660 89.930 57.830 90.100 ;
        RECT 59.690 89.930 59.860 90.100 ;
        RECT 62.120 89.930 62.290 90.100 ;
        RECT 62.480 89.930 62.650 90.100 ;
        RECT 62.840 89.930 63.010 90.100 ;
        RECT 64.460 89.930 64.630 90.100 ;
        RECT 64.820 89.930 64.990 90.100 ;
        RECT 65.180 89.930 65.350 90.100 ;
        RECT 67.160 89.930 67.330 90.100 ;
        RECT 67.520 89.930 67.690 90.100 ;
        RECT 67.880 89.930 68.050 90.100 ;
        RECT 68.910 89.930 69.080 90.100 ;
        RECT 69.270 89.930 69.440 90.100 ;
        RECT 69.630 89.930 69.800 90.100 ;
        RECT 70.440 89.930 70.610 90.100 ;
        RECT 70.800 89.930 70.970 90.100 ;
        RECT 71.160 89.930 71.330 90.100 ;
        RECT 72.500 89.880 72.670 90.050 ;
        RECT 72.860 89.880 73.030 90.050 ;
        RECT 73.300 89.880 73.470 90.050 ;
        RECT 75.000 89.930 75.170 90.100 ;
        RECT 75.360 89.930 75.530 90.100 ;
        RECT 75.720 89.930 75.890 90.100 ;
        RECT 76.560 89.930 76.730 90.100 ;
        RECT 76.920 89.930 77.090 90.100 ;
        RECT 77.280 89.930 77.450 90.100 ;
        RECT 78.200 89.930 78.370 90.100 ;
        RECT 78.560 89.930 78.730 90.100 ;
        RECT 78.920 89.930 79.090 90.100 ;
        RECT 80.180 89.880 80.350 90.050 ;
        RECT 80.540 89.880 80.710 90.050 ;
        RECT 80.980 89.880 81.150 90.050 ;
        RECT 81.720 89.930 81.890 90.100 ;
        RECT 82.080 89.930 82.250 90.100 ;
        RECT 82.440 89.930 82.610 90.100 ;
        RECT 83.280 89.930 83.450 90.100 ;
        RECT 83.640 89.930 83.810 90.100 ;
        RECT 84.000 89.930 84.170 90.100 ;
        RECT 84.920 89.930 85.090 90.100 ;
        RECT 85.280 89.930 85.450 90.100 ;
        RECT 85.640 89.930 85.810 90.100 ;
        RECT 86.900 89.880 87.070 90.050 ;
        RECT 87.260 89.880 87.430 90.050 ;
        RECT 87.700 89.880 87.870 90.050 ;
        RECT 88.440 89.930 88.610 90.100 ;
        RECT 88.800 89.930 88.970 90.100 ;
        RECT 89.160 89.930 89.330 90.100 ;
        RECT 90.000 89.930 90.170 90.100 ;
        RECT 90.360 89.930 90.530 90.100 ;
        RECT 90.720 89.930 90.890 90.100 ;
        RECT 91.640 89.930 91.810 90.100 ;
        RECT 92.000 89.930 92.170 90.100 ;
        RECT 92.360 89.930 92.530 90.100 ;
        RECT 93.620 89.880 93.790 90.050 ;
        RECT 93.980 89.880 94.150 90.050 ;
        RECT 94.420 89.880 94.590 90.050 ;
        RECT 95.160 89.930 95.330 90.100 ;
        RECT 95.520 89.930 95.690 90.100 ;
        RECT 95.880 89.930 96.050 90.100 ;
        RECT 96.720 89.930 96.890 90.100 ;
        RECT 97.080 89.930 97.250 90.100 ;
        RECT 97.440 89.930 97.610 90.100 ;
        RECT 98.360 89.930 98.530 90.100 ;
        RECT 98.720 89.930 98.890 90.100 ;
        RECT 99.080 89.930 99.250 90.100 ;
        RECT 100.340 89.880 100.510 90.050 ;
        RECT 100.700 89.880 100.870 90.050 ;
        RECT 101.140 89.880 101.310 90.050 ;
        RECT 101.880 89.930 102.050 90.100 ;
        RECT 102.240 89.930 102.410 90.100 ;
        RECT 102.600 89.930 102.770 90.100 ;
        RECT 103.440 89.930 103.610 90.100 ;
        RECT 103.800 89.930 103.970 90.100 ;
        RECT 104.160 89.930 104.330 90.100 ;
        RECT 105.080 89.930 105.250 90.100 ;
        RECT 105.440 89.930 105.610 90.100 ;
        RECT 105.800 89.930 105.970 90.100 ;
        RECT 107.060 89.880 107.230 90.050 ;
        RECT 107.420 89.880 107.590 90.050 ;
        RECT 107.860 89.880 108.030 90.050 ;
        RECT 108.600 89.930 108.770 90.100 ;
        RECT 108.960 89.930 109.130 90.100 ;
        RECT 109.320 89.930 109.490 90.100 ;
        RECT 110.730 89.930 110.900 90.100 ;
        RECT 111.090 89.930 111.260 90.100 ;
        RECT 111.450 89.930 111.620 90.100 ;
        RECT 112.340 89.880 112.510 90.050 ;
        RECT 112.700 89.880 112.870 90.050 ;
        RECT 113.140 89.880 113.310 90.050 ;
        RECT 113.880 89.930 114.050 90.100 ;
        RECT 114.240 89.930 114.410 90.100 ;
        RECT 115.700 89.880 115.870 90.050 ;
        RECT 116.060 89.880 116.230 90.050 ;
        RECT 116.500 89.880 116.670 90.050 ;
        RECT 117.860 89.930 118.030 90.100 ;
        RECT 118.220 89.930 118.390 90.100 ;
        RECT 120.020 89.880 120.190 90.050 ;
        RECT 120.380 89.880 120.550 90.050 ;
        RECT 120.820 89.880 120.990 90.050 ;
        RECT 121.560 89.930 121.730 90.100 ;
        RECT 121.920 89.930 122.090 90.100 ;
        RECT 122.280 89.930 122.450 90.100 ;
        RECT 123.120 89.930 123.290 90.100 ;
        RECT 123.480 89.930 123.650 90.100 ;
        RECT 123.840 89.930 124.010 90.100 ;
        RECT 124.760 89.930 124.930 90.100 ;
        RECT 125.120 89.930 125.290 90.100 ;
        RECT 125.480 89.930 125.650 90.100 ;
        RECT 126.950 89.880 127.120 90.050 ;
        RECT 127.390 89.880 127.560 90.050 ;
        RECT 127.800 89.880 127.970 90.050 ;
        RECT 128.230 89.880 128.400 90.050 ;
        RECT 128.670 89.880 128.840 90.050 ;
        RECT 129.080 89.880 129.250 90.050 ;
        RECT 130.790 89.880 130.960 90.050 ;
        RECT 131.230 89.880 131.400 90.050 ;
        RECT 131.640 89.880 131.810 90.050 ;
        RECT 132.070 89.880 132.240 90.050 ;
        RECT 132.510 89.880 132.680 90.050 ;
        RECT 132.920 89.880 133.090 90.050 ;
        RECT 134.630 89.880 134.800 90.050 ;
        RECT 135.070 89.880 135.240 90.050 ;
        RECT 135.480 89.880 135.650 90.050 ;
        RECT 135.910 89.880 136.080 90.050 ;
        RECT 136.350 89.880 136.520 90.050 ;
        RECT 136.760 89.880 136.930 90.050 ;
        RECT 138.470 89.880 138.640 90.050 ;
        RECT 138.910 89.880 139.080 90.050 ;
        RECT 139.320 89.880 139.490 90.050 ;
        RECT 139.750 89.880 139.920 90.050 ;
        RECT 140.190 89.880 140.360 90.050 ;
        RECT 140.600 89.880 140.770 90.050 ;
        RECT 5.920 89.450 6.090 89.630 ;
        RECT 6.400 89.450 6.570 89.630 ;
        RECT 6.880 89.450 7.050 89.630 ;
        RECT 7.360 89.450 7.530 89.630 ;
        RECT 7.840 89.450 8.010 89.630 ;
        RECT 8.320 89.450 8.490 89.630 ;
        RECT 8.800 89.450 8.970 89.630 ;
        RECT 9.280 89.450 9.450 89.630 ;
        RECT 9.760 89.450 9.930 89.630 ;
        RECT 10.240 89.450 10.410 89.630 ;
        RECT 10.720 89.450 10.890 89.630 ;
        RECT 11.200 89.450 11.370 89.630 ;
        RECT 11.680 89.450 11.850 89.630 ;
        RECT 12.160 89.450 12.330 89.630 ;
        RECT 12.640 89.620 12.810 89.630 ;
      LAYER li1 ;
        RECT 12.480 89.450 12.960 89.620 ;
      LAYER li1 ;
        RECT 13.120 89.450 13.290 89.630 ;
        RECT 13.600 89.450 13.770 89.630 ;
        RECT 14.080 89.450 14.250 89.630 ;
        RECT 14.560 89.450 14.730 89.630 ;
        RECT 15.040 89.450 15.210 89.630 ;
        RECT 15.520 89.450 15.690 89.630 ;
        RECT 16.000 89.450 16.170 89.630 ;
        RECT 16.480 89.450 16.650 89.630 ;
        RECT 16.960 89.450 17.130 89.630 ;
        RECT 17.440 89.450 17.610 89.630 ;
        RECT 17.920 89.450 18.090 89.630 ;
        RECT 18.400 89.450 18.570 89.630 ;
        RECT 18.880 89.450 19.050 89.630 ;
        RECT 19.360 89.450 19.530 89.630 ;
        RECT 19.840 89.450 20.010 89.630 ;
      LAYER li1 ;
        RECT 20.160 89.460 20.640 89.630 ;
      LAYER li1 ;
        RECT 20.320 89.450 20.490 89.460 ;
        RECT 20.800 89.450 20.970 89.630 ;
        RECT 21.280 89.450 21.450 89.630 ;
        RECT 21.760 89.450 21.930 89.630 ;
        RECT 22.240 89.450 22.410 89.630 ;
        RECT 22.720 89.450 22.890 89.630 ;
        RECT 23.200 89.450 23.370 89.630 ;
        RECT 23.680 89.450 23.850 89.630 ;
        RECT 24.160 89.450 24.330 89.630 ;
        RECT 24.640 89.450 24.810 89.630 ;
        RECT 25.120 89.450 25.290 89.630 ;
        RECT 25.600 89.450 25.770 89.630 ;
        RECT 26.080 89.450 26.250 89.630 ;
        RECT 26.560 89.450 26.730 89.630 ;
        RECT 27.040 89.450 27.210 89.630 ;
        RECT 27.520 89.450 27.690 89.630 ;
        RECT 28.000 89.450 28.170 89.630 ;
        RECT 28.480 89.450 28.650 89.630 ;
        RECT 28.960 89.450 29.130 89.630 ;
        RECT 29.440 89.450 29.610 89.630 ;
        RECT 29.920 89.450 30.090 89.630 ;
        RECT 30.400 89.450 30.570 89.630 ;
        RECT 30.880 89.450 31.050 89.630 ;
        RECT 31.360 89.450 31.530 89.630 ;
        RECT 31.840 89.450 32.010 89.630 ;
        RECT 32.320 89.450 32.490 89.630 ;
        RECT 32.800 89.450 32.970 89.630 ;
        RECT 33.280 89.450 33.450 89.630 ;
        RECT 33.760 89.450 33.930 89.630 ;
        RECT 34.240 89.450 34.410 89.630 ;
        RECT 34.720 89.450 34.890 89.630 ;
        RECT 35.200 89.450 35.370 89.630 ;
        RECT 35.680 89.450 35.850 89.630 ;
        RECT 36.160 89.450 36.330 89.630 ;
        RECT 36.640 89.450 36.810 89.630 ;
        RECT 37.120 89.450 37.290 89.630 ;
        RECT 37.600 89.450 37.770 89.630 ;
        RECT 38.080 89.450 38.250 89.630 ;
        RECT 38.560 89.450 38.730 89.630 ;
        RECT 39.040 89.450 39.210 89.630 ;
        RECT 39.520 89.450 39.690 89.630 ;
        RECT 40.000 89.450 40.170 89.630 ;
        RECT 40.480 89.450 40.650 89.630 ;
        RECT 40.960 89.450 41.130 89.630 ;
        RECT 41.440 89.450 41.610 89.630 ;
        RECT 41.920 89.450 42.090 89.630 ;
        RECT 42.400 89.450 42.570 89.630 ;
        RECT 42.880 89.450 43.050 89.630 ;
        RECT 43.360 89.450 43.530 89.630 ;
        RECT 43.840 89.450 44.010 89.630 ;
        RECT 44.320 89.450 44.490 89.630 ;
        RECT 44.800 89.450 44.970 89.630 ;
        RECT 45.280 89.450 45.450 89.630 ;
        RECT 45.760 89.450 45.930 89.630 ;
        RECT 46.240 89.450 46.410 89.630 ;
        RECT 46.720 89.450 46.890 89.630 ;
        RECT 47.200 89.450 47.370 89.630 ;
        RECT 47.680 89.450 47.850 89.630 ;
        RECT 48.160 89.450 48.330 89.630 ;
        RECT 48.640 89.450 48.810 89.630 ;
        RECT 49.120 89.450 49.290 89.630 ;
        RECT 49.600 89.450 49.770 89.630 ;
        RECT 50.080 89.450 50.250 89.630 ;
        RECT 50.560 89.450 50.730 89.630 ;
        RECT 51.040 89.450 51.210 89.630 ;
        RECT 51.520 89.450 51.690 89.630 ;
        RECT 52.000 89.450 52.170 89.630 ;
        RECT 52.480 89.450 52.650 89.630 ;
        RECT 52.960 89.450 53.130 89.630 ;
        RECT 53.440 89.450 53.610 89.630 ;
        RECT 53.920 89.450 54.090 89.630 ;
        RECT 54.400 89.450 54.570 89.630 ;
        RECT 54.880 89.450 55.050 89.630 ;
        RECT 55.360 89.450 55.530 89.630 ;
        RECT 55.840 89.450 56.010 89.630 ;
        RECT 56.320 89.620 56.490 89.630 ;
      LAYER li1 ;
        RECT 56.160 89.450 56.640 89.620 ;
      LAYER li1 ;
        RECT 56.800 89.450 56.970 89.630 ;
        RECT 57.280 89.450 57.450 89.630 ;
        RECT 57.760 89.450 57.930 89.630 ;
        RECT 58.240 89.450 58.410 89.630 ;
        RECT 58.720 89.450 58.890 89.630 ;
        RECT 59.200 89.450 59.370 89.630 ;
        RECT 59.680 89.450 59.850 89.630 ;
        RECT 60.160 89.450 60.330 89.630 ;
        RECT 60.640 89.450 60.810 89.630 ;
        RECT 61.120 89.450 61.290 89.630 ;
        RECT 61.600 89.450 61.770 89.630 ;
        RECT 62.080 89.450 62.250 89.630 ;
        RECT 62.560 89.450 62.730 89.630 ;
        RECT 63.040 89.450 63.210 89.630 ;
        RECT 63.520 89.450 63.690 89.630 ;
        RECT 64.000 89.450 64.170 89.630 ;
        RECT 64.480 89.450 64.650 89.630 ;
        RECT 64.960 89.450 65.130 89.630 ;
        RECT 65.440 89.450 65.610 89.630 ;
        RECT 65.920 89.450 66.090 89.630 ;
        RECT 66.400 89.450 66.570 89.630 ;
        RECT 66.880 89.450 67.050 89.630 ;
        RECT 67.360 89.450 67.530 89.630 ;
        RECT 67.840 89.450 68.010 89.630 ;
      LAYER li1 ;
        RECT 68.160 89.460 68.640 89.630 ;
      LAYER li1 ;
        RECT 68.320 89.450 68.490 89.460 ;
        RECT 68.800 89.450 68.970 89.630 ;
        RECT 69.280 89.450 69.450 89.630 ;
        RECT 69.760 89.450 69.930 89.630 ;
        RECT 70.240 89.450 70.410 89.630 ;
        RECT 70.720 89.450 70.890 89.630 ;
        RECT 71.200 89.450 71.370 89.630 ;
        RECT 71.680 89.450 71.850 89.630 ;
        RECT 72.160 89.450 72.330 89.630 ;
        RECT 72.640 89.450 72.810 89.630 ;
        RECT 73.120 89.450 73.290 89.630 ;
        RECT 73.600 89.450 73.770 89.630 ;
        RECT 74.080 89.450 74.250 89.630 ;
        RECT 74.560 89.450 74.730 89.630 ;
        RECT 75.040 89.450 75.210 89.630 ;
        RECT 75.520 89.450 75.690 89.630 ;
        RECT 76.000 89.450 76.170 89.630 ;
        RECT 76.480 89.450 76.650 89.630 ;
        RECT 76.960 89.450 77.130 89.630 ;
        RECT 77.440 89.450 77.610 89.630 ;
        RECT 77.920 89.450 78.090 89.630 ;
        RECT 78.400 89.450 78.570 89.630 ;
        RECT 78.880 89.450 79.050 89.630 ;
        RECT 79.360 89.450 79.530 89.630 ;
        RECT 79.840 89.450 80.010 89.630 ;
        RECT 80.320 89.450 80.490 89.630 ;
        RECT 80.800 89.450 80.970 89.630 ;
        RECT 81.280 89.450 81.450 89.630 ;
        RECT 81.760 89.450 81.930 89.630 ;
        RECT 82.240 89.450 82.410 89.630 ;
        RECT 82.720 89.450 82.890 89.630 ;
        RECT 83.200 89.450 83.370 89.630 ;
        RECT 83.680 89.450 83.850 89.630 ;
        RECT 84.160 89.450 84.330 89.630 ;
        RECT 84.640 89.450 84.810 89.630 ;
        RECT 85.120 89.450 85.290 89.630 ;
        RECT 85.600 89.450 85.770 89.630 ;
        RECT 86.080 89.450 86.250 89.630 ;
        RECT 86.560 89.450 86.730 89.630 ;
        RECT 87.040 89.450 87.210 89.630 ;
        RECT 87.520 89.450 87.690 89.630 ;
        RECT 88.000 89.450 88.170 89.630 ;
        RECT 88.480 89.450 88.650 89.630 ;
        RECT 88.960 89.450 89.130 89.630 ;
        RECT 89.440 89.450 89.610 89.630 ;
        RECT 89.920 89.450 90.090 89.630 ;
        RECT 90.400 89.450 90.570 89.630 ;
        RECT 90.880 89.450 91.050 89.630 ;
        RECT 91.360 89.450 91.530 89.630 ;
        RECT 91.840 89.450 92.010 89.630 ;
        RECT 92.320 89.450 92.490 89.630 ;
        RECT 92.800 89.450 92.970 89.630 ;
        RECT 93.280 89.450 93.450 89.630 ;
        RECT 93.760 89.450 93.930 89.630 ;
        RECT 94.240 89.450 94.410 89.630 ;
        RECT 94.720 89.450 94.890 89.630 ;
        RECT 95.200 89.450 95.370 89.630 ;
        RECT 95.680 89.450 95.850 89.630 ;
        RECT 96.160 89.450 96.330 89.630 ;
        RECT 96.640 89.450 96.810 89.630 ;
        RECT 97.120 89.450 97.290 89.630 ;
        RECT 97.600 89.450 97.770 89.630 ;
        RECT 98.080 89.450 98.250 89.630 ;
        RECT 98.560 89.450 98.730 89.630 ;
        RECT 99.040 89.450 99.210 89.630 ;
        RECT 99.520 89.450 99.690 89.630 ;
        RECT 100.000 89.450 100.170 89.630 ;
        RECT 100.480 89.450 100.650 89.630 ;
        RECT 100.960 89.450 101.130 89.630 ;
      LAYER li1 ;
        RECT 101.280 89.460 101.760 89.630 ;
      LAYER li1 ;
        RECT 101.440 89.450 101.610 89.460 ;
        RECT 101.920 89.450 102.090 89.630 ;
        RECT 102.400 89.450 102.570 89.630 ;
        RECT 102.880 89.450 103.050 89.630 ;
        RECT 103.360 89.450 103.530 89.630 ;
        RECT 103.840 89.450 104.010 89.630 ;
        RECT 104.320 89.450 104.490 89.630 ;
        RECT 104.800 89.450 104.970 89.630 ;
        RECT 105.280 89.450 105.450 89.630 ;
        RECT 105.760 89.450 105.930 89.630 ;
        RECT 106.240 89.450 106.410 89.630 ;
        RECT 106.720 89.450 106.890 89.630 ;
        RECT 107.200 89.450 107.370 89.630 ;
        RECT 107.680 89.450 107.850 89.630 ;
        RECT 108.160 89.450 108.330 89.630 ;
        RECT 108.640 89.450 108.810 89.630 ;
        RECT 109.120 89.450 109.290 89.630 ;
        RECT 109.600 89.450 109.770 89.630 ;
        RECT 110.080 89.450 110.250 89.630 ;
        RECT 110.560 89.450 110.730 89.630 ;
        RECT 111.040 89.450 111.210 89.630 ;
        RECT 111.520 89.450 111.690 89.630 ;
        RECT 112.000 89.450 112.170 89.630 ;
        RECT 112.480 89.450 112.650 89.630 ;
        RECT 112.960 89.450 113.130 89.630 ;
        RECT 113.440 89.450 113.610 89.630 ;
        RECT 113.920 89.450 114.090 89.630 ;
        RECT 114.400 89.450 114.570 89.630 ;
        RECT 114.880 89.450 115.050 89.630 ;
        RECT 115.360 89.450 115.530 89.630 ;
        RECT 115.840 89.450 116.010 89.630 ;
        RECT 116.320 89.450 116.490 89.630 ;
        RECT 116.800 89.450 116.970 89.630 ;
        RECT 117.280 89.450 117.450 89.630 ;
      LAYER li1 ;
        RECT 117.600 89.620 118.080 89.630 ;
      LAYER li1 ;
        RECT 117.760 89.450 117.930 89.620 ;
        RECT 118.240 89.450 118.410 89.630 ;
        RECT 118.720 89.450 118.890 89.630 ;
        RECT 119.200 89.450 119.370 89.630 ;
        RECT 119.680 89.450 119.850 89.630 ;
        RECT 120.160 89.450 120.330 89.630 ;
        RECT 120.640 89.450 120.810 89.630 ;
        RECT 121.120 89.450 121.290 89.630 ;
        RECT 121.600 89.450 121.770 89.630 ;
        RECT 122.080 89.450 122.250 89.630 ;
        RECT 122.560 89.450 122.730 89.630 ;
        RECT 123.040 89.450 123.210 89.630 ;
        RECT 123.520 89.450 123.690 89.630 ;
        RECT 124.000 89.450 124.170 89.630 ;
        RECT 124.480 89.450 124.650 89.630 ;
        RECT 124.960 89.450 125.130 89.630 ;
        RECT 125.440 89.450 125.610 89.630 ;
        RECT 125.920 89.450 126.090 89.630 ;
        RECT 126.400 89.450 126.570 89.630 ;
        RECT 126.880 89.450 127.050 89.630 ;
        RECT 127.360 89.450 127.530 89.630 ;
        RECT 127.840 89.450 128.010 89.630 ;
        RECT 128.320 89.450 128.490 89.630 ;
        RECT 128.800 89.450 128.970 89.630 ;
        RECT 129.280 89.450 129.450 89.630 ;
        RECT 129.760 89.450 129.930 89.630 ;
        RECT 130.240 89.450 130.410 89.630 ;
        RECT 130.720 89.450 130.890 89.630 ;
        RECT 131.200 89.450 131.370 89.630 ;
        RECT 131.680 89.450 131.850 89.630 ;
        RECT 132.160 89.450 132.330 89.630 ;
        RECT 132.640 89.450 132.810 89.630 ;
        RECT 133.120 89.450 133.290 89.630 ;
        RECT 133.600 89.450 133.770 89.630 ;
      LAYER li1 ;
        RECT 133.920 89.460 134.400 89.630 ;
      LAYER li1 ;
        RECT 134.080 89.450 134.250 89.460 ;
        RECT 134.560 89.450 134.730 89.630 ;
        RECT 135.040 89.450 135.210 89.630 ;
        RECT 135.520 89.450 135.690 89.630 ;
        RECT 136.000 89.450 136.170 89.630 ;
        RECT 136.480 89.450 136.650 89.630 ;
        RECT 136.960 89.450 137.130 89.630 ;
        RECT 137.440 89.450 137.610 89.630 ;
        RECT 137.920 89.450 138.090 89.630 ;
        RECT 138.400 89.450 138.570 89.630 ;
        RECT 138.880 89.450 139.050 89.630 ;
        RECT 139.360 89.450 139.530 89.630 ;
        RECT 139.840 89.450 140.010 89.630 ;
        RECT 140.320 89.450 140.490 89.630 ;
        RECT 140.800 89.450 140.970 89.630 ;
        RECT 141.280 89.450 141.450 89.630 ;
      LAYER li1 ;
        RECT 141.600 89.450 142.080 89.630 ;
      LAYER li1 ;
        RECT 6.470 89.030 6.640 89.200 ;
        RECT 6.910 89.030 7.080 89.200 ;
        RECT 7.320 89.030 7.490 89.200 ;
        RECT 7.750 89.030 7.920 89.200 ;
        RECT 8.190 89.030 8.360 89.200 ;
        RECT 8.600 89.030 8.770 89.200 ;
        RECT 10.310 89.030 10.480 89.200 ;
        RECT 10.750 89.030 10.920 89.200 ;
        RECT 11.160 89.030 11.330 89.200 ;
        RECT 11.590 89.030 11.760 89.200 ;
        RECT 12.030 89.030 12.200 89.200 ;
        RECT 12.440 89.030 12.610 89.200 ;
        RECT 14.150 89.030 14.320 89.200 ;
        RECT 14.590 89.030 14.760 89.200 ;
        RECT 15.000 89.030 15.170 89.200 ;
        RECT 15.430 89.030 15.600 89.200 ;
        RECT 15.870 89.030 16.040 89.200 ;
        RECT 16.280 89.030 16.450 89.200 ;
        RECT 17.780 89.030 17.950 89.200 ;
        RECT 18.140 89.030 18.310 89.200 ;
        RECT 18.580 89.030 18.750 89.200 ;
        RECT 20.760 88.980 20.930 89.150 ;
        RECT 21.120 88.980 21.290 89.150 ;
        RECT 22.580 89.030 22.750 89.200 ;
        RECT 22.940 89.030 23.110 89.200 ;
        RECT 23.380 89.030 23.550 89.200 ;
        RECT 24.120 88.980 24.290 89.150 ;
        RECT 24.480 88.980 24.650 89.150 ;
        RECT 25.940 89.030 26.110 89.200 ;
        RECT 26.300 89.030 26.470 89.200 ;
        RECT 26.740 89.030 26.910 89.200 ;
        RECT 28.100 88.980 28.270 89.150 ;
        RECT 28.460 88.980 28.630 89.150 ;
        RECT 30.260 89.030 30.430 89.200 ;
        RECT 30.620 89.030 30.790 89.200 ;
        RECT 31.060 89.030 31.230 89.200 ;
        RECT 31.800 88.980 31.970 89.150 ;
        RECT 32.160 88.980 32.330 89.150 ;
        RECT 32.520 88.980 32.690 89.150 ;
        RECT 33.360 88.980 33.530 89.150 ;
        RECT 33.720 88.980 33.890 89.150 ;
        RECT 34.080 88.980 34.250 89.150 ;
        RECT 35.000 88.980 35.170 89.150 ;
        RECT 35.360 88.980 35.530 89.150 ;
        RECT 35.720 88.980 35.890 89.150 ;
        RECT 36.980 89.030 37.150 89.200 ;
        RECT 37.340 89.030 37.510 89.200 ;
        RECT 37.780 89.030 37.950 89.200 ;
        RECT 38.520 88.980 38.690 89.150 ;
        RECT 38.880 88.980 39.050 89.150 ;
        RECT 39.240 88.980 39.410 89.150 ;
        RECT 40.080 88.980 40.250 89.150 ;
        RECT 40.440 88.980 40.610 89.150 ;
        RECT 40.800 88.980 40.970 89.150 ;
        RECT 41.720 88.980 41.890 89.150 ;
        RECT 42.080 88.980 42.250 89.150 ;
        RECT 42.440 88.980 42.610 89.150 ;
        RECT 43.700 89.030 43.870 89.200 ;
        RECT 44.060 89.030 44.230 89.200 ;
        RECT 44.500 89.030 44.670 89.200 ;
        RECT 45.240 88.980 45.410 89.150 ;
        RECT 45.600 88.980 45.770 89.150 ;
        RECT 45.960 88.980 46.130 89.150 ;
        RECT 46.800 88.980 46.970 89.150 ;
        RECT 47.160 88.980 47.330 89.150 ;
        RECT 47.520 88.980 47.690 89.150 ;
        RECT 48.440 88.980 48.610 89.150 ;
        RECT 48.800 88.980 48.970 89.150 ;
        RECT 49.160 88.980 49.330 89.150 ;
        RECT 50.420 89.030 50.590 89.200 ;
        RECT 50.780 89.030 50.950 89.200 ;
        RECT 51.220 89.030 51.390 89.200 ;
        RECT 51.940 88.980 52.110 89.150 ;
        RECT 52.300 88.980 52.470 89.150 ;
        RECT 52.660 88.980 52.830 89.150 ;
        RECT 53.020 88.980 53.190 89.150 ;
        RECT 54.180 88.980 54.350 89.150 ;
        RECT 54.540 88.980 54.710 89.150 ;
        RECT 54.900 88.980 55.070 89.150 ;
        RECT 55.260 88.980 55.430 89.150 ;
        RECT 56.180 89.030 56.350 89.200 ;
        RECT 56.540 89.030 56.710 89.200 ;
        RECT 56.980 89.030 57.150 89.200 ;
        RECT 58.380 88.980 58.550 89.150 ;
        RECT 58.740 88.980 58.910 89.150 ;
        RECT 59.100 88.980 59.270 89.150 ;
        RECT 59.460 88.980 59.630 89.150 ;
        RECT 60.570 88.980 60.740 89.150 ;
        RECT 60.930 88.980 61.100 89.150 ;
        RECT 61.290 88.980 61.460 89.150 ;
        RECT 61.650 88.980 61.820 89.150 ;
        RECT 62.420 89.030 62.590 89.200 ;
        RECT 62.780 89.030 62.950 89.200 ;
        RECT 63.220 89.030 63.390 89.200 ;
        RECT 64.580 88.980 64.750 89.150 ;
        RECT 64.940 88.980 65.110 89.150 ;
        RECT 66.740 89.030 66.910 89.200 ;
        RECT 67.100 89.030 67.270 89.200 ;
        RECT 67.540 89.030 67.710 89.200 ;
        RECT 68.760 88.980 68.930 89.150 ;
        RECT 69.120 88.980 69.290 89.150 ;
        RECT 70.580 89.030 70.750 89.200 ;
        RECT 70.940 89.030 71.110 89.200 ;
        RECT 71.380 89.030 71.550 89.200 ;
        RECT 72.110 88.980 72.280 89.150 ;
        RECT 72.470 88.980 72.640 89.150 ;
        RECT 72.830 88.980 73.000 89.150 ;
        RECT 73.550 88.980 73.720 89.150 ;
        RECT 73.910 88.980 74.080 89.150 ;
        RECT 74.270 88.980 74.440 89.150 ;
        RECT 74.630 88.980 74.800 89.150 ;
        RECT 75.860 89.030 76.030 89.200 ;
        RECT 76.220 89.030 76.390 89.200 ;
        RECT 76.660 89.030 76.830 89.200 ;
        RECT 77.400 88.980 77.570 89.150 ;
        RECT 77.760 88.980 77.930 89.150 ;
        RECT 78.120 88.980 78.290 89.150 ;
        RECT 78.960 88.980 79.130 89.150 ;
        RECT 79.320 88.980 79.490 89.150 ;
        RECT 79.680 88.980 79.850 89.150 ;
        RECT 80.600 88.980 80.770 89.150 ;
        RECT 80.960 88.980 81.130 89.150 ;
        RECT 81.320 88.980 81.490 89.150 ;
        RECT 82.580 89.030 82.750 89.200 ;
        RECT 82.940 89.030 83.110 89.200 ;
        RECT 83.380 89.030 83.550 89.200 ;
        RECT 84.120 88.980 84.290 89.150 ;
        RECT 84.480 88.980 84.650 89.150 ;
        RECT 84.840 88.980 85.010 89.150 ;
        RECT 85.680 88.980 85.850 89.150 ;
        RECT 86.040 88.980 86.210 89.150 ;
        RECT 86.400 88.980 86.570 89.150 ;
        RECT 87.320 88.980 87.490 89.150 ;
        RECT 87.680 88.980 87.850 89.150 ;
        RECT 88.040 88.980 88.210 89.150 ;
        RECT 89.510 89.030 89.680 89.200 ;
        RECT 89.950 89.030 90.120 89.200 ;
        RECT 90.360 89.030 90.530 89.200 ;
        RECT 90.790 89.030 90.960 89.200 ;
        RECT 91.230 89.030 91.400 89.200 ;
        RECT 91.640 89.030 91.810 89.200 ;
        RECT 93.720 88.980 93.890 89.150 ;
        RECT 94.080 88.980 94.250 89.150 ;
        RECT 94.440 88.980 94.610 89.150 ;
        RECT 95.280 88.980 95.450 89.150 ;
        RECT 95.640 88.980 95.810 89.150 ;
        RECT 96.000 88.980 96.170 89.150 ;
        RECT 96.920 88.980 97.090 89.150 ;
        RECT 97.280 88.980 97.450 89.150 ;
        RECT 97.640 88.980 97.810 89.150 ;
        RECT 98.900 89.030 99.070 89.200 ;
        RECT 99.260 89.030 99.430 89.200 ;
        RECT 99.700 89.030 99.870 89.200 ;
        RECT 102.460 88.980 102.630 89.150 ;
        RECT 102.820 88.980 102.990 89.150 ;
        RECT 105.200 88.980 105.370 89.150 ;
        RECT 105.560 88.980 105.730 89.150 ;
        RECT 105.920 88.980 106.090 89.150 ;
        RECT 106.280 88.980 106.450 89.150 ;
        RECT 107.540 89.030 107.710 89.200 ;
        RECT 107.900 89.030 108.070 89.200 ;
        RECT 108.340 89.030 108.510 89.200 ;
        RECT 109.080 88.980 109.250 89.150 ;
        RECT 109.440 88.980 109.610 89.150 ;
        RECT 109.800 88.980 109.970 89.150 ;
        RECT 110.160 88.980 110.330 89.150 ;
        RECT 110.520 88.980 110.690 89.150 ;
        RECT 111.860 89.030 112.030 89.200 ;
        RECT 112.220 89.030 112.390 89.200 ;
        RECT 112.660 89.030 112.830 89.200 ;
        RECT 114.020 88.980 114.190 89.150 ;
        RECT 114.380 88.980 114.550 89.150 ;
        RECT 116.180 89.030 116.350 89.200 ;
        RECT 116.540 89.030 116.710 89.200 ;
        RECT 116.980 89.030 117.150 89.200 ;
        RECT 118.820 88.980 118.990 89.150 ;
        RECT 119.180 88.980 119.350 89.150 ;
        RECT 121.190 89.030 121.360 89.200 ;
        RECT 121.630 89.030 121.800 89.200 ;
        RECT 122.040 89.030 122.210 89.200 ;
        RECT 122.470 89.030 122.640 89.200 ;
        RECT 122.910 89.030 123.080 89.200 ;
        RECT 123.320 89.030 123.490 89.200 ;
        RECT 125.030 89.030 125.200 89.200 ;
        RECT 125.470 89.030 125.640 89.200 ;
        RECT 125.880 89.030 126.050 89.200 ;
        RECT 126.310 89.030 126.480 89.200 ;
        RECT 126.750 89.030 126.920 89.200 ;
        RECT 127.160 89.030 127.330 89.200 ;
        RECT 128.870 89.030 129.040 89.200 ;
        RECT 129.310 89.030 129.480 89.200 ;
        RECT 129.720 89.030 129.890 89.200 ;
        RECT 130.150 89.030 130.320 89.200 ;
        RECT 130.590 89.030 130.760 89.200 ;
        RECT 131.000 89.030 131.170 89.200 ;
        RECT 132.500 89.030 132.670 89.200 ;
        RECT 132.860 89.030 133.030 89.200 ;
        RECT 133.300 89.030 133.470 89.200 ;
        RECT 134.680 88.980 134.850 89.150 ;
        RECT 135.040 88.980 135.210 89.150 ;
        RECT 137.510 89.030 137.680 89.200 ;
        RECT 137.950 89.030 138.120 89.200 ;
        RECT 138.360 89.030 138.530 89.200 ;
        RECT 138.790 89.030 138.960 89.200 ;
        RECT 139.230 89.030 139.400 89.200 ;
        RECT 139.640 89.030 139.810 89.200 ;
        RECT 6.260 81.740 6.430 81.910 ;
        RECT 6.620 81.740 6.790 81.910 ;
        RECT 7.060 81.740 7.230 81.910 ;
        RECT 8.340 81.790 8.510 81.960 ;
        RECT 8.700 81.790 8.870 81.960 ;
        RECT 10.730 81.790 10.900 81.960 ;
        RECT 13.160 81.790 13.330 81.960 ;
        RECT 13.520 81.790 13.690 81.960 ;
        RECT 13.880 81.790 14.050 81.960 ;
        RECT 15.500 81.790 15.670 81.960 ;
        RECT 15.860 81.790 16.030 81.960 ;
        RECT 16.220 81.790 16.390 81.960 ;
        RECT 18.200 81.790 18.370 81.960 ;
        RECT 18.560 81.790 18.730 81.960 ;
        RECT 18.920 81.790 19.090 81.960 ;
        RECT 19.950 81.790 20.120 81.960 ;
        RECT 20.310 81.790 20.480 81.960 ;
        RECT 20.670 81.790 20.840 81.960 ;
        RECT 21.480 81.790 21.650 81.960 ;
        RECT 21.840 81.790 22.010 81.960 ;
        RECT 22.200 81.790 22.370 81.960 ;
        RECT 23.540 81.740 23.710 81.910 ;
        RECT 23.900 81.740 24.070 81.910 ;
        RECT 24.340 81.740 24.510 81.910 ;
        RECT 25.700 81.790 25.870 81.960 ;
        RECT 26.060 81.790 26.230 81.960 ;
        RECT 27.860 81.740 28.030 81.910 ;
        RECT 28.220 81.740 28.390 81.910 ;
        RECT 28.660 81.740 28.830 81.910 ;
        RECT 29.380 81.790 29.550 81.960 ;
        RECT 29.740 81.790 29.910 81.960 ;
        RECT 30.100 81.790 30.270 81.960 ;
        RECT 30.460 81.790 30.630 81.960 ;
        RECT 31.620 81.790 31.790 81.960 ;
        RECT 31.980 81.790 32.150 81.960 ;
        RECT 32.340 81.790 32.510 81.960 ;
        RECT 32.700 81.790 32.870 81.960 ;
        RECT 33.620 81.740 33.790 81.910 ;
        RECT 33.980 81.740 34.150 81.910 ;
        RECT 34.420 81.740 34.590 81.910 ;
        RECT 35.780 81.790 35.950 81.960 ;
        RECT 36.140 81.790 36.310 81.960 ;
        RECT 37.940 81.740 38.110 81.910 ;
        RECT 38.300 81.740 38.470 81.910 ;
        RECT 38.740 81.740 38.910 81.910 ;
        RECT 39.480 81.790 39.650 81.960 ;
        RECT 39.840 81.790 40.010 81.960 ;
        RECT 40.200 81.790 40.370 81.960 ;
        RECT 41.040 81.790 41.210 81.960 ;
        RECT 41.400 81.790 41.570 81.960 ;
        RECT 41.760 81.790 41.930 81.960 ;
        RECT 42.680 81.790 42.850 81.960 ;
        RECT 43.040 81.790 43.210 81.960 ;
        RECT 43.400 81.790 43.570 81.960 ;
        RECT 44.870 81.740 45.040 81.910 ;
        RECT 45.310 81.740 45.480 81.910 ;
        RECT 45.720 81.740 45.890 81.910 ;
        RECT 46.150 81.740 46.320 81.910 ;
        RECT 46.590 81.740 46.760 81.910 ;
        RECT 47.000 81.740 47.170 81.910 ;
        RECT 49.080 81.790 49.250 81.960 ;
        RECT 49.440 81.790 49.610 81.960 ;
        RECT 49.800 81.790 49.970 81.960 ;
        RECT 50.640 81.790 50.810 81.960 ;
        RECT 51.000 81.790 51.170 81.960 ;
        RECT 51.360 81.790 51.530 81.960 ;
        RECT 52.280 81.790 52.450 81.960 ;
        RECT 52.640 81.790 52.810 81.960 ;
        RECT 53.000 81.790 53.170 81.960 ;
        RECT 54.260 81.740 54.430 81.910 ;
        RECT 54.620 81.740 54.790 81.910 ;
        RECT 55.060 81.740 55.230 81.910 ;
        RECT 55.800 81.790 55.970 81.960 ;
        RECT 56.160 81.790 56.330 81.960 ;
        RECT 56.520 81.790 56.690 81.960 ;
        RECT 57.360 81.790 57.530 81.960 ;
        RECT 57.720 81.790 57.890 81.960 ;
        RECT 58.080 81.790 58.250 81.960 ;
        RECT 59.000 81.790 59.170 81.960 ;
        RECT 59.360 81.790 59.530 81.960 ;
        RECT 59.720 81.790 59.890 81.960 ;
        RECT 61.190 81.740 61.360 81.910 ;
        RECT 61.630 81.740 61.800 81.910 ;
        RECT 62.040 81.740 62.210 81.910 ;
        RECT 62.470 81.740 62.640 81.910 ;
        RECT 62.910 81.740 63.080 81.910 ;
        RECT 63.320 81.740 63.490 81.910 ;
        RECT 65.540 81.790 65.710 81.960 ;
        RECT 65.900 81.790 66.070 81.960 ;
        RECT 67.910 81.740 68.080 81.910 ;
        RECT 68.350 81.740 68.520 81.910 ;
        RECT 68.760 81.740 68.930 81.910 ;
        RECT 69.190 81.740 69.360 81.910 ;
        RECT 69.630 81.740 69.800 81.910 ;
        RECT 70.040 81.740 70.210 81.910 ;
        RECT 72.120 81.790 72.290 81.960 ;
        RECT 72.480 81.790 72.650 81.960 ;
        RECT 72.840 81.790 73.010 81.960 ;
        RECT 73.690 81.790 73.860 81.960 ;
        RECT 74.050 81.790 74.220 81.960 ;
        RECT 74.900 81.740 75.070 81.910 ;
        RECT 75.260 81.740 75.430 81.910 ;
        RECT 75.700 81.740 75.870 81.910 ;
        RECT 77.990 81.790 78.160 81.960 ;
        RECT 78.350 81.790 78.520 81.960 ;
        RECT 78.710 81.790 78.880 81.960 ;
        RECT 79.070 81.790 79.240 81.960 ;
        RECT 79.430 81.790 79.600 81.960 ;
        RECT 80.660 81.740 80.830 81.910 ;
        RECT 81.020 81.740 81.190 81.910 ;
        RECT 81.460 81.740 81.630 81.910 ;
        RECT 84.250 81.790 84.420 81.960 ;
        RECT 84.610 81.790 84.780 81.960 ;
        RECT 84.970 81.790 85.140 81.960 ;
        RECT 86.420 81.740 86.590 81.910 ;
        RECT 86.780 81.740 86.950 81.910 ;
        RECT 87.220 81.740 87.390 81.910 ;
        RECT 87.960 81.790 88.130 81.960 ;
        RECT 88.320 81.790 88.490 81.960 ;
        RECT 88.680 81.790 88.850 81.960 ;
        RECT 89.520 81.790 89.690 81.960 ;
        RECT 89.880 81.790 90.050 81.960 ;
        RECT 90.240 81.790 90.410 81.960 ;
        RECT 91.160 81.790 91.330 81.960 ;
        RECT 91.520 81.790 91.690 81.960 ;
        RECT 91.880 81.790 92.050 81.960 ;
        RECT 93.140 81.740 93.310 81.910 ;
        RECT 93.500 81.740 93.670 81.910 ;
        RECT 93.940 81.740 94.110 81.910 ;
        RECT 94.680 81.790 94.850 81.960 ;
        RECT 95.040 81.790 95.210 81.960 ;
        RECT 95.400 81.790 95.570 81.960 ;
        RECT 96.240 81.790 96.410 81.960 ;
        RECT 96.600 81.790 96.770 81.960 ;
        RECT 96.960 81.790 97.130 81.960 ;
        RECT 97.880 81.790 98.050 81.960 ;
        RECT 98.240 81.790 98.410 81.960 ;
        RECT 98.600 81.790 98.770 81.960 ;
        RECT 99.860 81.740 100.030 81.910 ;
        RECT 100.220 81.740 100.390 81.910 ;
        RECT 100.660 81.740 100.830 81.910 ;
        RECT 101.400 81.790 101.570 81.960 ;
        RECT 101.760 81.790 101.930 81.960 ;
        RECT 103.220 81.740 103.390 81.910 ;
        RECT 103.580 81.740 103.750 81.910 ;
        RECT 104.020 81.740 104.190 81.910 ;
        RECT 105.780 81.790 105.950 81.960 ;
        RECT 106.140 81.790 106.310 81.960 ;
        RECT 108.170 81.790 108.340 81.960 ;
        RECT 110.600 81.790 110.770 81.960 ;
        RECT 110.960 81.790 111.130 81.960 ;
        RECT 111.320 81.790 111.490 81.960 ;
        RECT 112.940 81.790 113.110 81.960 ;
        RECT 113.300 81.790 113.470 81.960 ;
        RECT 113.660 81.790 113.830 81.960 ;
        RECT 115.640 81.790 115.810 81.960 ;
        RECT 116.000 81.790 116.170 81.960 ;
        RECT 116.360 81.790 116.530 81.960 ;
        RECT 117.390 81.790 117.560 81.960 ;
        RECT 117.750 81.790 117.920 81.960 ;
        RECT 118.110 81.790 118.280 81.960 ;
        RECT 118.920 81.790 119.090 81.960 ;
        RECT 119.280 81.790 119.450 81.960 ;
        RECT 119.640 81.790 119.810 81.960 ;
        RECT 121.190 81.740 121.360 81.910 ;
        RECT 121.630 81.740 121.800 81.910 ;
        RECT 122.040 81.740 122.210 81.910 ;
        RECT 122.470 81.740 122.640 81.910 ;
        RECT 122.910 81.740 123.080 81.910 ;
        RECT 123.320 81.740 123.490 81.910 ;
        RECT 125.030 81.740 125.200 81.910 ;
        RECT 125.470 81.740 125.640 81.910 ;
        RECT 125.880 81.740 126.050 81.910 ;
        RECT 126.310 81.740 126.480 81.910 ;
        RECT 126.750 81.740 126.920 81.910 ;
        RECT 127.160 81.740 127.330 81.910 ;
        RECT 128.870 81.740 129.040 81.910 ;
        RECT 129.310 81.740 129.480 81.910 ;
        RECT 129.720 81.740 129.890 81.910 ;
        RECT 130.150 81.740 130.320 81.910 ;
        RECT 130.590 81.740 130.760 81.910 ;
        RECT 131.000 81.740 131.170 81.910 ;
        RECT 132.710 81.740 132.880 81.910 ;
        RECT 133.150 81.740 133.320 81.910 ;
        RECT 133.560 81.740 133.730 81.910 ;
        RECT 133.990 81.740 134.160 81.910 ;
        RECT 134.430 81.740 134.600 81.910 ;
        RECT 134.840 81.740 135.010 81.910 ;
        RECT 136.550 81.740 136.720 81.910 ;
        RECT 136.990 81.740 137.160 81.910 ;
        RECT 137.400 81.740 137.570 81.910 ;
        RECT 137.830 81.740 138.000 81.910 ;
        RECT 138.270 81.740 138.440 81.910 ;
        RECT 138.680 81.740 138.850 81.910 ;
        RECT 140.180 81.740 140.350 81.910 ;
        RECT 140.540 81.740 140.710 81.910 ;
        RECT 140.980 81.740 141.150 81.910 ;
        RECT 5.920 81.310 6.090 81.490 ;
        RECT 6.400 81.310 6.570 81.490 ;
        RECT 6.880 81.310 7.050 81.490 ;
        RECT 7.360 81.310 7.530 81.490 ;
        RECT 7.840 81.310 8.010 81.490 ;
        RECT 8.320 81.310 8.490 81.490 ;
        RECT 8.800 81.310 8.970 81.490 ;
        RECT 9.280 81.310 9.450 81.490 ;
        RECT 9.760 81.310 9.930 81.490 ;
        RECT 10.240 81.310 10.410 81.490 ;
        RECT 10.720 81.310 10.890 81.490 ;
        RECT 11.200 81.310 11.370 81.490 ;
        RECT 11.680 81.310 11.850 81.490 ;
        RECT 12.160 81.310 12.330 81.490 ;
        RECT 12.640 81.310 12.810 81.490 ;
        RECT 13.120 81.310 13.290 81.490 ;
        RECT 13.600 81.310 13.770 81.490 ;
        RECT 14.080 81.310 14.250 81.490 ;
      LAYER li1 ;
        RECT 14.400 81.480 14.880 81.490 ;
      LAYER li1 ;
        RECT 14.560 81.310 14.730 81.480 ;
        RECT 15.040 81.310 15.210 81.490 ;
        RECT 15.520 81.310 15.690 81.490 ;
        RECT 16.000 81.310 16.170 81.490 ;
        RECT 16.480 81.310 16.650 81.490 ;
        RECT 16.960 81.310 17.130 81.490 ;
        RECT 17.440 81.310 17.610 81.490 ;
        RECT 17.920 81.310 18.090 81.490 ;
        RECT 18.400 81.310 18.570 81.490 ;
        RECT 18.880 81.310 19.050 81.490 ;
        RECT 19.360 81.310 19.530 81.490 ;
        RECT 19.840 81.310 20.010 81.490 ;
        RECT 20.320 81.310 20.490 81.490 ;
        RECT 20.800 81.310 20.970 81.490 ;
        RECT 21.280 81.310 21.450 81.490 ;
        RECT 21.760 81.310 21.930 81.490 ;
        RECT 22.240 81.310 22.410 81.490 ;
        RECT 22.720 81.310 22.890 81.490 ;
        RECT 23.200 81.310 23.370 81.490 ;
        RECT 23.680 81.310 23.850 81.490 ;
        RECT 24.160 81.310 24.330 81.490 ;
        RECT 24.640 81.310 24.810 81.490 ;
        RECT 25.120 81.310 25.290 81.490 ;
        RECT 25.600 81.310 25.770 81.490 ;
        RECT 26.080 81.310 26.250 81.490 ;
        RECT 26.560 81.310 26.730 81.490 ;
        RECT 27.040 81.310 27.210 81.490 ;
        RECT 27.520 81.310 27.690 81.490 ;
        RECT 28.000 81.310 28.170 81.490 ;
        RECT 28.480 81.310 28.650 81.490 ;
        RECT 28.960 81.310 29.130 81.490 ;
        RECT 29.440 81.310 29.610 81.490 ;
        RECT 29.920 81.310 30.090 81.490 ;
        RECT 30.400 81.310 30.570 81.490 ;
        RECT 30.880 81.310 31.050 81.490 ;
        RECT 31.360 81.310 31.530 81.490 ;
        RECT 31.840 81.310 32.010 81.490 ;
        RECT 32.320 81.310 32.490 81.490 ;
        RECT 32.800 81.310 32.970 81.490 ;
        RECT 33.280 81.310 33.450 81.490 ;
        RECT 33.760 81.310 33.930 81.490 ;
        RECT 34.240 81.310 34.410 81.490 ;
        RECT 34.720 81.310 34.890 81.490 ;
        RECT 35.200 81.310 35.370 81.490 ;
        RECT 35.680 81.310 35.850 81.490 ;
        RECT 36.160 81.310 36.330 81.490 ;
        RECT 36.640 81.310 36.810 81.490 ;
        RECT 37.120 81.310 37.290 81.490 ;
        RECT 37.600 81.310 37.770 81.490 ;
        RECT 38.080 81.310 38.250 81.490 ;
        RECT 38.560 81.310 38.730 81.490 ;
        RECT 39.040 81.310 39.210 81.490 ;
        RECT 39.520 81.310 39.690 81.490 ;
        RECT 40.000 81.310 40.170 81.490 ;
        RECT 40.480 81.310 40.650 81.490 ;
        RECT 40.960 81.310 41.130 81.490 ;
        RECT 41.440 81.310 41.610 81.490 ;
        RECT 41.920 81.310 42.090 81.490 ;
        RECT 42.400 81.310 42.570 81.490 ;
        RECT 42.880 81.310 43.050 81.490 ;
        RECT 43.360 81.310 43.530 81.490 ;
        RECT 43.840 81.310 44.010 81.490 ;
        RECT 44.320 81.310 44.490 81.490 ;
        RECT 44.800 81.310 44.970 81.490 ;
        RECT 45.280 81.310 45.450 81.490 ;
        RECT 45.760 81.310 45.930 81.490 ;
        RECT 46.240 81.310 46.410 81.490 ;
        RECT 46.720 81.310 46.890 81.490 ;
        RECT 47.200 81.310 47.370 81.490 ;
        RECT 47.680 81.310 47.850 81.490 ;
        RECT 48.160 81.310 48.330 81.490 ;
        RECT 48.640 81.310 48.810 81.490 ;
        RECT 49.120 81.310 49.290 81.490 ;
        RECT 49.600 81.310 49.770 81.490 ;
        RECT 50.080 81.310 50.250 81.490 ;
        RECT 50.560 81.310 50.730 81.490 ;
        RECT 51.040 81.310 51.210 81.490 ;
        RECT 51.520 81.310 51.690 81.490 ;
        RECT 52.000 81.310 52.170 81.490 ;
        RECT 52.480 81.310 52.650 81.490 ;
        RECT 52.960 81.310 53.130 81.490 ;
        RECT 53.440 81.310 53.610 81.490 ;
        RECT 53.920 81.310 54.090 81.490 ;
        RECT 54.400 81.310 54.570 81.490 ;
        RECT 54.880 81.310 55.050 81.490 ;
        RECT 55.360 81.310 55.530 81.490 ;
        RECT 55.840 81.310 56.010 81.490 ;
        RECT 56.320 81.310 56.490 81.490 ;
        RECT 56.800 81.310 56.970 81.490 ;
        RECT 57.280 81.310 57.450 81.490 ;
        RECT 57.760 81.310 57.930 81.490 ;
        RECT 58.240 81.310 58.410 81.490 ;
        RECT 58.720 81.310 58.890 81.490 ;
        RECT 59.200 81.310 59.370 81.490 ;
        RECT 59.680 81.310 59.850 81.490 ;
        RECT 60.160 81.310 60.330 81.490 ;
        RECT 60.640 81.310 60.810 81.490 ;
        RECT 61.120 81.310 61.290 81.490 ;
        RECT 61.600 81.310 61.770 81.490 ;
        RECT 62.080 81.310 62.250 81.490 ;
        RECT 62.560 81.310 62.730 81.490 ;
        RECT 63.040 81.310 63.210 81.490 ;
        RECT 63.520 81.310 63.690 81.490 ;
        RECT 64.000 81.310 64.170 81.490 ;
        RECT 64.480 81.480 64.650 81.490 ;
      LAYER li1 ;
        RECT 64.320 81.310 64.800 81.480 ;
      LAYER li1 ;
        RECT 64.960 81.310 65.130 81.490 ;
        RECT 65.440 81.310 65.610 81.490 ;
        RECT 65.920 81.310 66.090 81.490 ;
        RECT 66.400 81.310 66.570 81.490 ;
        RECT 66.880 81.310 67.050 81.490 ;
        RECT 67.360 81.310 67.530 81.490 ;
        RECT 67.840 81.310 68.010 81.490 ;
        RECT 68.320 81.310 68.490 81.490 ;
        RECT 68.800 81.310 68.970 81.490 ;
        RECT 69.280 81.310 69.450 81.490 ;
        RECT 69.760 81.310 69.930 81.490 ;
        RECT 70.240 81.310 70.410 81.490 ;
        RECT 70.720 81.310 70.890 81.490 ;
      LAYER li1 ;
        RECT 71.040 81.480 71.520 81.490 ;
      LAYER li1 ;
        RECT 71.200 81.310 71.370 81.480 ;
        RECT 71.680 81.310 71.850 81.490 ;
        RECT 72.160 81.310 72.330 81.490 ;
        RECT 72.640 81.310 72.810 81.490 ;
        RECT 73.120 81.310 73.290 81.490 ;
        RECT 73.600 81.310 73.770 81.490 ;
        RECT 74.080 81.310 74.250 81.490 ;
        RECT 74.560 81.310 74.730 81.490 ;
        RECT 75.040 81.310 75.210 81.490 ;
        RECT 75.520 81.310 75.690 81.490 ;
        RECT 76.000 81.310 76.170 81.490 ;
        RECT 76.480 81.310 76.650 81.490 ;
        RECT 76.960 81.310 77.130 81.490 ;
        RECT 77.440 81.310 77.610 81.490 ;
        RECT 77.920 81.310 78.090 81.490 ;
        RECT 78.400 81.310 78.570 81.490 ;
        RECT 78.880 81.310 79.050 81.490 ;
        RECT 79.360 81.310 79.530 81.490 ;
        RECT 79.840 81.310 80.010 81.490 ;
        RECT 80.320 81.310 80.490 81.490 ;
      LAYER li1 ;
        RECT 80.640 81.480 81.120 81.490 ;
      LAYER li1 ;
        RECT 80.800 81.310 80.970 81.480 ;
        RECT 81.280 81.310 81.450 81.490 ;
        RECT 81.760 81.310 81.930 81.490 ;
        RECT 82.240 81.310 82.410 81.490 ;
        RECT 82.720 81.310 82.890 81.490 ;
        RECT 83.200 81.310 83.370 81.490 ;
        RECT 83.680 81.310 83.850 81.490 ;
        RECT 84.160 81.310 84.330 81.490 ;
        RECT 84.640 81.310 84.810 81.490 ;
        RECT 85.120 81.310 85.290 81.490 ;
        RECT 85.600 81.310 85.770 81.490 ;
        RECT 86.080 81.310 86.250 81.490 ;
        RECT 86.560 81.310 86.730 81.490 ;
        RECT 87.040 81.310 87.210 81.490 ;
        RECT 87.520 81.310 87.690 81.490 ;
        RECT 88.000 81.310 88.170 81.490 ;
        RECT 88.480 81.310 88.650 81.490 ;
        RECT 88.960 81.310 89.130 81.490 ;
        RECT 89.440 81.310 89.610 81.490 ;
        RECT 89.920 81.310 90.090 81.490 ;
        RECT 90.400 81.310 90.570 81.490 ;
        RECT 90.880 81.310 91.050 81.490 ;
        RECT 91.360 81.310 91.530 81.490 ;
        RECT 91.840 81.310 92.010 81.490 ;
        RECT 92.320 81.310 92.490 81.490 ;
        RECT 92.800 81.310 92.970 81.490 ;
        RECT 93.280 81.310 93.450 81.490 ;
        RECT 93.760 81.310 93.930 81.490 ;
        RECT 94.240 81.310 94.410 81.490 ;
        RECT 94.720 81.310 94.890 81.490 ;
        RECT 95.200 81.310 95.370 81.490 ;
        RECT 95.680 81.310 95.850 81.490 ;
        RECT 96.160 81.310 96.330 81.490 ;
        RECT 96.640 81.310 96.810 81.490 ;
        RECT 97.120 81.310 97.290 81.490 ;
        RECT 97.600 81.310 97.770 81.490 ;
        RECT 98.080 81.310 98.250 81.490 ;
        RECT 98.560 81.310 98.730 81.490 ;
        RECT 99.040 81.310 99.210 81.490 ;
        RECT 99.520 81.310 99.690 81.490 ;
        RECT 100.000 81.310 100.170 81.490 ;
        RECT 100.480 81.310 100.650 81.490 ;
        RECT 100.960 81.310 101.130 81.490 ;
        RECT 101.440 81.310 101.610 81.490 ;
        RECT 101.920 81.310 102.090 81.490 ;
        RECT 102.400 81.310 102.570 81.490 ;
        RECT 102.880 81.310 103.050 81.490 ;
        RECT 103.360 81.310 103.530 81.490 ;
        RECT 103.840 81.310 104.010 81.490 ;
        RECT 104.320 81.310 104.490 81.490 ;
        RECT 104.800 81.480 104.970 81.490 ;
      LAYER li1 ;
        RECT 104.640 81.310 105.120 81.480 ;
      LAYER li1 ;
        RECT 105.280 81.310 105.450 81.490 ;
        RECT 105.760 81.310 105.930 81.490 ;
        RECT 106.240 81.310 106.410 81.490 ;
        RECT 106.720 81.310 106.890 81.490 ;
        RECT 107.200 81.310 107.370 81.490 ;
        RECT 107.680 81.310 107.850 81.490 ;
        RECT 108.160 81.310 108.330 81.490 ;
        RECT 108.640 81.310 108.810 81.490 ;
        RECT 109.120 81.310 109.290 81.490 ;
        RECT 109.600 81.310 109.770 81.490 ;
        RECT 110.080 81.310 110.250 81.490 ;
        RECT 110.560 81.310 110.730 81.490 ;
        RECT 111.040 81.310 111.210 81.490 ;
        RECT 111.520 81.310 111.690 81.490 ;
        RECT 112.000 81.310 112.170 81.490 ;
        RECT 112.480 81.310 112.650 81.490 ;
        RECT 112.960 81.310 113.130 81.490 ;
        RECT 113.440 81.310 113.610 81.490 ;
        RECT 113.920 81.310 114.090 81.490 ;
        RECT 114.400 81.310 114.570 81.490 ;
        RECT 114.880 81.310 115.050 81.490 ;
        RECT 115.360 81.310 115.530 81.490 ;
        RECT 115.840 81.310 116.010 81.490 ;
        RECT 116.320 81.310 116.490 81.490 ;
        RECT 116.800 81.310 116.970 81.490 ;
        RECT 117.280 81.310 117.450 81.490 ;
        RECT 117.760 81.310 117.930 81.490 ;
        RECT 118.240 81.310 118.410 81.490 ;
        RECT 118.720 81.310 118.890 81.490 ;
        RECT 119.200 81.310 119.370 81.490 ;
        RECT 119.680 81.310 119.850 81.490 ;
        RECT 120.160 81.310 120.330 81.490 ;
        RECT 120.640 81.310 120.810 81.490 ;
        RECT 121.120 81.310 121.290 81.490 ;
        RECT 121.600 81.310 121.770 81.490 ;
        RECT 122.080 81.310 122.250 81.490 ;
        RECT 122.560 81.310 122.730 81.490 ;
        RECT 123.040 81.310 123.210 81.490 ;
        RECT 123.520 81.310 123.690 81.490 ;
        RECT 124.000 81.310 124.170 81.490 ;
        RECT 124.480 81.310 124.650 81.490 ;
        RECT 124.960 81.310 125.130 81.490 ;
        RECT 125.440 81.310 125.610 81.490 ;
        RECT 125.920 81.310 126.090 81.490 ;
        RECT 126.400 81.310 126.570 81.490 ;
        RECT 126.880 81.310 127.050 81.490 ;
        RECT 127.360 81.310 127.530 81.490 ;
        RECT 127.840 81.310 128.010 81.490 ;
        RECT 128.320 81.310 128.490 81.490 ;
        RECT 128.800 81.310 128.970 81.490 ;
        RECT 129.280 81.310 129.450 81.490 ;
        RECT 129.760 81.310 129.930 81.490 ;
        RECT 130.240 81.310 130.410 81.490 ;
        RECT 130.720 81.310 130.890 81.490 ;
        RECT 131.200 81.310 131.370 81.490 ;
        RECT 131.680 81.310 131.850 81.490 ;
        RECT 132.160 81.310 132.330 81.490 ;
        RECT 132.640 81.310 132.810 81.490 ;
        RECT 133.120 81.310 133.290 81.490 ;
        RECT 133.600 81.310 133.770 81.490 ;
        RECT 134.080 81.310 134.250 81.490 ;
        RECT 134.560 81.310 134.730 81.490 ;
        RECT 135.040 81.310 135.210 81.490 ;
        RECT 135.520 81.310 135.690 81.490 ;
        RECT 136.000 81.310 136.170 81.490 ;
        RECT 136.480 81.310 136.650 81.490 ;
        RECT 136.960 81.310 137.130 81.490 ;
        RECT 137.440 81.310 137.610 81.490 ;
        RECT 137.920 81.310 138.090 81.490 ;
        RECT 138.400 81.310 138.570 81.490 ;
        RECT 138.880 81.310 139.050 81.490 ;
        RECT 139.360 81.310 139.530 81.490 ;
        RECT 139.840 81.310 140.010 81.490 ;
        RECT 140.320 81.310 140.490 81.490 ;
        RECT 140.800 81.310 140.970 81.490 ;
        RECT 141.280 81.310 141.450 81.490 ;
        RECT 141.760 81.480 141.930 81.490 ;
      LAYER li1 ;
        RECT 141.600 81.310 142.080 81.480 ;
      LAYER li1 ;
        RECT 6.470 80.890 6.640 81.060 ;
        RECT 6.910 80.890 7.080 81.060 ;
        RECT 7.320 80.890 7.490 81.060 ;
        RECT 7.750 80.890 7.920 81.060 ;
        RECT 8.190 80.890 8.360 81.060 ;
        RECT 8.600 80.890 8.770 81.060 ;
        RECT 10.310 80.890 10.480 81.060 ;
        RECT 10.750 80.890 10.920 81.060 ;
        RECT 11.160 80.890 11.330 81.060 ;
        RECT 11.590 80.890 11.760 81.060 ;
        RECT 12.030 80.890 12.200 81.060 ;
        RECT 12.440 80.890 12.610 81.060 ;
        RECT 15.620 80.840 15.790 81.010 ;
        RECT 15.980 80.840 16.150 81.010 ;
        RECT 17.990 80.890 18.160 81.060 ;
        RECT 18.430 80.890 18.600 81.060 ;
        RECT 18.840 80.890 19.010 81.060 ;
        RECT 19.270 80.890 19.440 81.060 ;
        RECT 19.710 80.890 19.880 81.060 ;
        RECT 20.120 80.890 20.290 81.060 ;
        RECT 21.620 80.890 21.790 81.060 ;
        RECT 21.980 80.890 22.150 81.060 ;
        RECT 22.420 80.890 22.590 81.060 ;
        RECT 23.700 80.840 23.870 81.010 ;
        RECT 24.060 80.840 24.230 81.010 ;
        RECT 26.090 80.840 26.260 81.010 ;
        RECT 28.520 80.840 28.690 81.010 ;
        RECT 28.880 80.840 29.050 81.010 ;
        RECT 29.240 80.840 29.410 81.010 ;
        RECT 30.860 80.840 31.030 81.010 ;
        RECT 31.220 80.840 31.390 81.010 ;
        RECT 31.580 80.840 31.750 81.010 ;
        RECT 33.560 80.840 33.730 81.010 ;
        RECT 33.920 80.840 34.090 81.010 ;
        RECT 34.280 80.840 34.450 81.010 ;
        RECT 35.310 80.840 35.480 81.010 ;
        RECT 35.670 80.840 35.840 81.010 ;
        RECT 36.030 80.840 36.200 81.010 ;
        RECT 36.840 80.840 37.010 81.010 ;
        RECT 37.200 80.840 37.370 81.010 ;
        RECT 37.560 80.840 37.730 81.010 ;
        RECT 39.110 80.890 39.280 81.060 ;
        RECT 39.550 80.890 39.720 81.060 ;
        RECT 39.960 80.890 40.130 81.060 ;
        RECT 40.390 80.890 40.560 81.060 ;
        RECT 40.830 80.890 41.000 81.060 ;
        RECT 41.240 80.890 41.410 81.060 ;
        RECT 42.900 80.840 43.070 81.010 ;
        RECT 43.260 80.840 43.430 81.010 ;
        RECT 45.290 80.840 45.460 81.010 ;
        RECT 47.720 80.840 47.890 81.010 ;
        RECT 48.080 80.840 48.250 81.010 ;
        RECT 48.440 80.840 48.610 81.010 ;
        RECT 50.060 80.840 50.230 81.010 ;
        RECT 50.420 80.840 50.590 81.010 ;
        RECT 50.780 80.840 50.950 81.010 ;
        RECT 52.760 80.840 52.930 81.010 ;
        RECT 53.120 80.840 53.290 81.010 ;
        RECT 53.480 80.840 53.650 81.010 ;
        RECT 54.510 80.840 54.680 81.010 ;
        RECT 54.870 80.840 55.040 81.010 ;
        RECT 55.230 80.840 55.400 81.010 ;
        RECT 56.040 80.840 56.210 81.010 ;
        RECT 56.400 80.840 56.570 81.010 ;
        RECT 56.760 80.840 56.930 81.010 ;
        RECT 58.310 80.890 58.480 81.060 ;
        RECT 58.750 80.890 58.920 81.060 ;
        RECT 59.160 80.890 59.330 81.060 ;
        RECT 59.590 80.890 59.760 81.060 ;
        RECT 60.030 80.890 60.200 81.060 ;
        RECT 60.440 80.890 60.610 81.060 ;
        RECT 61.560 80.840 61.730 81.010 ;
        RECT 61.920 80.840 62.090 81.010 ;
        RECT 62.280 80.840 62.450 81.010 ;
        RECT 63.120 80.840 63.290 81.010 ;
        RECT 63.480 80.840 63.650 81.010 ;
        RECT 63.840 80.840 64.010 81.010 ;
        RECT 64.760 80.840 64.930 81.010 ;
        RECT 65.120 80.840 65.290 81.010 ;
        RECT 65.480 80.840 65.650 81.010 ;
        RECT 66.950 80.890 67.120 81.060 ;
        RECT 67.390 80.890 67.560 81.060 ;
        RECT 67.800 80.890 67.970 81.060 ;
        RECT 68.230 80.890 68.400 81.060 ;
        RECT 68.670 80.890 68.840 81.060 ;
        RECT 69.080 80.890 69.250 81.060 ;
        RECT 72.220 80.840 72.390 81.010 ;
        RECT 72.580 80.840 72.750 81.010 ;
        RECT 74.960 80.840 75.130 81.010 ;
        RECT 75.320 80.840 75.490 81.010 ;
        RECT 75.680 80.840 75.850 81.010 ;
        RECT 76.040 80.840 76.210 81.010 ;
        RECT 77.510 80.890 77.680 81.060 ;
        RECT 77.950 80.890 78.120 81.060 ;
        RECT 78.360 80.890 78.530 81.060 ;
        RECT 78.790 80.890 78.960 81.060 ;
        RECT 79.230 80.890 79.400 81.060 ;
        RECT 79.640 80.890 79.810 81.060 ;
        RECT 81.240 80.840 81.410 81.010 ;
        RECT 81.600 80.840 81.770 81.010 ;
        RECT 81.960 80.840 82.130 81.010 ;
        RECT 82.800 80.840 82.970 81.010 ;
        RECT 83.160 80.840 83.330 81.010 ;
        RECT 83.520 80.840 83.690 81.010 ;
        RECT 84.440 80.840 84.610 81.010 ;
        RECT 84.800 80.840 84.970 81.010 ;
        RECT 85.160 80.840 85.330 81.010 ;
        RECT 86.420 80.890 86.590 81.060 ;
        RECT 86.780 80.890 86.950 81.060 ;
        RECT 87.220 80.890 87.390 81.060 ;
        RECT 87.960 80.840 88.130 81.010 ;
        RECT 88.320 80.840 88.490 81.010 ;
        RECT 88.680 80.840 88.850 81.010 ;
        RECT 89.520 80.840 89.690 81.010 ;
        RECT 89.880 80.840 90.050 81.010 ;
        RECT 90.240 80.840 90.410 81.010 ;
        RECT 91.160 80.840 91.330 81.010 ;
        RECT 91.520 80.840 91.690 81.010 ;
        RECT 91.880 80.840 92.050 81.010 ;
        RECT 93.140 80.890 93.310 81.060 ;
        RECT 93.500 80.890 93.670 81.060 ;
        RECT 93.940 80.890 94.110 81.060 ;
        RECT 95.390 80.840 95.560 81.010 ;
        RECT 95.750 80.840 95.920 81.010 ;
        RECT 96.110 80.840 96.280 81.010 ;
        RECT 96.470 80.840 96.640 81.010 ;
        RECT 96.830 80.840 97.000 81.010 ;
        RECT 97.190 80.840 97.360 81.010 ;
        RECT 98.420 80.890 98.590 81.060 ;
        RECT 98.780 80.890 98.950 81.060 ;
        RECT 99.220 80.890 99.390 81.060 ;
        RECT 100.670 80.840 100.840 81.010 ;
        RECT 101.030 80.840 101.200 81.010 ;
        RECT 101.390 80.840 101.560 81.010 ;
        RECT 101.750 80.840 101.920 81.010 ;
        RECT 102.110 80.840 102.280 81.010 ;
        RECT 102.470 80.840 102.640 81.010 ;
        RECT 103.700 80.890 103.870 81.060 ;
        RECT 104.060 80.890 104.230 81.060 ;
        RECT 104.500 80.890 104.670 81.060 ;
        RECT 105.950 80.840 106.120 81.010 ;
        RECT 106.310 80.840 106.480 81.010 ;
        RECT 106.670 80.840 106.840 81.010 ;
        RECT 107.030 80.840 107.200 81.010 ;
        RECT 107.390 80.840 107.560 81.010 ;
        RECT 107.750 80.840 107.920 81.010 ;
        RECT 108.980 80.890 109.150 81.060 ;
        RECT 109.340 80.890 109.510 81.060 ;
        RECT 109.780 80.890 109.950 81.060 ;
        RECT 111.140 80.840 111.310 81.010 ;
        RECT 111.500 80.840 111.670 81.010 ;
        RECT 113.300 80.890 113.470 81.060 ;
        RECT 113.660 80.890 113.830 81.060 ;
        RECT 114.100 80.890 114.270 81.060 ;
        RECT 115.460 80.840 115.630 81.010 ;
        RECT 115.820 80.840 115.990 81.010 ;
        RECT 117.620 80.890 117.790 81.060 ;
        RECT 117.980 80.890 118.150 81.060 ;
        RECT 118.420 80.890 118.590 81.060 ;
        RECT 119.780 80.840 119.950 81.010 ;
        RECT 120.140 80.840 120.310 81.010 ;
        RECT 121.940 80.890 122.110 81.060 ;
        RECT 122.300 80.890 122.470 81.060 ;
        RECT 122.740 80.890 122.910 81.060 ;
        RECT 124.100 80.840 124.270 81.010 ;
        RECT 124.460 80.840 124.630 81.010 ;
        RECT 126.470 80.890 126.640 81.060 ;
        RECT 126.910 80.890 127.080 81.060 ;
        RECT 127.320 80.890 127.490 81.060 ;
        RECT 127.750 80.890 127.920 81.060 ;
        RECT 128.190 80.890 128.360 81.060 ;
        RECT 128.600 80.890 128.770 81.060 ;
        RECT 130.310 80.890 130.480 81.060 ;
        RECT 130.750 80.890 130.920 81.060 ;
        RECT 131.160 80.890 131.330 81.060 ;
        RECT 131.590 80.890 131.760 81.060 ;
        RECT 132.030 80.890 132.200 81.060 ;
        RECT 132.440 80.890 132.610 81.060 ;
        RECT 134.150 80.890 134.320 81.060 ;
        RECT 134.590 80.890 134.760 81.060 ;
        RECT 135.000 80.890 135.170 81.060 ;
        RECT 135.430 80.890 135.600 81.060 ;
        RECT 135.870 80.890 136.040 81.060 ;
        RECT 136.280 80.890 136.450 81.060 ;
        RECT 137.990 80.890 138.160 81.060 ;
        RECT 138.430 80.890 138.600 81.060 ;
        RECT 138.840 80.890 139.010 81.060 ;
        RECT 139.270 80.890 139.440 81.060 ;
        RECT 139.710 80.890 139.880 81.060 ;
        RECT 140.120 80.890 140.290 81.060 ;
        RECT 6.470 73.600 6.640 73.770 ;
        RECT 6.910 73.600 7.080 73.770 ;
        RECT 7.320 73.600 7.490 73.770 ;
        RECT 7.750 73.600 7.920 73.770 ;
        RECT 8.190 73.600 8.360 73.770 ;
        RECT 8.600 73.600 8.770 73.770 ;
        RECT 10.310 73.600 10.480 73.770 ;
        RECT 10.750 73.600 10.920 73.770 ;
        RECT 11.160 73.600 11.330 73.770 ;
        RECT 11.590 73.600 11.760 73.770 ;
        RECT 12.030 73.600 12.200 73.770 ;
        RECT 12.440 73.600 12.610 73.770 ;
        RECT 14.150 73.600 14.320 73.770 ;
        RECT 14.590 73.600 14.760 73.770 ;
        RECT 15.000 73.600 15.170 73.770 ;
        RECT 15.430 73.600 15.600 73.770 ;
        RECT 15.870 73.600 16.040 73.770 ;
        RECT 16.280 73.600 16.450 73.770 ;
        RECT 18.020 73.650 18.190 73.820 ;
        RECT 18.380 73.650 18.550 73.820 ;
        RECT 20.180 73.600 20.350 73.770 ;
        RECT 20.540 73.600 20.710 73.770 ;
        RECT 20.980 73.600 21.150 73.770 ;
        RECT 22.340 73.650 22.510 73.820 ;
        RECT 22.700 73.650 22.870 73.820 ;
        RECT 24.500 73.600 24.670 73.770 ;
        RECT 24.860 73.600 25.030 73.770 ;
        RECT 25.300 73.600 25.470 73.770 ;
        RECT 26.040 73.650 26.210 73.820 ;
        RECT 26.400 73.650 26.570 73.820 ;
        RECT 26.760 73.650 26.930 73.820 ;
        RECT 27.600 73.650 27.770 73.820 ;
        RECT 27.960 73.650 28.130 73.820 ;
        RECT 28.320 73.650 28.490 73.820 ;
        RECT 29.240 73.650 29.410 73.820 ;
        RECT 29.600 73.650 29.770 73.820 ;
        RECT 29.960 73.650 30.130 73.820 ;
        RECT 31.220 73.600 31.390 73.770 ;
        RECT 31.580 73.600 31.750 73.770 ;
        RECT 32.020 73.600 32.190 73.770 ;
        RECT 32.760 73.650 32.930 73.820 ;
        RECT 33.120 73.650 33.290 73.820 ;
        RECT 33.480 73.650 33.650 73.820 ;
        RECT 34.320 73.650 34.490 73.820 ;
        RECT 34.680 73.650 34.850 73.820 ;
        RECT 35.040 73.650 35.210 73.820 ;
        RECT 35.960 73.650 36.130 73.820 ;
        RECT 36.320 73.650 36.490 73.820 ;
        RECT 36.680 73.650 36.850 73.820 ;
        RECT 37.940 73.600 38.110 73.770 ;
        RECT 38.300 73.600 38.470 73.770 ;
        RECT 38.740 73.600 38.910 73.770 ;
        RECT 39.480 73.650 39.650 73.820 ;
        RECT 39.840 73.650 40.010 73.820 ;
        RECT 40.200 73.650 40.370 73.820 ;
        RECT 41.040 73.650 41.210 73.820 ;
        RECT 41.400 73.650 41.570 73.820 ;
        RECT 41.760 73.650 41.930 73.820 ;
        RECT 42.680 73.650 42.850 73.820 ;
        RECT 43.040 73.650 43.210 73.820 ;
        RECT 43.400 73.650 43.570 73.820 ;
        RECT 44.660 73.600 44.830 73.770 ;
        RECT 45.020 73.600 45.190 73.770 ;
        RECT 45.460 73.600 45.630 73.770 ;
        RECT 47.640 73.650 47.810 73.820 ;
        RECT 48.000 73.650 48.170 73.820 ;
        RECT 48.360 73.650 48.530 73.820 ;
        RECT 49.200 73.650 49.370 73.820 ;
        RECT 49.560 73.650 49.730 73.820 ;
        RECT 49.920 73.650 50.090 73.820 ;
        RECT 50.840 73.650 51.010 73.820 ;
        RECT 51.200 73.650 51.370 73.820 ;
        RECT 51.560 73.650 51.730 73.820 ;
        RECT 52.820 73.600 52.990 73.770 ;
        RECT 53.180 73.600 53.350 73.770 ;
        RECT 53.620 73.600 53.790 73.770 ;
        RECT 54.940 73.650 55.110 73.820 ;
        RECT 55.300 73.650 55.470 73.820 ;
        RECT 57.680 73.650 57.850 73.820 ;
        RECT 58.040 73.650 58.210 73.820 ;
        RECT 58.400 73.650 58.570 73.820 ;
        RECT 58.760 73.650 58.930 73.820 ;
        RECT 60.020 73.600 60.190 73.770 ;
        RECT 60.380 73.600 60.550 73.770 ;
        RECT 60.820 73.600 60.990 73.770 ;
        RECT 62.100 73.650 62.270 73.820 ;
        RECT 62.460 73.650 62.630 73.820 ;
        RECT 64.490 73.650 64.660 73.820 ;
        RECT 66.920 73.650 67.090 73.820 ;
        RECT 67.280 73.650 67.450 73.820 ;
        RECT 67.640 73.650 67.810 73.820 ;
        RECT 69.260 73.650 69.430 73.820 ;
        RECT 69.620 73.650 69.790 73.820 ;
        RECT 69.980 73.650 70.150 73.820 ;
        RECT 71.960 73.650 72.130 73.820 ;
        RECT 72.320 73.650 72.490 73.820 ;
        RECT 72.680 73.650 72.850 73.820 ;
        RECT 73.710 73.650 73.880 73.820 ;
        RECT 74.070 73.650 74.240 73.820 ;
        RECT 74.430 73.650 74.600 73.820 ;
        RECT 75.240 73.650 75.410 73.820 ;
        RECT 75.600 73.650 75.770 73.820 ;
        RECT 75.960 73.650 76.130 73.820 ;
        RECT 77.300 73.600 77.470 73.770 ;
        RECT 77.660 73.600 77.830 73.770 ;
        RECT 78.100 73.600 78.270 73.770 ;
        RECT 79.320 73.650 79.490 73.820 ;
        RECT 79.680 73.650 79.850 73.820 ;
        RECT 81.140 73.600 81.310 73.770 ;
        RECT 81.500 73.600 81.670 73.770 ;
        RECT 81.940 73.600 82.110 73.770 ;
        RECT 83.120 73.650 83.290 73.820 ;
        RECT 83.480 73.650 83.650 73.820 ;
        RECT 83.840 73.650 84.010 73.820 ;
        RECT 84.200 73.650 84.370 73.820 ;
        RECT 84.560 73.650 84.730 73.820 ;
        RECT 84.920 73.650 85.090 73.820 ;
        RECT 85.280 73.650 85.450 73.820 ;
        RECT 85.640 73.650 85.810 73.820 ;
        RECT 86.450 73.650 86.620 73.820 ;
        RECT 86.810 73.650 86.980 73.820 ;
        RECT 87.170 73.650 87.340 73.820 ;
        RECT 87.530 73.650 87.700 73.820 ;
        RECT 88.340 73.600 88.510 73.770 ;
        RECT 88.700 73.600 88.870 73.770 ;
        RECT 89.140 73.600 89.310 73.770 ;
        RECT 90.540 73.650 90.710 73.820 ;
        RECT 90.900 73.650 91.070 73.820 ;
        RECT 91.260 73.650 91.430 73.820 ;
        RECT 91.620 73.650 91.790 73.820 ;
        RECT 92.730 73.650 92.900 73.820 ;
        RECT 93.090 73.650 93.260 73.820 ;
        RECT 93.450 73.650 93.620 73.820 ;
        RECT 93.810 73.650 93.980 73.820 ;
        RECT 94.580 73.600 94.750 73.770 ;
        RECT 94.940 73.600 95.110 73.770 ;
        RECT 95.380 73.600 95.550 73.770 ;
        RECT 96.120 73.650 96.290 73.820 ;
        RECT 96.480 73.650 96.650 73.820 ;
        RECT 96.840 73.650 97.010 73.820 ;
        RECT 98.250 73.650 98.420 73.820 ;
        RECT 98.610 73.650 98.780 73.820 ;
        RECT 98.970 73.650 99.140 73.820 ;
        RECT 99.860 73.600 100.030 73.770 ;
        RECT 100.220 73.600 100.390 73.770 ;
        RECT 100.660 73.600 100.830 73.770 ;
        RECT 101.980 73.650 102.150 73.820 ;
        RECT 102.340 73.650 102.510 73.820 ;
        RECT 104.720 73.650 104.890 73.820 ;
        RECT 105.080 73.650 105.250 73.820 ;
        RECT 105.440 73.650 105.610 73.820 ;
        RECT 105.800 73.650 105.970 73.820 ;
        RECT 107.060 73.600 107.230 73.770 ;
        RECT 107.420 73.600 107.590 73.770 ;
        RECT 107.860 73.600 108.030 73.770 ;
        RECT 109.560 73.650 109.730 73.820 ;
        RECT 109.920 73.650 110.090 73.820 ;
        RECT 110.280 73.650 110.450 73.820 ;
        RECT 111.130 73.650 111.300 73.820 ;
        RECT 111.490 73.650 111.660 73.820 ;
        RECT 112.340 73.600 112.510 73.770 ;
        RECT 112.700 73.600 112.870 73.770 ;
        RECT 113.140 73.600 113.310 73.770 ;
        RECT 114.420 73.650 114.590 73.820 ;
        RECT 114.780 73.650 114.950 73.820 ;
        RECT 116.810 73.650 116.980 73.820 ;
        RECT 119.240 73.650 119.410 73.820 ;
        RECT 119.600 73.650 119.770 73.820 ;
        RECT 119.960 73.650 120.130 73.820 ;
        RECT 121.580 73.650 121.750 73.820 ;
        RECT 121.940 73.650 122.110 73.820 ;
        RECT 122.300 73.650 122.470 73.820 ;
        RECT 124.280 73.650 124.450 73.820 ;
        RECT 124.640 73.650 124.810 73.820 ;
        RECT 125.000 73.650 125.170 73.820 ;
        RECT 126.030 73.650 126.200 73.820 ;
        RECT 126.390 73.650 126.560 73.820 ;
        RECT 126.750 73.650 126.920 73.820 ;
        RECT 127.560 73.650 127.730 73.820 ;
        RECT 127.920 73.650 128.090 73.820 ;
        RECT 128.280 73.650 128.450 73.820 ;
        RECT 129.830 73.600 130.000 73.770 ;
        RECT 130.270 73.600 130.440 73.770 ;
        RECT 130.680 73.600 130.850 73.770 ;
        RECT 131.110 73.600 131.280 73.770 ;
        RECT 131.550 73.600 131.720 73.770 ;
        RECT 131.960 73.600 132.130 73.770 ;
        RECT 134.680 73.650 134.850 73.820 ;
        RECT 135.040 73.650 135.210 73.820 ;
        RECT 137.510 73.600 137.680 73.770 ;
        RECT 137.950 73.600 138.120 73.770 ;
        RECT 138.360 73.600 138.530 73.770 ;
        RECT 138.790 73.600 138.960 73.770 ;
        RECT 139.230 73.600 139.400 73.770 ;
        RECT 139.640 73.600 139.810 73.770 ;
        RECT 5.920 73.170 6.090 73.350 ;
        RECT 6.400 73.170 6.570 73.350 ;
        RECT 6.880 73.170 7.050 73.350 ;
        RECT 7.360 73.170 7.530 73.350 ;
        RECT 7.840 73.170 8.010 73.350 ;
        RECT 8.320 73.170 8.490 73.350 ;
        RECT 8.800 73.170 8.970 73.350 ;
        RECT 9.280 73.170 9.450 73.350 ;
        RECT 9.760 73.170 9.930 73.350 ;
        RECT 10.240 73.170 10.410 73.350 ;
        RECT 10.720 73.170 10.890 73.350 ;
        RECT 11.200 73.170 11.370 73.350 ;
        RECT 11.680 73.170 11.850 73.350 ;
        RECT 12.160 73.170 12.330 73.350 ;
        RECT 12.640 73.170 12.810 73.350 ;
        RECT 13.120 73.170 13.290 73.350 ;
        RECT 13.600 73.170 13.770 73.350 ;
        RECT 14.080 73.170 14.250 73.350 ;
        RECT 14.560 73.170 14.730 73.350 ;
        RECT 15.040 73.170 15.210 73.350 ;
        RECT 15.520 73.170 15.690 73.350 ;
        RECT 16.000 73.170 16.170 73.350 ;
        RECT 16.480 73.170 16.650 73.350 ;
        RECT 16.960 73.170 17.130 73.350 ;
        RECT 17.440 73.170 17.610 73.350 ;
        RECT 17.920 73.170 18.090 73.350 ;
        RECT 18.400 73.170 18.570 73.350 ;
        RECT 18.880 73.170 19.050 73.350 ;
        RECT 19.360 73.170 19.530 73.350 ;
        RECT 19.840 73.170 20.010 73.350 ;
        RECT 20.320 73.170 20.490 73.350 ;
        RECT 20.800 73.170 20.970 73.350 ;
        RECT 21.280 73.170 21.450 73.350 ;
        RECT 21.760 73.170 21.930 73.350 ;
        RECT 22.240 73.170 22.410 73.350 ;
        RECT 22.720 73.170 22.890 73.350 ;
        RECT 23.200 73.170 23.370 73.350 ;
        RECT 23.680 73.170 23.850 73.350 ;
        RECT 24.160 73.170 24.330 73.350 ;
        RECT 24.640 73.170 24.810 73.350 ;
        RECT 25.120 73.170 25.290 73.350 ;
        RECT 25.600 73.170 25.770 73.350 ;
        RECT 26.080 73.170 26.250 73.350 ;
        RECT 26.560 73.170 26.730 73.350 ;
        RECT 27.040 73.170 27.210 73.350 ;
        RECT 27.520 73.170 27.690 73.350 ;
        RECT 28.000 73.170 28.170 73.350 ;
        RECT 28.480 73.170 28.650 73.350 ;
        RECT 28.960 73.170 29.130 73.350 ;
        RECT 29.440 73.170 29.610 73.350 ;
        RECT 29.920 73.170 30.090 73.350 ;
        RECT 30.400 73.170 30.570 73.350 ;
        RECT 30.880 73.170 31.050 73.350 ;
        RECT 31.360 73.170 31.530 73.350 ;
        RECT 31.840 73.170 32.010 73.350 ;
        RECT 32.320 73.170 32.490 73.350 ;
        RECT 32.800 73.170 32.970 73.350 ;
        RECT 33.280 73.170 33.450 73.350 ;
        RECT 33.760 73.170 33.930 73.350 ;
        RECT 34.240 73.170 34.410 73.350 ;
        RECT 34.720 73.170 34.890 73.350 ;
        RECT 35.200 73.170 35.370 73.350 ;
        RECT 35.680 73.170 35.850 73.350 ;
        RECT 36.160 73.170 36.330 73.350 ;
        RECT 36.640 73.170 36.810 73.350 ;
        RECT 37.120 73.170 37.290 73.350 ;
        RECT 37.600 73.170 37.770 73.350 ;
        RECT 38.080 73.170 38.250 73.350 ;
        RECT 38.560 73.170 38.730 73.350 ;
        RECT 39.040 73.170 39.210 73.350 ;
        RECT 39.520 73.170 39.690 73.350 ;
        RECT 40.000 73.170 40.170 73.350 ;
        RECT 40.480 73.170 40.650 73.350 ;
        RECT 40.960 73.170 41.130 73.350 ;
        RECT 41.440 73.170 41.610 73.350 ;
        RECT 41.920 73.170 42.090 73.350 ;
        RECT 42.400 73.170 42.570 73.350 ;
        RECT 42.880 73.170 43.050 73.350 ;
        RECT 43.360 73.170 43.530 73.350 ;
        RECT 43.840 73.170 44.010 73.350 ;
        RECT 44.320 73.170 44.490 73.350 ;
        RECT 44.800 73.170 44.970 73.350 ;
        RECT 45.280 73.170 45.450 73.350 ;
        RECT 45.760 73.170 45.930 73.350 ;
        RECT 46.240 73.170 46.410 73.350 ;
        RECT 46.720 73.170 46.890 73.350 ;
        RECT 47.200 73.340 47.370 73.350 ;
      LAYER li1 ;
        RECT 47.520 73.340 48.000 73.350 ;
        RECT 47.040 73.170 47.520 73.340 ;
      LAYER li1 ;
        RECT 47.680 73.170 47.850 73.340 ;
        RECT 48.160 73.170 48.330 73.350 ;
        RECT 48.640 73.170 48.810 73.350 ;
        RECT 49.120 73.170 49.290 73.350 ;
        RECT 49.600 73.170 49.770 73.350 ;
        RECT 50.080 73.170 50.250 73.350 ;
        RECT 50.560 73.170 50.730 73.350 ;
        RECT 51.040 73.170 51.210 73.350 ;
        RECT 51.520 73.170 51.690 73.350 ;
        RECT 52.000 73.170 52.170 73.350 ;
        RECT 52.480 73.170 52.650 73.350 ;
        RECT 52.960 73.170 53.130 73.350 ;
        RECT 53.440 73.170 53.610 73.350 ;
        RECT 53.920 73.170 54.090 73.350 ;
        RECT 54.400 73.170 54.570 73.350 ;
        RECT 54.880 73.170 55.050 73.350 ;
        RECT 55.360 73.170 55.530 73.350 ;
        RECT 55.840 73.170 56.010 73.350 ;
        RECT 56.320 73.170 56.490 73.350 ;
        RECT 56.800 73.170 56.970 73.350 ;
        RECT 57.280 73.170 57.450 73.350 ;
        RECT 57.760 73.170 57.930 73.350 ;
        RECT 58.240 73.170 58.410 73.350 ;
        RECT 58.720 73.170 58.890 73.350 ;
      LAYER li1 ;
        RECT 59.040 73.340 59.520 73.350 ;
      LAYER li1 ;
        RECT 59.200 73.170 59.370 73.340 ;
        RECT 59.680 73.170 59.850 73.350 ;
        RECT 60.160 73.170 60.330 73.350 ;
        RECT 60.640 73.170 60.810 73.350 ;
        RECT 61.120 73.170 61.290 73.350 ;
        RECT 61.600 73.170 61.770 73.350 ;
        RECT 62.080 73.170 62.250 73.350 ;
        RECT 62.560 73.170 62.730 73.350 ;
        RECT 63.040 73.170 63.210 73.350 ;
        RECT 63.520 73.170 63.690 73.350 ;
        RECT 64.000 73.170 64.170 73.350 ;
        RECT 64.480 73.170 64.650 73.350 ;
        RECT 64.960 73.170 65.130 73.350 ;
        RECT 65.440 73.170 65.610 73.350 ;
        RECT 65.920 73.170 66.090 73.350 ;
        RECT 66.400 73.170 66.570 73.350 ;
        RECT 66.880 73.170 67.050 73.350 ;
        RECT 67.360 73.170 67.530 73.350 ;
        RECT 67.840 73.170 68.010 73.350 ;
        RECT 68.320 73.170 68.490 73.350 ;
        RECT 68.800 73.170 68.970 73.350 ;
        RECT 69.280 73.170 69.450 73.350 ;
        RECT 69.760 73.170 69.930 73.350 ;
        RECT 70.240 73.170 70.410 73.350 ;
        RECT 70.720 73.170 70.890 73.350 ;
        RECT 71.200 73.170 71.370 73.350 ;
        RECT 71.680 73.170 71.850 73.350 ;
        RECT 72.160 73.170 72.330 73.350 ;
        RECT 72.640 73.170 72.810 73.350 ;
        RECT 73.120 73.170 73.290 73.350 ;
        RECT 73.600 73.170 73.770 73.350 ;
        RECT 74.080 73.170 74.250 73.350 ;
        RECT 74.560 73.170 74.730 73.350 ;
        RECT 75.040 73.170 75.210 73.350 ;
        RECT 75.520 73.170 75.690 73.350 ;
        RECT 76.000 73.170 76.170 73.350 ;
      LAYER li1 ;
        RECT 76.320 73.340 76.800 73.350 ;
      LAYER li1 ;
        RECT 76.480 73.170 76.650 73.340 ;
        RECT 76.960 73.170 77.130 73.350 ;
        RECT 77.440 73.170 77.610 73.350 ;
        RECT 77.920 73.170 78.090 73.350 ;
        RECT 78.400 73.170 78.570 73.350 ;
        RECT 78.880 73.340 79.050 73.350 ;
      LAYER li1 ;
        RECT 78.720 73.170 79.200 73.340 ;
      LAYER li1 ;
        RECT 79.360 73.170 79.530 73.350 ;
        RECT 79.840 73.170 80.010 73.350 ;
        RECT 80.320 73.170 80.490 73.350 ;
        RECT 80.800 73.170 80.970 73.350 ;
        RECT 81.280 73.170 81.450 73.350 ;
        RECT 81.760 73.170 81.930 73.350 ;
        RECT 82.240 73.170 82.410 73.350 ;
        RECT 82.720 73.170 82.890 73.350 ;
        RECT 83.200 73.170 83.370 73.350 ;
        RECT 83.680 73.170 83.850 73.350 ;
        RECT 84.160 73.170 84.330 73.350 ;
        RECT 84.640 73.170 84.810 73.350 ;
        RECT 85.120 73.170 85.290 73.350 ;
        RECT 85.600 73.170 85.770 73.350 ;
        RECT 86.080 73.170 86.250 73.350 ;
        RECT 86.560 73.170 86.730 73.350 ;
        RECT 87.040 73.170 87.210 73.350 ;
        RECT 87.520 73.170 87.690 73.350 ;
        RECT 88.000 73.170 88.170 73.350 ;
        RECT 88.480 73.170 88.650 73.350 ;
        RECT 88.960 73.170 89.130 73.350 ;
        RECT 89.440 73.170 89.610 73.350 ;
        RECT 89.920 73.170 90.090 73.350 ;
        RECT 90.400 73.170 90.570 73.350 ;
        RECT 90.880 73.170 91.050 73.350 ;
        RECT 91.360 73.170 91.530 73.350 ;
        RECT 91.840 73.170 92.010 73.350 ;
        RECT 92.320 73.170 92.490 73.350 ;
        RECT 92.800 73.170 92.970 73.350 ;
        RECT 93.280 73.170 93.450 73.350 ;
        RECT 93.760 73.170 93.930 73.350 ;
        RECT 94.240 73.170 94.410 73.350 ;
        RECT 94.720 73.170 94.890 73.350 ;
        RECT 95.200 73.170 95.370 73.350 ;
        RECT 95.680 73.170 95.850 73.350 ;
        RECT 96.160 73.170 96.330 73.350 ;
        RECT 96.640 73.170 96.810 73.350 ;
        RECT 97.120 73.170 97.290 73.350 ;
        RECT 97.600 73.170 97.770 73.350 ;
        RECT 98.080 73.170 98.250 73.350 ;
        RECT 98.560 73.170 98.730 73.350 ;
        RECT 99.040 73.170 99.210 73.350 ;
        RECT 99.520 73.170 99.690 73.350 ;
        RECT 100.000 73.170 100.170 73.350 ;
        RECT 100.480 73.170 100.650 73.350 ;
        RECT 100.960 73.170 101.130 73.350 ;
        RECT 101.440 73.170 101.610 73.350 ;
        RECT 101.920 73.170 102.090 73.350 ;
        RECT 102.400 73.170 102.570 73.350 ;
        RECT 102.880 73.170 103.050 73.350 ;
        RECT 103.360 73.170 103.530 73.350 ;
        RECT 103.840 73.170 104.010 73.350 ;
        RECT 104.320 73.170 104.490 73.350 ;
        RECT 104.800 73.170 104.970 73.350 ;
        RECT 105.280 73.170 105.450 73.350 ;
        RECT 105.760 73.170 105.930 73.350 ;
        RECT 106.240 73.170 106.410 73.350 ;
        RECT 106.720 73.170 106.890 73.350 ;
        RECT 107.200 73.170 107.370 73.350 ;
        RECT 107.680 73.170 107.850 73.350 ;
        RECT 108.160 73.170 108.330 73.350 ;
        RECT 108.640 73.170 108.810 73.350 ;
        RECT 109.120 73.170 109.290 73.350 ;
        RECT 109.600 73.170 109.770 73.350 ;
        RECT 110.080 73.170 110.250 73.350 ;
        RECT 110.560 73.170 110.730 73.350 ;
        RECT 111.040 73.170 111.210 73.350 ;
        RECT 111.520 73.170 111.690 73.350 ;
        RECT 112.000 73.170 112.170 73.350 ;
        RECT 112.480 73.170 112.650 73.350 ;
        RECT 112.960 73.170 113.130 73.350 ;
        RECT 113.440 73.170 113.610 73.350 ;
        RECT 113.920 73.170 114.090 73.350 ;
        RECT 114.400 73.170 114.570 73.350 ;
        RECT 114.880 73.170 115.050 73.350 ;
        RECT 115.360 73.170 115.530 73.350 ;
        RECT 115.840 73.170 116.010 73.350 ;
        RECT 116.320 73.170 116.490 73.350 ;
        RECT 116.800 73.170 116.970 73.350 ;
        RECT 117.280 73.170 117.450 73.350 ;
        RECT 117.760 73.170 117.930 73.350 ;
        RECT 118.240 73.170 118.410 73.350 ;
        RECT 118.720 73.170 118.890 73.350 ;
        RECT 119.200 73.170 119.370 73.350 ;
        RECT 119.680 73.170 119.850 73.350 ;
        RECT 120.160 73.170 120.330 73.350 ;
        RECT 120.640 73.170 120.810 73.350 ;
        RECT 121.120 73.170 121.290 73.350 ;
        RECT 121.600 73.170 121.770 73.350 ;
        RECT 122.080 73.170 122.250 73.350 ;
        RECT 122.560 73.170 122.730 73.350 ;
        RECT 123.040 73.170 123.210 73.350 ;
        RECT 123.520 73.170 123.690 73.350 ;
        RECT 124.000 73.170 124.170 73.350 ;
        RECT 124.480 73.170 124.650 73.350 ;
        RECT 124.960 73.170 125.130 73.350 ;
        RECT 125.440 73.170 125.610 73.350 ;
        RECT 125.920 73.170 126.090 73.350 ;
        RECT 126.400 73.170 126.570 73.350 ;
        RECT 126.880 73.170 127.050 73.350 ;
        RECT 127.360 73.170 127.530 73.350 ;
        RECT 127.840 73.170 128.010 73.350 ;
        RECT 128.320 73.170 128.490 73.350 ;
        RECT 128.800 73.170 128.970 73.350 ;
        RECT 129.280 73.170 129.450 73.350 ;
        RECT 129.760 73.170 129.930 73.350 ;
        RECT 130.240 73.170 130.410 73.350 ;
        RECT 130.720 73.170 130.890 73.350 ;
        RECT 131.200 73.170 131.370 73.350 ;
        RECT 131.680 73.170 131.850 73.350 ;
        RECT 132.160 73.170 132.330 73.350 ;
        RECT 132.640 73.170 132.810 73.350 ;
        RECT 133.120 73.170 133.290 73.350 ;
        RECT 133.600 73.170 133.770 73.350 ;
        RECT 134.080 73.340 134.250 73.350 ;
      LAYER li1 ;
        RECT 133.920 73.170 134.400 73.340 ;
      LAYER li1 ;
        RECT 134.560 73.170 134.730 73.350 ;
        RECT 135.040 73.170 135.210 73.350 ;
        RECT 135.520 73.170 135.690 73.350 ;
        RECT 136.000 73.170 136.170 73.350 ;
        RECT 136.480 73.170 136.650 73.350 ;
        RECT 136.960 73.170 137.130 73.350 ;
        RECT 137.440 73.170 137.610 73.350 ;
        RECT 137.920 73.170 138.090 73.350 ;
        RECT 138.400 73.170 138.570 73.350 ;
        RECT 138.880 73.170 139.050 73.350 ;
        RECT 139.360 73.170 139.530 73.350 ;
        RECT 139.840 73.170 140.010 73.350 ;
        RECT 140.320 73.170 140.490 73.350 ;
        RECT 140.800 73.170 140.970 73.350 ;
        RECT 141.280 73.170 141.450 73.350 ;
        RECT 141.760 73.340 141.930 73.350 ;
      LAYER li1 ;
        RECT 141.600 73.170 142.080 73.340 ;
      LAYER li1 ;
        RECT 6.470 72.750 6.640 72.920 ;
        RECT 6.910 72.750 7.080 72.920 ;
        RECT 7.320 72.750 7.490 72.920 ;
        RECT 7.750 72.750 7.920 72.920 ;
        RECT 8.190 72.750 8.360 72.920 ;
        RECT 8.600 72.750 8.770 72.920 ;
        RECT 10.100 72.750 10.270 72.920 ;
        RECT 10.460 72.750 10.630 72.920 ;
        RECT 10.900 72.750 11.070 72.920 ;
        RECT 13.220 72.700 13.390 72.870 ;
        RECT 13.580 72.700 13.750 72.870 ;
        RECT 15.380 72.750 15.550 72.920 ;
        RECT 15.740 72.750 15.910 72.920 ;
        RECT 16.180 72.750 16.350 72.920 ;
        RECT 17.540 72.700 17.710 72.870 ;
        RECT 17.900 72.700 18.070 72.870 ;
        RECT 19.700 72.750 19.870 72.920 ;
        RECT 20.060 72.750 20.230 72.920 ;
        RECT 20.500 72.750 20.670 72.920 ;
        RECT 21.810 72.700 21.980 72.870 ;
        RECT 22.170 72.700 22.340 72.870 ;
        RECT 22.530 72.700 22.700 72.870 ;
        RECT 22.890 72.700 23.060 72.870 ;
        RECT 24.980 72.750 25.150 72.920 ;
        RECT 25.340 72.750 25.510 72.920 ;
        RECT 25.780 72.750 25.950 72.920 ;
        RECT 26.520 72.700 26.690 72.870 ;
        RECT 26.880 72.700 27.050 72.870 ;
        RECT 27.240 72.700 27.410 72.870 ;
        RECT 28.080 72.700 28.250 72.870 ;
        RECT 28.440 72.700 28.610 72.870 ;
        RECT 28.800 72.700 28.970 72.870 ;
        RECT 29.720 72.700 29.890 72.870 ;
        RECT 30.080 72.700 30.250 72.870 ;
        RECT 30.440 72.700 30.610 72.870 ;
        RECT 31.700 72.750 31.870 72.920 ;
        RECT 32.060 72.750 32.230 72.920 ;
        RECT 32.500 72.750 32.670 72.920 ;
        RECT 33.240 72.700 33.410 72.870 ;
        RECT 33.600 72.700 33.770 72.870 ;
        RECT 33.960 72.700 34.130 72.870 ;
        RECT 34.800 72.700 34.970 72.870 ;
        RECT 35.160 72.700 35.330 72.870 ;
        RECT 35.520 72.700 35.690 72.870 ;
        RECT 36.440 72.700 36.610 72.870 ;
        RECT 36.800 72.700 36.970 72.870 ;
        RECT 37.160 72.700 37.330 72.870 ;
        RECT 38.420 72.750 38.590 72.920 ;
        RECT 38.780 72.750 38.950 72.920 ;
        RECT 39.220 72.750 39.390 72.920 ;
        RECT 39.960 72.700 40.130 72.870 ;
        RECT 40.320 72.700 40.490 72.870 ;
        RECT 40.680 72.700 40.850 72.870 ;
        RECT 41.520 72.700 41.690 72.870 ;
        RECT 41.880 72.700 42.050 72.870 ;
        RECT 42.240 72.700 42.410 72.870 ;
        RECT 43.160 72.700 43.330 72.870 ;
        RECT 43.520 72.700 43.690 72.870 ;
        RECT 43.880 72.700 44.050 72.870 ;
        RECT 45.140 72.750 45.310 72.920 ;
        RECT 45.500 72.750 45.670 72.920 ;
        RECT 45.940 72.750 46.110 72.920 ;
        RECT 48.120 72.700 48.290 72.870 ;
        RECT 48.480 72.700 48.650 72.870 ;
        RECT 48.840 72.700 49.010 72.870 ;
        RECT 49.680 72.700 49.850 72.870 ;
        RECT 50.040 72.700 50.210 72.870 ;
        RECT 50.400 72.700 50.570 72.870 ;
        RECT 51.320 72.700 51.490 72.870 ;
        RECT 51.680 72.700 51.850 72.870 ;
        RECT 52.040 72.700 52.210 72.870 ;
        RECT 53.300 72.750 53.470 72.920 ;
        RECT 53.660 72.750 53.830 72.920 ;
        RECT 54.100 72.750 54.270 72.920 ;
        RECT 54.840 72.700 55.010 72.870 ;
        RECT 55.200 72.700 55.370 72.870 ;
        RECT 55.560 72.700 55.730 72.870 ;
        RECT 55.920 72.700 56.090 72.870 ;
        RECT 56.280 72.700 56.450 72.870 ;
        RECT 57.620 72.750 57.790 72.920 ;
        RECT 57.980 72.750 58.150 72.920 ;
        RECT 58.420 72.750 58.590 72.920 ;
        RECT 59.640 72.700 59.810 72.870 ;
        RECT 60.000 72.700 60.170 72.870 ;
        RECT 60.360 72.700 60.530 72.870 ;
        RECT 61.200 72.700 61.370 72.870 ;
        RECT 61.560 72.700 61.730 72.870 ;
        RECT 61.920 72.700 62.090 72.870 ;
        RECT 62.840 72.700 63.010 72.870 ;
        RECT 63.200 72.700 63.370 72.870 ;
        RECT 63.560 72.700 63.730 72.870 ;
        RECT 64.820 72.750 64.990 72.920 ;
        RECT 65.180 72.750 65.350 72.920 ;
        RECT 65.620 72.750 65.790 72.920 ;
        RECT 66.360 72.700 66.530 72.870 ;
        RECT 66.720 72.700 66.890 72.870 ;
        RECT 67.080 72.700 67.250 72.870 ;
        RECT 67.920 72.700 68.090 72.870 ;
        RECT 68.280 72.700 68.450 72.870 ;
        RECT 68.640 72.700 68.810 72.870 ;
        RECT 69.560 72.700 69.730 72.870 ;
        RECT 69.920 72.700 70.090 72.870 ;
        RECT 70.280 72.700 70.450 72.870 ;
        RECT 71.540 72.750 71.710 72.920 ;
        RECT 71.900 72.750 72.070 72.920 ;
        RECT 72.340 72.750 72.510 72.920 ;
        RECT 73.080 72.700 73.250 72.870 ;
        RECT 73.440 72.700 73.610 72.870 ;
        RECT 74.900 72.750 75.070 72.920 ;
        RECT 75.260 72.750 75.430 72.920 ;
        RECT 75.700 72.750 75.870 72.920 ;
        RECT 77.490 72.700 77.660 72.870 ;
        RECT 77.850 72.700 78.020 72.870 ;
        RECT 78.210 72.700 78.380 72.870 ;
        RECT 78.570 72.700 78.740 72.870 ;
        RECT 80.660 72.750 80.830 72.920 ;
        RECT 81.020 72.750 81.190 72.920 ;
        RECT 81.460 72.750 81.630 72.920 ;
        RECT 82.200 72.700 82.370 72.870 ;
        RECT 82.560 72.700 82.730 72.870 ;
        RECT 82.920 72.700 83.090 72.870 ;
        RECT 83.760 72.700 83.930 72.870 ;
        RECT 84.120 72.700 84.290 72.870 ;
        RECT 84.480 72.700 84.650 72.870 ;
        RECT 85.400 72.700 85.570 72.870 ;
        RECT 85.760 72.700 85.930 72.870 ;
        RECT 86.120 72.700 86.290 72.870 ;
        RECT 87.380 72.750 87.550 72.920 ;
        RECT 87.740 72.750 87.910 72.920 ;
        RECT 88.180 72.750 88.350 72.920 ;
        RECT 88.920 72.700 89.090 72.870 ;
        RECT 89.280 72.700 89.450 72.870 ;
        RECT 89.640 72.700 89.810 72.870 ;
        RECT 90.480 72.700 90.650 72.870 ;
        RECT 90.840 72.700 91.010 72.870 ;
        RECT 91.200 72.700 91.370 72.870 ;
        RECT 92.120 72.700 92.290 72.870 ;
        RECT 92.480 72.700 92.650 72.870 ;
        RECT 92.840 72.700 93.010 72.870 ;
        RECT 94.100 72.750 94.270 72.920 ;
        RECT 94.460 72.750 94.630 72.920 ;
        RECT 94.900 72.750 95.070 72.920 ;
        RECT 95.640 72.700 95.810 72.870 ;
        RECT 96.000 72.700 96.170 72.870 ;
        RECT 97.460 72.750 97.630 72.920 ;
        RECT 97.820 72.750 97.990 72.920 ;
        RECT 98.260 72.750 98.430 72.920 ;
        RECT 99.570 72.700 99.740 72.870 ;
        RECT 99.930 72.700 100.100 72.870 ;
        RECT 100.290 72.700 100.460 72.870 ;
        RECT 100.650 72.700 100.820 72.870 ;
        RECT 102.740 72.750 102.910 72.920 ;
        RECT 103.100 72.750 103.270 72.920 ;
        RECT 103.540 72.750 103.710 72.920 ;
        RECT 104.280 72.700 104.450 72.870 ;
        RECT 104.640 72.700 104.810 72.870 ;
        RECT 105.000 72.700 105.170 72.870 ;
        RECT 105.850 72.700 106.020 72.870 ;
        RECT 106.210 72.700 106.380 72.870 ;
        RECT 107.060 72.750 107.230 72.920 ;
        RECT 107.420 72.750 107.590 72.920 ;
        RECT 107.860 72.750 108.030 72.920 ;
        RECT 108.600 72.700 108.770 72.870 ;
        RECT 108.960 72.700 109.130 72.870 ;
        RECT 109.320 72.700 109.490 72.870 ;
        RECT 109.680 72.700 109.850 72.870 ;
        RECT 110.040 72.700 110.210 72.870 ;
        RECT 111.380 72.750 111.550 72.920 ;
        RECT 111.740 72.750 111.910 72.920 ;
        RECT 112.180 72.750 112.350 72.920 ;
        RECT 112.920 72.700 113.090 72.870 ;
        RECT 113.280 72.700 113.450 72.870 ;
        RECT 114.740 72.750 114.910 72.920 ;
        RECT 115.100 72.750 115.270 72.920 ;
        RECT 115.540 72.750 115.710 72.920 ;
        RECT 116.280 72.700 116.450 72.870 ;
        RECT 116.640 72.700 116.810 72.870 ;
        RECT 117.000 72.700 117.170 72.870 ;
        RECT 117.840 72.700 118.010 72.870 ;
        RECT 118.200 72.700 118.370 72.870 ;
        RECT 118.560 72.700 118.730 72.870 ;
        RECT 119.480 72.700 119.650 72.870 ;
        RECT 119.840 72.700 120.010 72.870 ;
        RECT 120.200 72.700 120.370 72.870 ;
        RECT 121.460 72.750 121.630 72.920 ;
        RECT 121.820 72.750 121.990 72.920 ;
        RECT 122.260 72.750 122.430 72.920 ;
        RECT 123.620 72.700 123.790 72.870 ;
        RECT 123.980 72.700 124.150 72.870 ;
        RECT 125.990 72.750 126.160 72.920 ;
        RECT 126.430 72.750 126.600 72.920 ;
        RECT 126.840 72.750 127.010 72.920 ;
        RECT 127.270 72.750 127.440 72.920 ;
        RECT 127.710 72.750 127.880 72.920 ;
        RECT 128.120 72.750 128.290 72.920 ;
        RECT 129.860 72.700 130.030 72.870 ;
        RECT 130.220 72.700 130.390 72.870 ;
        RECT 132.230 72.750 132.400 72.920 ;
        RECT 132.670 72.750 132.840 72.920 ;
        RECT 133.080 72.750 133.250 72.920 ;
        RECT 133.510 72.750 133.680 72.920 ;
        RECT 133.950 72.750 134.120 72.920 ;
        RECT 134.360 72.750 134.530 72.920 ;
        RECT 136.070 72.750 136.240 72.920 ;
        RECT 136.510 72.750 136.680 72.920 ;
        RECT 136.920 72.750 137.090 72.920 ;
        RECT 137.350 72.750 137.520 72.920 ;
        RECT 137.790 72.750 137.960 72.920 ;
        RECT 138.200 72.750 138.370 72.920 ;
        RECT 139.700 72.750 139.870 72.920 ;
        RECT 140.060 72.750 140.230 72.920 ;
        RECT 140.500 72.750 140.670 72.920 ;
        RECT 6.260 65.460 6.430 65.630 ;
        RECT 6.620 65.460 6.790 65.630 ;
        RECT 7.060 65.460 7.230 65.630 ;
        RECT 9.860 65.510 10.030 65.680 ;
        RECT 10.220 65.510 10.390 65.680 ;
        RECT 12.020 65.460 12.190 65.630 ;
        RECT 12.380 65.460 12.550 65.630 ;
        RECT 12.820 65.460 12.990 65.630 ;
        RECT 13.560 65.510 13.730 65.680 ;
        RECT 13.920 65.510 14.090 65.680 ;
        RECT 14.280 65.510 14.450 65.680 ;
        RECT 14.640 65.510 14.810 65.680 ;
        RECT 15.000 65.510 15.170 65.680 ;
        RECT 16.340 65.460 16.510 65.630 ;
        RECT 16.700 65.460 16.870 65.630 ;
        RECT 17.140 65.460 17.310 65.630 ;
        RECT 17.880 65.510 18.050 65.680 ;
        RECT 18.240 65.510 18.410 65.680 ;
        RECT 18.600 65.510 18.770 65.680 ;
        RECT 19.450 65.510 19.620 65.680 ;
        RECT 19.810 65.510 19.980 65.680 ;
        RECT 20.660 65.460 20.830 65.630 ;
        RECT 21.020 65.460 21.190 65.630 ;
        RECT 21.460 65.460 21.630 65.630 ;
        RECT 22.200 65.510 22.370 65.680 ;
        RECT 22.560 65.510 22.730 65.680 ;
        RECT 22.920 65.510 23.090 65.680 ;
        RECT 23.760 65.510 23.930 65.680 ;
        RECT 24.120 65.510 24.290 65.680 ;
        RECT 24.480 65.510 24.650 65.680 ;
        RECT 25.400 65.510 25.570 65.680 ;
        RECT 25.760 65.510 25.930 65.680 ;
        RECT 26.120 65.510 26.290 65.680 ;
        RECT 27.380 65.460 27.550 65.630 ;
        RECT 27.740 65.460 27.910 65.630 ;
        RECT 28.180 65.460 28.350 65.630 ;
        RECT 28.920 65.510 29.090 65.680 ;
        RECT 29.280 65.510 29.450 65.680 ;
        RECT 29.640 65.510 29.810 65.680 ;
        RECT 30.480 65.510 30.650 65.680 ;
        RECT 30.840 65.510 31.010 65.680 ;
        RECT 31.200 65.510 31.370 65.680 ;
        RECT 32.120 65.510 32.290 65.680 ;
        RECT 32.480 65.510 32.650 65.680 ;
        RECT 32.840 65.510 33.010 65.680 ;
        RECT 34.100 65.460 34.270 65.630 ;
        RECT 34.460 65.460 34.630 65.630 ;
        RECT 34.900 65.460 35.070 65.630 ;
        RECT 35.640 65.510 35.810 65.680 ;
        RECT 36.000 65.510 36.170 65.680 ;
        RECT 37.460 65.460 37.630 65.630 ;
        RECT 37.820 65.460 37.990 65.630 ;
        RECT 38.260 65.460 38.430 65.630 ;
        RECT 39.000 65.510 39.170 65.680 ;
        RECT 39.360 65.510 39.530 65.680 ;
        RECT 39.720 65.510 39.890 65.680 ;
        RECT 40.560 65.510 40.730 65.680 ;
        RECT 40.920 65.510 41.090 65.680 ;
        RECT 41.280 65.510 41.450 65.680 ;
        RECT 42.200 65.510 42.370 65.680 ;
        RECT 42.560 65.510 42.730 65.680 ;
        RECT 42.920 65.510 43.090 65.680 ;
        RECT 44.390 65.460 44.560 65.630 ;
        RECT 44.830 65.460 45.000 65.630 ;
        RECT 45.240 65.460 45.410 65.630 ;
        RECT 45.670 65.460 45.840 65.630 ;
        RECT 46.110 65.460 46.280 65.630 ;
        RECT 46.520 65.460 46.690 65.630 ;
        RECT 48.120 65.510 48.290 65.680 ;
        RECT 48.480 65.510 48.650 65.680 ;
        RECT 48.840 65.510 49.010 65.680 ;
        RECT 49.680 65.510 49.850 65.680 ;
        RECT 50.040 65.510 50.210 65.680 ;
        RECT 50.400 65.510 50.570 65.680 ;
        RECT 51.320 65.510 51.490 65.680 ;
        RECT 51.680 65.510 51.850 65.680 ;
        RECT 52.040 65.510 52.210 65.680 ;
        RECT 53.510 65.460 53.680 65.630 ;
        RECT 53.950 65.460 54.120 65.630 ;
        RECT 54.360 65.460 54.530 65.630 ;
        RECT 54.790 65.460 54.960 65.630 ;
        RECT 55.230 65.460 55.400 65.630 ;
        RECT 55.640 65.460 55.810 65.630 ;
        RECT 57.720 65.510 57.890 65.680 ;
        RECT 58.080 65.510 58.250 65.680 ;
        RECT 58.440 65.510 58.610 65.680 ;
        RECT 59.280 65.510 59.450 65.680 ;
        RECT 59.640 65.510 59.810 65.680 ;
        RECT 60.000 65.510 60.170 65.680 ;
        RECT 60.920 65.510 61.090 65.680 ;
        RECT 61.280 65.510 61.450 65.680 ;
        RECT 61.640 65.510 61.810 65.680 ;
        RECT 62.900 65.460 63.070 65.630 ;
        RECT 63.260 65.460 63.430 65.630 ;
        RECT 63.700 65.460 63.870 65.630 ;
        RECT 64.440 65.510 64.610 65.680 ;
        RECT 64.800 65.510 64.970 65.680 ;
        RECT 65.160 65.510 65.330 65.680 ;
        RECT 66.000 65.510 66.170 65.680 ;
        RECT 66.360 65.510 66.530 65.680 ;
        RECT 66.720 65.510 66.890 65.680 ;
        RECT 67.640 65.510 67.810 65.680 ;
        RECT 68.000 65.510 68.170 65.680 ;
        RECT 68.360 65.510 68.530 65.680 ;
        RECT 69.620 65.460 69.790 65.630 ;
        RECT 69.980 65.460 70.150 65.630 ;
        RECT 70.420 65.460 70.590 65.630 ;
        RECT 71.160 65.510 71.330 65.680 ;
        RECT 71.520 65.510 71.690 65.680 ;
        RECT 71.880 65.510 72.050 65.680 ;
        RECT 72.720 65.510 72.890 65.680 ;
        RECT 73.080 65.510 73.250 65.680 ;
        RECT 73.440 65.510 73.610 65.680 ;
        RECT 74.360 65.510 74.530 65.680 ;
        RECT 74.720 65.510 74.890 65.680 ;
        RECT 75.080 65.510 75.250 65.680 ;
        RECT 76.340 65.460 76.510 65.630 ;
        RECT 76.700 65.460 76.870 65.630 ;
        RECT 77.140 65.460 77.310 65.630 ;
        RECT 77.870 65.510 78.040 65.680 ;
        RECT 78.230 65.510 78.400 65.680 ;
        RECT 78.590 65.510 78.760 65.680 ;
        RECT 79.310 65.510 79.480 65.680 ;
        RECT 79.670 65.510 79.840 65.680 ;
        RECT 80.030 65.510 80.200 65.680 ;
        RECT 80.390 65.510 80.560 65.680 ;
        RECT 81.620 65.460 81.790 65.630 ;
        RECT 81.980 65.460 82.150 65.630 ;
        RECT 82.420 65.460 82.590 65.630 ;
        RECT 83.590 65.510 83.760 65.680 ;
        RECT 83.950 65.510 84.120 65.680 ;
        RECT 84.310 65.510 84.480 65.680 ;
        RECT 85.900 65.510 86.070 65.680 ;
        RECT 86.260 65.510 86.430 65.680 ;
        RECT 86.620 65.510 86.790 65.680 ;
        RECT 88.070 65.460 88.240 65.630 ;
        RECT 88.510 65.460 88.680 65.630 ;
        RECT 88.920 65.460 89.090 65.630 ;
        RECT 89.350 65.460 89.520 65.630 ;
        RECT 89.790 65.460 89.960 65.630 ;
        RECT 90.200 65.460 90.370 65.630 ;
        RECT 92.340 65.510 92.510 65.680 ;
        RECT 92.700 65.510 92.870 65.680 ;
        RECT 94.730 65.510 94.900 65.680 ;
        RECT 97.160 65.510 97.330 65.680 ;
        RECT 97.520 65.510 97.690 65.680 ;
        RECT 97.880 65.510 98.050 65.680 ;
        RECT 99.500 65.510 99.670 65.680 ;
        RECT 99.860 65.510 100.030 65.680 ;
        RECT 100.220 65.510 100.390 65.680 ;
        RECT 102.200 65.510 102.370 65.680 ;
        RECT 102.560 65.510 102.730 65.680 ;
        RECT 102.920 65.510 103.090 65.680 ;
        RECT 103.950 65.510 104.120 65.680 ;
        RECT 104.310 65.510 104.480 65.680 ;
        RECT 104.670 65.510 104.840 65.680 ;
        RECT 105.480 65.510 105.650 65.680 ;
        RECT 105.840 65.510 106.010 65.680 ;
        RECT 106.200 65.510 106.370 65.680 ;
        RECT 107.750 65.460 107.920 65.630 ;
        RECT 108.190 65.460 108.360 65.630 ;
        RECT 108.600 65.460 108.770 65.630 ;
        RECT 109.030 65.460 109.200 65.630 ;
        RECT 109.470 65.460 109.640 65.630 ;
        RECT 109.880 65.460 110.050 65.630 ;
        RECT 111.000 65.510 111.170 65.680 ;
        RECT 111.360 65.510 111.530 65.680 ;
        RECT 111.720 65.510 111.890 65.680 ;
        RECT 113.130 65.510 113.300 65.680 ;
        RECT 113.490 65.510 113.660 65.680 ;
        RECT 113.850 65.510 114.020 65.680 ;
        RECT 114.740 65.460 114.910 65.630 ;
        RECT 115.100 65.460 115.270 65.630 ;
        RECT 115.540 65.460 115.710 65.630 ;
        RECT 116.280 65.510 116.450 65.680 ;
        RECT 116.640 65.510 116.810 65.680 ;
        RECT 117.000 65.510 117.170 65.680 ;
        RECT 117.840 65.510 118.010 65.680 ;
        RECT 118.200 65.510 118.370 65.680 ;
        RECT 118.560 65.510 118.730 65.680 ;
        RECT 119.480 65.510 119.650 65.680 ;
        RECT 119.840 65.510 120.010 65.680 ;
        RECT 120.200 65.510 120.370 65.680 ;
        RECT 121.460 65.460 121.630 65.630 ;
        RECT 121.820 65.460 121.990 65.630 ;
        RECT 122.260 65.460 122.430 65.630 ;
        RECT 123.000 65.510 123.170 65.680 ;
        RECT 123.360 65.510 123.530 65.680 ;
        RECT 123.720 65.510 123.890 65.680 ;
        RECT 124.080 65.510 124.250 65.680 ;
        RECT 124.440 65.510 124.610 65.680 ;
        RECT 126.950 65.460 127.120 65.630 ;
        RECT 127.390 65.460 127.560 65.630 ;
        RECT 127.800 65.460 127.970 65.630 ;
        RECT 128.230 65.460 128.400 65.630 ;
        RECT 128.670 65.460 128.840 65.630 ;
        RECT 129.080 65.460 129.250 65.630 ;
        RECT 131.300 65.510 131.470 65.680 ;
        RECT 131.660 65.510 131.830 65.680 ;
        RECT 133.460 65.460 133.630 65.630 ;
        RECT 133.820 65.460 133.990 65.630 ;
        RECT 134.260 65.460 134.430 65.630 ;
        RECT 135.000 65.510 135.170 65.680 ;
        RECT 135.360 65.510 135.530 65.680 ;
        RECT 137.030 65.460 137.200 65.630 ;
        RECT 137.470 65.460 137.640 65.630 ;
        RECT 137.880 65.460 138.050 65.630 ;
        RECT 138.310 65.460 138.480 65.630 ;
        RECT 138.750 65.460 138.920 65.630 ;
        RECT 139.160 65.460 139.330 65.630 ;
        RECT 140.660 65.460 140.830 65.630 ;
        RECT 141.020 65.460 141.190 65.630 ;
        RECT 141.460 65.460 141.630 65.630 ;
        RECT 5.920 65.030 6.090 65.210 ;
        RECT 6.400 65.030 6.570 65.210 ;
        RECT 6.880 65.030 7.050 65.210 ;
        RECT 7.360 65.030 7.530 65.210 ;
        RECT 7.840 65.030 8.010 65.210 ;
        RECT 8.320 65.030 8.490 65.210 ;
        RECT 8.800 65.200 8.970 65.210 ;
      LAYER li1 ;
        RECT 8.640 65.030 9.120 65.200 ;
      LAYER li1 ;
        RECT 9.280 65.030 9.450 65.210 ;
        RECT 9.760 65.030 9.930 65.210 ;
        RECT 10.240 65.030 10.410 65.210 ;
        RECT 10.720 65.030 10.890 65.210 ;
        RECT 11.200 65.030 11.370 65.210 ;
        RECT 11.680 65.030 11.850 65.210 ;
        RECT 12.160 65.030 12.330 65.210 ;
        RECT 12.640 65.030 12.810 65.210 ;
        RECT 13.120 65.030 13.290 65.210 ;
        RECT 13.600 65.030 13.770 65.210 ;
        RECT 14.080 65.030 14.250 65.210 ;
        RECT 14.560 65.030 14.730 65.210 ;
        RECT 15.040 65.030 15.210 65.210 ;
        RECT 15.520 65.030 15.690 65.210 ;
        RECT 16.000 65.030 16.170 65.210 ;
        RECT 16.480 65.030 16.650 65.210 ;
        RECT 16.960 65.030 17.130 65.210 ;
        RECT 17.440 65.030 17.610 65.210 ;
        RECT 17.920 65.030 18.090 65.210 ;
        RECT 18.400 65.030 18.570 65.210 ;
        RECT 18.880 65.030 19.050 65.210 ;
        RECT 19.360 65.030 19.530 65.210 ;
        RECT 19.840 65.030 20.010 65.210 ;
        RECT 20.320 65.030 20.490 65.210 ;
        RECT 20.800 65.030 20.970 65.210 ;
        RECT 21.280 65.030 21.450 65.210 ;
        RECT 21.760 65.030 21.930 65.210 ;
        RECT 22.240 65.030 22.410 65.210 ;
        RECT 22.720 65.030 22.890 65.210 ;
        RECT 23.200 65.030 23.370 65.210 ;
        RECT 23.680 65.030 23.850 65.210 ;
        RECT 24.160 65.030 24.330 65.210 ;
        RECT 24.640 65.030 24.810 65.210 ;
        RECT 25.120 65.030 25.290 65.210 ;
        RECT 25.600 65.030 25.770 65.210 ;
        RECT 26.080 65.030 26.250 65.210 ;
        RECT 26.560 65.030 26.730 65.210 ;
        RECT 27.040 65.030 27.210 65.210 ;
        RECT 27.520 65.030 27.690 65.210 ;
        RECT 28.000 65.030 28.170 65.210 ;
        RECT 28.480 65.030 28.650 65.210 ;
        RECT 28.960 65.030 29.130 65.210 ;
        RECT 29.440 65.030 29.610 65.210 ;
        RECT 29.920 65.030 30.090 65.210 ;
        RECT 30.400 65.030 30.570 65.210 ;
        RECT 30.880 65.030 31.050 65.210 ;
        RECT 31.360 65.030 31.530 65.210 ;
        RECT 31.840 65.030 32.010 65.210 ;
        RECT 32.320 65.030 32.490 65.210 ;
        RECT 32.800 65.030 32.970 65.210 ;
        RECT 33.280 65.030 33.450 65.210 ;
        RECT 33.760 65.030 33.930 65.210 ;
        RECT 34.240 65.030 34.410 65.210 ;
        RECT 34.720 65.030 34.890 65.210 ;
        RECT 35.200 65.030 35.370 65.210 ;
        RECT 35.680 65.030 35.850 65.210 ;
        RECT 36.160 65.030 36.330 65.210 ;
        RECT 36.640 65.030 36.810 65.210 ;
        RECT 37.120 65.030 37.290 65.210 ;
        RECT 37.600 65.030 37.770 65.210 ;
        RECT 38.080 65.030 38.250 65.210 ;
        RECT 38.560 65.030 38.730 65.210 ;
        RECT 39.040 65.030 39.210 65.210 ;
        RECT 39.520 65.030 39.690 65.210 ;
        RECT 40.000 65.030 40.170 65.210 ;
        RECT 40.480 65.030 40.650 65.210 ;
        RECT 40.960 65.030 41.130 65.210 ;
        RECT 41.440 65.030 41.610 65.210 ;
        RECT 41.920 65.030 42.090 65.210 ;
        RECT 42.400 65.030 42.570 65.210 ;
        RECT 42.880 65.030 43.050 65.210 ;
        RECT 43.360 65.030 43.530 65.210 ;
        RECT 43.840 65.030 44.010 65.210 ;
        RECT 44.320 65.030 44.490 65.210 ;
        RECT 44.800 65.030 44.970 65.210 ;
        RECT 45.280 65.030 45.450 65.210 ;
        RECT 45.760 65.030 45.930 65.210 ;
        RECT 46.240 65.030 46.410 65.210 ;
        RECT 46.720 65.030 46.890 65.210 ;
        RECT 47.200 65.030 47.370 65.210 ;
        RECT 47.680 65.200 47.850 65.210 ;
      LAYER li1 ;
        RECT 47.520 65.030 48.000 65.200 ;
      LAYER li1 ;
        RECT 48.160 65.030 48.330 65.210 ;
        RECT 48.640 65.030 48.810 65.210 ;
        RECT 49.120 65.030 49.290 65.210 ;
        RECT 49.600 65.030 49.770 65.210 ;
        RECT 50.080 65.030 50.250 65.210 ;
        RECT 50.560 65.030 50.730 65.210 ;
        RECT 51.040 65.030 51.210 65.210 ;
        RECT 51.520 65.030 51.690 65.210 ;
        RECT 52.000 65.030 52.170 65.210 ;
        RECT 52.480 65.030 52.650 65.210 ;
        RECT 52.960 65.030 53.130 65.210 ;
        RECT 53.440 65.030 53.610 65.210 ;
        RECT 53.920 65.030 54.090 65.210 ;
        RECT 54.400 65.030 54.570 65.210 ;
        RECT 54.880 65.030 55.050 65.210 ;
        RECT 55.360 65.030 55.530 65.210 ;
        RECT 55.840 65.030 56.010 65.210 ;
        RECT 56.320 65.030 56.490 65.210 ;
        RECT 56.800 65.030 56.970 65.210 ;
        RECT 57.280 65.030 57.450 65.210 ;
        RECT 57.760 65.030 57.930 65.210 ;
        RECT 58.240 65.030 58.410 65.210 ;
        RECT 58.720 65.030 58.890 65.210 ;
        RECT 59.200 65.030 59.370 65.210 ;
        RECT 59.680 65.030 59.850 65.210 ;
        RECT 60.160 65.030 60.330 65.210 ;
        RECT 60.640 65.030 60.810 65.210 ;
        RECT 61.120 65.030 61.290 65.210 ;
        RECT 61.600 65.030 61.770 65.210 ;
        RECT 62.080 65.030 62.250 65.210 ;
        RECT 62.560 65.030 62.730 65.210 ;
        RECT 63.040 65.030 63.210 65.210 ;
        RECT 63.520 65.030 63.690 65.210 ;
        RECT 64.000 65.030 64.170 65.210 ;
        RECT 64.480 65.030 64.650 65.210 ;
        RECT 64.960 65.030 65.130 65.210 ;
        RECT 65.440 65.030 65.610 65.210 ;
        RECT 65.920 65.030 66.090 65.210 ;
        RECT 66.400 65.030 66.570 65.210 ;
        RECT 66.880 65.030 67.050 65.210 ;
        RECT 67.360 65.030 67.530 65.210 ;
        RECT 67.840 65.030 68.010 65.210 ;
        RECT 68.320 65.030 68.490 65.210 ;
        RECT 68.800 65.030 68.970 65.210 ;
        RECT 69.280 65.030 69.450 65.210 ;
        RECT 69.760 65.030 69.930 65.210 ;
        RECT 70.240 65.030 70.410 65.210 ;
        RECT 70.720 65.030 70.890 65.210 ;
        RECT 71.200 65.030 71.370 65.210 ;
        RECT 71.680 65.030 71.850 65.210 ;
        RECT 72.160 65.030 72.330 65.210 ;
        RECT 72.640 65.030 72.810 65.210 ;
        RECT 73.120 65.030 73.290 65.210 ;
        RECT 73.600 65.030 73.770 65.210 ;
        RECT 74.080 65.030 74.250 65.210 ;
        RECT 74.560 65.030 74.730 65.210 ;
        RECT 75.040 65.030 75.210 65.210 ;
        RECT 75.520 65.030 75.690 65.210 ;
        RECT 76.000 65.030 76.170 65.210 ;
        RECT 76.480 65.030 76.650 65.210 ;
        RECT 76.960 65.030 77.130 65.210 ;
        RECT 77.440 65.030 77.610 65.210 ;
        RECT 77.920 65.030 78.090 65.210 ;
        RECT 78.400 65.030 78.570 65.210 ;
        RECT 78.880 65.030 79.050 65.210 ;
        RECT 79.360 65.030 79.530 65.210 ;
        RECT 79.840 65.030 80.010 65.210 ;
        RECT 80.320 65.030 80.490 65.210 ;
        RECT 80.800 65.030 80.970 65.210 ;
        RECT 81.280 65.030 81.450 65.210 ;
        RECT 81.760 65.030 81.930 65.210 ;
        RECT 82.240 65.030 82.410 65.210 ;
        RECT 82.720 65.030 82.890 65.210 ;
        RECT 83.200 65.030 83.370 65.210 ;
        RECT 83.680 65.030 83.850 65.210 ;
        RECT 84.160 65.030 84.330 65.210 ;
        RECT 84.640 65.030 84.810 65.210 ;
        RECT 85.120 65.030 85.290 65.210 ;
        RECT 85.600 65.030 85.770 65.210 ;
        RECT 86.080 65.030 86.250 65.210 ;
        RECT 86.560 65.030 86.730 65.210 ;
        RECT 87.040 65.030 87.210 65.210 ;
        RECT 87.520 65.030 87.690 65.210 ;
        RECT 88.000 65.030 88.170 65.210 ;
        RECT 88.480 65.030 88.650 65.210 ;
        RECT 88.960 65.030 89.130 65.210 ;
        RECT 89.440 65.030 89.610 65.210 ;
        RECT 89.920 65.030 90.090 65.210 ;
        RECT 90.400 65.030 90.570 65.210 ;
        RECT 90.880 65.030 91.050 65.210 ;
      LAYER li1 ;
        RECT 91.200 65.030 91.680 65.210 ;
      LAYER li1 ;
        RECT 91.840 65.030 92.010 65.210 ;
        RECT 92.320 65.030 92.490 65.210 ;
        RECT 92.800 65.030 92.970 65.210 ;
        RECT 93.280 65.030 93.450 65.210 ;
        RECT 93.760 65.030 93.930 65.210 ;
        RECT 94.240 65.030 94.410 65.210 ;
        RECT 94.720 65.030 94.890 65.210 ;
        RECT 95.200 65.030 95.370 65.210 ;
        RECT 95.680 65.030 95.850 65.210 ;
        RECT 96.160 65.030 96.330 65.210 ;
        RECT 96.640 65.030 96.810 65.210 ;
        RECT 97.120 65.030 97.290 65.210 ;
        RECT 97.600 65.030 97.770 65.210 ;
        RECT 98.080 65.030 98.250 65.210 ;
        RECT 98.560 65.030 98.730 65.210 ;
        RECT 99.040 65.030 99.210 65.210 ;
        RECT 99.520 65.030 99.690 65.210 ;
        RECT 100.000 65.030 100.170 65.210 ;
        RECT 100.480 65.030 100.650 65.210 ;
        RECT 100.960 65.030 101.130 65.210 ;
        RECT 101.440 65.030 101.610 65.210 ;
        RECT 101.920 65.030 102.090 65.210 ;
        RECT 102.400 65.030 102.570 65.210 ;
        RECT 102.880 65.030 103.050 65.210 ;
        RECT 103.360 65.030 103.530 65.210 ;
        RECT 103.840 65.030 104.010 65.210 ;
        RECT 104.320 65.030 104.490 65.210 ;
        RECT 104.800 65.030 104.970 65.210 ;
        RECT 105.280 65.030 105.450 65.210 ;
      LAYER li1 ;
        RECT 105.600 65.200 106.080 65.210 ;
      LAYER li1 ;
        RECT 105.760 65.030 105.930 65.200 ;
        RECT 106.240 65.030 106.410 65.210 ;
        RECT 106.720 65.030 106.890 65.210 ;
        RECT 107.200 65.030 107.370 65.210 ;
        RECT 107.680 65.030 107.850 65.210 ;
        RECT 108.160 65.030 108.330 65.210 ;
        RECT 108.640 65.030 108.810 65.210 ;
        RECT 109.120 65.030 109.290 65.210 ;
        RECT 109.600 65.030 109.770 65.210 ;
        RECT 110.080 65.030 110.250 65.210 ;
        RECT 110.560 65.030 110.730 65.210 ;
        RECT 111.040 65.030 111.210 65.210 ;
        RECT 111.520 65.030 111.690 65.210 ;
        RECT 112.000 65.030 112.170 65.210 ;
        RECT 112.480 65.030 112.650 65.210 ;
        RECT 112.960 65.030 113.130 65.210 ;
        RECT 113.440 65.030 113.610 65.210 ;
        RECT 113.920 65.030 114.090 65.210 ;
        RECT 114.400 65.030 114.570 65.210 ;
        RECT 114.880 65.030 115.050 65.210 ;
        RECT 115.360 65.030 115.530 65.210 ;
        RECT 115.840 65.030 116.010 65.210 ;
        RECT 116.320 65.030 116.490 65.210 ;
        RECT 116.800 65.030 116.970 65.210 ;
        RECT 117.280 65.030 117.450 65.210 ;
        RECT 117.760 65.030 117.930 65.210 ;
        RECT 118.240 65.030 118.410 65.210 ;
        RECT 118.720 65.030 118.890 65.210 ;
        RECT 119.200 65.030 119.370 65.210 ;
        RECT 119.680 65.030 119.850 65.210 ;
        RECT 120.160 65.030 120.330 65.210 ;
        RECT 120.640 65.030 120.810 65.210 ;
        RECT 121.120 65.030 121.290 65.210 ;
        RECT 121.600 65.030 121.770 65.210 ;
        RECT 122.080 65.030 122.250 65.210 ;
        RECT 122.560 65.030 122.730 65.210 ;
        RECT 123.040 65.030 123.210 65.210 ;
        RECT 123.520 65.030 123.690 65.210 ;
        RECT 124.000 65.030 124.170 65.210 ;
        RECT 124.480 65.030 124.650 65.210 ;
        RECT 124.960 65.030 125.130 65.210 ;
        RECT 125.440 65.030 125.610 65.210 ;
        RECT 125.920 65.030 126.090 65.210 ;
        RECT 126.400 65.030 126.570 65.210 ;
        RECT 126.880 65.030 127.050 65.210 ;
        RECT 127.360 65.030 127.530 65.210 ;
        RECT 127.840 65.030 128.010 65.210 ;
        RECT 128.320 65.030 128.490 65.210 ;
        RECT 128.800 65.030 128.970 65.210 ;
        RECT 129.280 65.030 129.450 65.210 ;
        RECT 129.760 65.030 129.930 65.210 ;
        RECT 130.240 65.200 130.410 65.210 ;
      LAYER li1 ;
        RECT 130.080 65.030 130.560 65.200 ;
      LAYER li1 ;
        RECT 130.720 65.030 130.890 65.210 ;
        RECT 131.200 65.030 131.370 65.210 ;
        RECT 131.680 65.030 131.850 65.210 ;
        RECT 132.160 65.030 132.330 65.210 ;
        RECT 132.640 65.030 132.810 65.210 ;
        RECT 133.120 65.030 133.290 65.210 ;
        RECT 133.600 65.030 133.770 65.210 ;
        RECT 134.080 65.030 134.250 65.210 ;
        RECT 134.560 65.030 134.730 65.210 ;
        RECT 135.040 65.030 135.210 65.210 ;
        RECT 135.520 65.030 135.690 65.210 ;
        RECT 136.000 65.030 136.170 65.210 ;
        RECT 136.480 65.030 136.650 65.210 ;
        RECT 136.960 65.030 137.130 65.210 ;
        RECT 137.440 65.030 137.610 65.210 ;
        RECT 137.920 65.030 138.090 65.210 ;
        RECT 138.400 65.030 138.570 65.210 ;
        RECT 138.880 65.030 139.050 65.210 ;
        RECT 139.360 65.030 139.530 65.210 ;
        RECT 139.840 65.030 140.010 65.210 ;
        RECT 140.320 65.030 140.490 65.210 ;
        RECT 140.800 65.030 140.970 65.210 ;
        RECT 141.280 65.030 141.450 65.210 ;
      LAYER li1 ;
        RECT 141.600 65.200 142.080 65.210 ;
      LAYER li1 ;
        RECT 141.760 65.030 141.930 65.200 ;
        RECT 6.260 64.610 6.430 64.780 ;
        RECT 6.620 64.610 6.790 64.780 ;
        RECT 7.060 64.610 7.230 64.780 ;
        RECT 7.800 64.560 7.970 64.730 ;
        RECT 8.160 64.560 8.330 64.730 ;
        RECT 8.520 64.560 8.690 64.730 ;
        RECT 8.880 64.560 9.050 64.730 ;
        RECT 9.240 64.560 9.410 64.730 ;
        RECT 10.580 64.610 10.750 64.780 ;
        RECT 10.940 64.610 11.110 64.780 ;
        RECT 11.380 64.610 11.550 64.780 ;
        RECT 12.120 64.560 12.290 64.730 ;
        RECT 12.480 64.560 12.650 64.730 ;
        RECT 12.840 64.560 13.010 64.730 ;
        RECT 13.690 64.560 13.860 64.730 ;
        RECT 14.050 64.560 14.220 64.730 ;
        RECT 14.900 64.610 15.070 64.780 ;
        RECT 15.260 64.610 15.430 64.780 ;
        RECT 15.700 64.610 15.870 64.780 ;
        RECT 17.010 64.560 17.180 64.730 ;
        RECT 17.370 64.560 17.540 64.730 ;
        RECT 17.730 64.560 17.900 64.730 ;
        RECT 18.090 64.560 18.260 64.730 ;
        RECT 20.180 64.610 20.350 64.780 ;
        RECT 20.540 64.610 20.710 64.780 ;
        RECT 20.980 64.610 21.150 64.780 ;
        RECT 22.260 64.560 22.430 64.730 ;
        RECT 22.620 64.560 22.790 64.730 ;
        RECT 24.650 64.560 24.820 64.730 ;
        RECT 27.080 64.560 27.250 64.730 ;
        RECT 27.440 64.560 27.610 64.730 ;
        RECT 27.800 64.560 27.970 64.730 ;
        RECT 29.420 64.560 29.590 64.730 ;
        RECT 29.780 64.560 29.950 64.730 ;
        RECT 30.140 64.560 30.310 64.730 ;
        RECT 32.120 64.560 32.290 64.730 ;
        RECT 32.480 64.560 32.650 64.730 ;
        RECT 32.840 64.560 33.010 64.730 ;
        RECT 33.870 64.560 34.040 64.730 ;
        RECT 34.230 64.560 34.400 64.730 ;
        RECT 34.590 64.560 34.760 64.730 ;
        RECT 35.400 64.560 35.570 64.730 ;
        RECT 35.760 64.560 35.930 64.730 ;
        RECT 36.120 64.560 36.290 64.730 ;
        RECT 37.460 64.610 37.630 64.780 ;
        RECT 37.820 64.610 37.990 64.780 ;
        RECT 38.260 64.610 38.430 64.780 ;
        RECT 39.000 64.560 39.170 64.730 ;
        RECT 39.360 64.560 39.530 64.730 ;
        RECT 39.720 64.560 39.890 64.730 ;
        RECT 40.560 64.560 40.730 64.730 ;
        RECT 40.920 64.560 41.090 64.730 ;
        RECT 41.280 64.560 41.450 64.730 ;
        RECT 42.200 64.560 42.370 64.730 ;
        RECT 42.560 64.560 42.730 64.730 ;
        RECT 42.920 64.560 43.090 64.730 ;
        RECT 44.180 64.610 44.350 64.780 ;
        RECT 44.540 64.610 44.710 64.780 ;
        RECT 44.980 64.610 45.150 64.780 ;
        RECT 47.220 64.560 47.390 64.730 ;
        RECT 47.580 64.560 47.750 64.730 ;
        RECT 49.610 64.560 49.780 64.730 ;
        RECT 52.040 64.560 52.210 64.730 ;
        RECT 52.400 64.560 52.570 64.730 ;
        RECT 52.760 64.560 52.930 64.730 ;
        RECT 54.380 64.560 54.550 64.730 ;
        RECT 54.740 64.560 54.910 64.730 ;
        RECT 55.100 64.560 55.270 64.730 ;
        RECT 57.080 64.560 57.250 64.730 ;
        RECT 57.440 64.560 57.610 64.730 ;
        RECT 57.800 64.560 57.970 64.730 ;
        RECT 58.830 64.560 59.000 64.730 ;
        RECT 59.190 64.560 59.360 64.730 ;
        RECT 59.550 64.560 59.720 64.730 ;
        RECT 60.360 64.560 60.530 64.730 ;
        RECT 60.720 64.560 60.890 64.730 ;
        RECT 61.080 64.560 61.250 64.730 ;
        RECT 62.420 64.610 62.590 64.780 ;
        RECT 62.780 64.610 62.950 64.780 ;
        RECT 63.220 64.610 63.390 64.780 ;
        RECT 63.960 64.560 64.130 64.730 ;
        RECT 64.320 64.560 64.490 64.730 ;
        RECT 64.680 64.560 64.850 64.730 ;
        RECT 65.530 64.560 65.700 64.730 ;
        RECT 65.890 64.560 66.060 64.730 ;
        RECT 66.740 64.610 66.910 64.780 ;
        RECT 67.100 64.610 67.270 64.780 ;
        RECT 67.540 64.610 67.710 64.780 ;
        RECT 68.860 64.560 69.030 64.730 ;
        RECT 69.220 64.560 69.390 64.730 ;
        RECT 71.600 64.560 71.770 64.730 ;
        RECT 71.960 64.560 72.130 64.730 ;
        RECT 72.320 64.560 72.490 64.730 ;
        RECT 72.680 64.560 72.850 64.730 ;
        RECT 73.940 64.610 74.110 64.780 ;
        RECT 74.300 64.610 74.470 64.780 ;
        RECT 74.740 64.610 74.910 64.780 ;
        RECT 75.480 64.560 75.650 64.730 ;
        RECT 75.840 64.560 76.010 64.730 ;
        RECT 76.200 64.560 76.370 64.730 ;
        RECT 77.040 64.560 77.210 64.730 ;
        RECT 77.400 64.560 77.570 64.730 ;
        RECT 77.760 64.560 77.930 64.730 ;
        RECT 78.680 64.560 78.850 64.730 ;
        RECT 79.040 64.560 79.210 64.730 ;
        RECT 79.400 64.560 79.570 64.730 ;
        RECT 80.660 64.610 80.830 64.780 ;
        RECT 81.020 64.610 81.190 64.780 ;
        RECT 81.460 64.610 81.630 64.780 ;
        RECT 82.200 64.560 82.370 64.730 ;
        RECT 82.560 64.560 82.730 64.730 ;
        RECT 84.020 64.610 84.190 64.780 ;
        RECT 84.380 64.610 84.550 64.780 ;
        RECT 84.820 64.610 84.990 64.780 ;
        RECT 85.540 64.560 85.710 64.730 ;
        RECT 85.900 64.560 86.070 64.730 ;
        RECT 86.260 64.560 86.430 64.730 ;
        RECT 86.620 64.560 86.790 64.730 ;
        RECT 87.780 64.560 87.950 64.730 ;
        RECT 88.140 64.560 88.310 64.730 ;
        RECT 88.500 64.560 88.670 64.730 ;
        RECT 88.860 64.560 89.030 64.730 ;
        RECT 89.780 64.610 89.950 64.780 ;
        RECT 90.140 64.610 90.310 64.780 ;
        RECT 90.580 64.610 90.750 64.780 ;
        RECT 91.800 64.560 91.970 64.730 ;
        RECT 92.160 64.560 92.330 64.730 ;
        RECT 92.520 64.560 92.690 64.730 ;
        RECT 93.360 64.560 93.530 64.730 ;
        RECT 93.720 64.560 93.890 64.730 ;
        RECT 94.080 64.560 94.250 64.730 ;
        RECT 95.000 64.560 95.170 64.730 ;
        RECT 95.360 64.560 95.530 64.730 ;
        RECT 95.720 64.560 95.890 64.730 ;
        RECT 96.980 64.610 97.150 64.780 ;
        RECT 97.340 64.610 97.510 64.780 ;
        RECT 97.780 64.610 97.950 64.780 ;
        RECT 99.090 64.560 99.260 64.730 ;
        RECT 99.450 64.560 99.620 64.730 ;
        RECT 99.810 64.560 99.980 64.730 ;
        RECT 100.170 64.560 100.340 64.730 ;
        RECT 102.470 64.610 102.640 64.780 ;
        RECT 102.910 64.610 103.080 64.780 ;
        RECT 103.320 64.610 103.490 64.780 ;
        RECT 103.750 64.610 103.920 64.780 ;
        RECT 104.190 64.610 104.360 64.780 ;
        RECT 104.600 64.610 104.770 64.780 ;
        RECT 106.740 64.560 106.910 64.730 ;
        RECT 107.100 64.560 107.270 64.730 ;
        RECT 109.130 64.560 109.300 64.730 ;
        RECT 111.560 64.560 111.730 64.730 ;
        RECT 111.920 64.560 112.090 64.730 ;
        RECT 112.280 64.560 112.450 64.730 ;
        RECT 113.900 64.560 114.070 64.730 ;
        RECT 114.260 64.560 114.430 64.730 ;
        RECT 114.620 64.560 114.790 64.730 ;
        RECT 116.600 64.560 116.770 64.730 ;
        RECT 116.960 64.560 117.130 64.730 ;
        RECT 117.320 64.560 117.490 64.730 ;
        RECT 118.350 64.560 118.520 64.730 ;
        RECT 118.710 64.560 118.880 64.730 ;
        RECT 119.070 64.560 119.240 64.730 ;
        RECT 119.880 64.560 120.050 64.730 ;
        RECT 120.240 64.560 120.410 64.730 ;
        RECT 120.600 64.560 120.770 64.730 ;
        RECT 121.940 64.610 122.110 64.780 ;
        RECT 122.300 64.610 122.470 64.780 ;
        RECT 122.740 64.610 122.910 64.780 ;
        RECT 124.020 64.560 124.190 64.730 ;
        RECT 124.380 64.560 124.550 64.730 ;
        RECT 126.410 64.560 126.580 64.730 ;
        RECT 128.840 64.560 129.010 64.730 ;
        RECT 129.200 64.560 129.370 64.730 ;
        RECT 129.560 64.560 129.730 64.730 ;
        RECT 131.180 64.560 131.350 64.730 ;
        RECT 131.540 64.560 131.710 64.730 ;
        RECT 131.900 64.560 132.070 64.730 ;
        RECT 133.880 64.560 134.050 64.730 ;
        RECT 134.240 64.560 134.410 64.730 ;
        RECT 134.600 64.560 134.770 64.730 ;
        RECT 135.630 64.560 135.800 64.730 ;
        RECT 135.990 64.560 136.160 64.730 ;
        RECT 136.350 64.560 136.520 64.730 ;
        RECT 137.160 64.560 137.330 64.730 ;
        RECT 137.520 64.560 137.690 64.730 ;
        RECT 137.880 64.560 138.050 64.730 ;
        RECT 139.220 64.610 139.390 64.780 ;
        RECT 139.580 64.610 139.750 64.780 ;
        RECT 140.020 64.610 140.190 64.780 ;
        RECT 6.260 57.320 6.430 57.490 ;
        RECT 6.620 57.320 6.790 57.490 ;
        RECT 7.060 57.320 7.230 57.490 ;
        RECT 8.340 57.370 8.510 57.540 ;
        RECT 8.700 57.370 8.870 57.540 ;
        RECT 10.730 57.370 10.900 57.540 ;
        RECT 13.160 57.370 13.330 57.540 ;
        RECT 13.520 57.370 13.690 57.540 ;
        RECT 13.880 57.370 14.050 57.540 ;
        RECT 15.500 57.370 15.670 57.540 ;
        RECT 15.860 57.370 16.030 57.540 ;
        RECT 16.220 57.370 16.390 57.540 ;
        RECT 18.200 57.370 18.370 57.540 ;
        RECT 18.560 57.370 18.730 57.540 ;
        RECT 18.920 57.370 19.090 57.540 ;
        RECT 19.950 57.370 20.120 57.540 ;
        RECT 20.310 57.370 20.480 57.540 ;
        RECT 20.670 57.370 20.840 57.540 ;
        RECT 21.480 57.370 21.650 57.540 ;
        RECT 21.840 57.370 22.010 57.540 ;
        RECT 22.200 57.370 22.370 57.540 ;
        RECT 23.540 57.320 23.710 57.490 ;
        RECT 23.900 57.320 24.070 57.490 ;
        RECT 24.340 57.320 24.510 57.490 ;
        RECT 25.700 57.370 25.870 57.540 ;
        RECT 26.060 57.370 26.230 57.540 ;
        RECT 27.860 57.320 28.030 57.490 ;
        RECT 28.220 57.320 28.390 57.490 ;
        RECT 28.660 57.320 28.830 57.490 ;
        RECT 29.400 57.370 29.570 57.540 ;
        RECT 29.760 57.370 29.930 57.540 ;
        RECT 30.120 57.370 30.290 57.540 ;
        RECT 30.960 57.370 31.130 57.540 ;
        RECT 31.320 57.370 31.490 57.540 ;
        RECT 31.680 57.370 31.850 57.540 ;
        RECT 32.600 57.370 32.770 57.540 ;
        RECT 32.960 57.370 33.130 57.540 ;
        RECT 33.320 57.370 33.490 57.540 ;
        RECT 34.580 57.320 34.750 57.490 ;
        RECT 34.940 57.320 35.110 57.490 ;
        RECT 35.380 57.320 35.550 57.490 ;
        RECT 36.120 57.370 36.290 57.540 ;
        RECT 36.480 57.370 36.650 57.540 ;
        RECT 36.840 57.370 37.010 57.540 ;
        RECT 37.680 57.370 37.850 57.540 ;
        RECT 38.040 57.370 38.210 57.540 ;
        RECT 38.400 57.370 38.570 57.540 ;
        RECT 39.320 57.370 39.490 57.540 ;
        RECT 39.680 57.370 39.850 57.540 ;
        RECT 40.040 57.370 40.210 57.540 ;
        RECT 41.300 57.320 41.470 57.490 ;
        RECT 41.660 57.320 41.830 57.490 ;
        RECT 42.100 57.320 42.270 57.490 ;
        RECT 42.840 57.370 43.010 57.540 ;
        RECT 43.200 57.370 43.370 57.540 ;
        RECT 43.560 57.370 43.730 57.540 ;
        RECT 44.400 57.370 44.570 57.540 ;
        RECT 44.760 57.370 44.930 57.540 ;
        RECT 45.120 57.370 45.290 57.540 ;
        RECT 46.040 57.370 46.210 57.540 ;
        RECT 46.400 57.370 46.570 57.540 ;
        RECT 46.760 57.370 46.930 57.540 ;
        RECT 48.020 57.320 48.190 57.490 ;
        RECT 48.380 57.320 48.550 57.490 ;
        RECT 48.820 57.320 48.990 57.490 ;
        RECT 50.040 57.370 50.210 57.540 ;
        RECT 50.400 57.370 50.570 57.540 ;
        RECT 50.760 57.370 50.930 57.540 ;
        RECT 51.600 57.370 51.770 57.540 ;
        RECT 51.960 57.370 52.130 57.540 ;
        RECT 52.320 57.370 52.490 57.540 ;
        RECT 53.240 57.370 53.410 57.540 ;
        RECT 53.600 57.370 53.770 57.540 ;
        RECT 53.960 57.370 54.130 57.540 ;
        RECT 55.220 57.320 55.390 57.490 ;
        RECT 55.580 57.320 55.750 57.490 ;
        RECT 56.020 57.320 56.190 57.490 ;
        RECT 56.760 57.370 56.930 57.540 ;
        RECT 57.120 57.370 57.290 57.540 ;
        RECT 57.480 57.370 57.650 57.540 ;
        RECT 57.840 57.370 58.010 57.540 ;
        RECT 58.200 57.370 58.370 57.540 ;
        RECT 60.500 57.320 60.670 57.490 ;
        RECT 60.860 57.320 61.030 57.490 ;
        RECT 61.300 57.320 61.470 57.490 ;
        RECT 62.580 57.370 62.750 57.540 ;
        RECT 62.940 57.370 63.110 57.540 ;
        RECT 64.970 57.370 65.140 57.540 ;
        RECT 67.400 57.370 67.570 57.540 ;
        RECT 67.760 57.370 67.930 57.540 ;
        RECT 68.120 57.370 68.290 57.540 ;
        RECT 69.740 57.370 69.910 57.540 ;
        RECT 70.100 57.370 70.270 57.540 ;
        RECT 70.460 57.370 70.630 57.540 ;
        RECT 72.440 57.370 72.610 57.540 ;
        RECT 72.800 57.370 72.970 57.540 ;
        RECT 73.160 57.370 73.330 57.540 ;
        RECT 74.190 57.370 74.360 57.540 ;
        RECT 74.550 57.370 74.720 57.540 ;
        RECT 74.910 57.370 75.080 57.540 ;
        RECT 75.720 57.370 75.890 57.540 ;
        RECT 76.080 57.370 76.250 57.540 ;
        RECT 76.440 57.370 76.610 57.540 ;
        RECT 77.780 57.320 77.950 57.490 ;
        RECT 78.140 57.320 78.310 57.490 ;
        RECT 78.580 57.320 78.750 57.490 ;
        RECT 79.320 57.370 79.490 57.540 ;
        RECT 79.680 57.370 79.850 57.540 ;
        RECT 80.040 57.370 80.210 57.540 ;
        RECT 80.880 57.370 81.050 57.540 ;
        RECT 81.240 57.370 81.410 57.540 ;
        RECT 81.600 57.370 81.770 57.540 ;
        RECT 82.520 57.370 82.690 57.540 ;
        RECT 82.880 57.370 83.050 57.540 ;
        RECT 83.240 57.370 83.410 57.540 ;
        RECT 84.710 57.320 84.880 57.490 ;
        RECT 85.150 57.320 85.320 57.490 ;
        RECT 85.560 57.320 85.730 57.490 ;
        RECT 85.990 57.320 86.160 57.490 ;
        RECT 86.430 57.320 86.600 57.490 ;
        RECT 86.840 57.320 87.010 57.490 ;
        RECT 87.960 57.370 88.130 57.540 ;
        RECT 88.320 57.370 88.490 57.540 ;
        RECT 88.680 57.370 88.850 57.540 ;
        RECT 89.520 57.370 89.690 57.540 ;
        RECT 89.880 57.370 90.050 57.540 ;
        RECT 90.240 57.370 90.410 57.540 ;
        RECT 91.160 57.370 91.330 57.540 ;
        RECT 91.520 57.370 91.690 57.540 ;
        RECT 91.880 57.370 92.050 57.540 ;
        RECT 93.140 57.320 93.310 57.490 ;
        RECT 93.500 57.320 93.670 57.490 ;
        RECT 93.940 57.320 94.110 57.490 ;
        RECT 94.680 57.370 94.850 57.540 ;
        RECT 95.040 57.370 95.210 57.540 ;
        RECT 95.400 57.370 95.570 57.540 ;
        RECT 96.240 57.370 96.410 57.540 ;
        RECT 96.600 57.370 96.770 57.540 ;
        RECT 96.960 57.370 97.130 57.540 ;
        RECT 97.880 57.370 98.050 57.540 ;
        RECT 98.240 57.370 98.410 57.540 ;
        RECT 98.600 57.370 98.770 57.540 ;
        RECT 99.860 57.320 100.030 57.490 ;
        RECT 100.220 57.320 100.390 57.490 ;
        RECT 100.660 57.320 100.830 57.490 ;
        RECT 102.340 57.370 102.510 57.540 ;
        RECT 102.700 57.370 102.870 57.540 ;
        RECT 103.060 57.370 103.230 57.540 ;
        RECT 103.760 57.370 103.930 57.540 ;
        RECT 104.120 57.370 104.290 57.540 ;
        RECT 104.480 57.370 104.650 57.540 ;
        RECT 104.840 57.370 105.010 57.540 ;
        RECT 105.200 57.370 105.370 57.540 ;
        RECT 105.560 57.370 105.730 57.540 ;
        RECT 105.920 57.370 106.090 57.540 ;
        RECT 106.740 57.370 106.910 57.540 ;
        RECT 107.100 57.370 107.270 57.540 ;
        RECT 108.020 57.320 108.190 57.490 ;
        RECT 108.380 57.320 108.550 57.490 ;
        RECT 108.820 57.320 108.990 57.490 ;
        RECT 109.560 57.370 109.730 57.540 ;
        RECT 109.920 57.370 110.090 57.540 ;
        RECT 110.280 57.370 110.450 57.540 ;
        RECT 111.120 57.370 111.290 57.540 ;
        RECT 111.480 57.370 111.650 57.540 ;
        RECT 111.840 57.370 112.010 57.540 ;
        RECT 112.760 57.370 112.930 57.540 ;
        RECT 113.120 57.370 113.290 57.540 ;
        RECT 113.480 57.370 113.650 57.540 ;
        RECT 114.740 57.320 114.910 57.490 ;
        RECT 115.100 57.320 115.270 57.490 ;
        RECT 115.540 57.320 115.710 57.490 ;
        RECT 116.280 57.370 116.450 57.540 ;
        RECT 116.640 57.370 116.810 57.540 ;
        RECT 117.000 57.370 117.170 57.540 ;
        RECT 117.840 57.370 118.010 57.540 ;
        RECT 118.200 57.370 118.370 57.540 ;
        RECT 118.560 57.370 118.730 57.540 ;
        RECT 119.480 57.370 119.650 57.540 ;
        RECT 119.840 57.370 120.010 57.540 ;
        RECT 120.200 57.370 120.370 57.540 ;
        RECT 121.460 57.320 121.630 57.490 ;
        RECT 121.820 57.320 121.990 57.490 ;
        RECT 122.260 57.320 122.430 57.490 ;
        RECT 123.000 57.370 123.170 57.540 ;
        RECT 123.360 57.370 123.530 57.540 ;
        RECT 123.720 57.370 123.890 57.540 ;
        RECT 124.560 57.370 124.730 57.540 ;
        RECT 124.920 57.370 125.090 57.540 ;
        RECT 125.280 57.370 125.450 57.540 ;
        RECT 126.200 57.370 126.370 57.540 ;
        RECT 126.560 57.370 126.730 57.540 ;
        RECT 126.920 57.370 127.090 57.540 ;
        RECT 128.180 57.320 128.350 57.490 ;
        RECT 128.540 57.320 128.710 57.490 ;
        RECT 128.980 57.320 129.150 57.490 ;
        RECT 129.720 57.370 129.890 57.540 ;
        RECT 130.080 57.370 130.250 57.540 ;
        RECT 130.440 57.370 130.610 57.540 ;
        RECT 131.280 57.370 131.450 57.540 ;
        RECT 131.640 57.370 131.810 57.540 ;
        RECT 132.000 57.370 132.170 57.540 ;
        RECT 132.920 57.370 133.090 57.540 ;
        RECT 133.280 57.370 133.450 57.540 ;
        RECT 133.640 57.370 133.810 57.540 ;
        RECT 134.900 57.320 135.070 57.490 ;
        RECT 135.260 57.320 135.430 57.490 ;
        RECT 135.700 57.320 135.870 57.490 ;
        RECT 136.600 57.370 136.770 57.540 ;
        RECT 136.960 57.370 137.130 57.540 ;
        RECT 139.220 57.320 139.390 57.490 ;
        RECT 139.580 57.320 139.750 57.490 ;
        RECT 140.020 57.320 140.190 57.490 ;
        RECT 5.920 56.890 6.090 57.070 ;
        RECT 6.400 56.890 6.570 57.070 ;
        RECT 6.880 56.890 7.050 57.070 ;
        RECT 7.360 56.890 7.530 57.070 ;
        RECT 7.840 56.890 8.010 57.070 ;
        RECT 8.320 56.890 8.490 57.070 ;
        RECT 8.800 56.890 8.970 57.070 ;
        RECT 9.280 56.890 9.450 57.070 ;
        RECT 9.760 56.890 9.930 57.070 ;
        RECT 10.240 56.890 10.410 57.070 ;
        RECT 10.720 56.890 10.890 57.070 ;
        RECT 11.200 56.890 11.370 57.070 ;
        RECT 11.680 56.890 11.850 57.070 ;
        RECT 12.160 56.890 12.330 57.070 ;
        RECT 12.640 56.890 12.810 57.070 ;
        RECT 13.120 56.890 13.290 57.070 ;
        RECT 13.600 56.890 13.770 57.070 ;
        RECT 14.080 56.890 14.250 57.070 ;
        RECT 14.560 56.890 14.730 57.070 ;
        RECT 15.040 56.890 15.210 57.070 ;
        RECT 15.520 56.890 15.690 57.070 ;
        RECT 16.000 56.890 16.170 57.070 ;
        RECT 16.480 56.890 16.650 57.070 ;
        RECT 16.960 56.890 17.130 57.070 ;
        RECT 17.440 56.890 17.610 57.070 ;
        RECT 17.920 56.890 18.090 57.070 ;
        RECT 18.400 56.890 18.570 57.070 ;
        RECT 18.880 56.890 19.050 57.070 ;
        RECT 19.360 56.890 19.530 57.070 ;
        RECT 19.840 56.890 20.010 57.070 ;
        RECT 20.320 56.890 20.490 57.070 ;
        RECT 20.800 56.890 20.970 57.070 ;
        RECT 21.280 56.890 21.450 57.070 ;
        RECT 21.760 56.890 21.930 57.070 ;
        RECT 22.240 56.890 22.410 57.070 ;
        RECT 22.720 56.890 22.890 57.070 ;
        RECT 23.200 56.890 23.370 57.070 ;
        RECT 23.680 56.890 23.850 57.070 ;
        RECT 24.160 56.890 24.330 57.070 ;
        RECT 24.640 56.890 24.810 57.070 ;
        RECT 25.120 56.890 25.290 57.070 ;
        RECT 25.600 56.890 25.770 57.070 ;
        RECT 26.080 56.890 26.250 57.070 ;
        RECT 26.560 56.890 26.730 57.070 ;
        RECT 27.040 56.890 27.210 57.070 ;
        RECT 27.520 56.890 27.690 57.070 ;
        RECT 28.000 56.890 28.170 57.070 ;
        RECT 28.480 56.890 28.650 57.070 ;
        RECT 28.960 56.890 29.130 57.070 ;
        RECT 29.440 56.890 29.610 57.070 ;
        RECT 29.920 56.890 30.090 57.070 ;
        RECT 30.400 56.890 30.570 57.070 ;
        RECT 30.880 56.890 31.050 57.070 ;
        RECT 31.360 56.890 31.530 57.070 ;
        RECT 31.840 56.890 32.010 57.070 ;
        RECT 32.320 56.890 32.490 57.070 ;
        RECT 32.800 56.890 32.970 57.070 ;
        RECT 33.280 56.890 33.450 57.070 ;
        RECT 33.760 56.890 33.930 57.070 ;
        RECT 34.240 56.890 34.410 57.070 ;
        RECT 34.720 56.890 34.890 57.070 ;
        RECT 35.200 56.890 35.370 57.070 ;
        RECT 35.680 56.890 35.850 57.070 ;
        RECT 36.160 56.890 36.330 57.070 ;
        RECT 36.640 56.890 36.810 57.070 ;
        RECT 37.120 56.890 37.290 57.070 ;
        RECT 37.600 56.890 37.770 57.070 ;
        RECT 38.080 56.890 38.250 57.070 ;
        RECT 38.560 56.890 38.730 57.070 ;
        RECT 39.040 56.890 39.210 57.070 ;
        RECT 39.520 56.890 39.690 57.070 ;
        RECT 40.000 56.890 40.170 57.070 ;
        RECT 40.480 56.890 40.650 57.070 ;
        RECT 40.960 56.890 41.130 57.070 ;
        RECT 41.440 56.890 41.610 57.070 ;
        RECT 41.920 56.890 42.090 57.070 ;
        RECT 42.400 56.890 42.570 57.070 ;
        RECT 42.880 56.890 43.050 57.070 ;
        RECT 43.360 56.890 43.530 57.070 ;
        RECT 43.840 56.890 44.010 57.070 ;
        RECT 44.320 56.890 44.490 57.070 ;
        RECT 44.800 56.890 44.970 57.070 ;
        RECT 45.280 56.890 45.450 57.070 ;
        RECT 45.760 56.890 45.930 57.070 ;
        RECT 46.240 56.890 46.410 57.070 ;
        RECT 46.720 56.890 46.890 57.070 ;
        RECT 47.200 56.890 47.370 57.070 ;
        RECT 47.680 56.890 47.850 57.070 ;
        RECT 48.160 56.890 48.330 57.070 ;
        RECT 48.640 56.890 48.810 57.070 ;
        RECT 49.120 56.890 49.290 57.070 ;
        RECT 49.600 57.060 49.770 57.070 ;
      LAYER li1 ;
        RECT 49.440 56.890 49.920 57.060 ;
      LAYER li1 ;
        RECT 50.080 56.890 50.250 57.070 ;
        RECT 50.560 56.890 50.730 57.070 ;
        RECT 51.040 56.890 51.210 57.070 ;
        RECT 51.520 56.890 51.690 57.070 ;
        RECT 52.000 56.890 52.170 57.070 ;
        RECT 52.480 56.890 52.650 57.070 ;
        RECT 52.960 56.890 53.130 57.070 ;
        RECT 53.440 56.890 53.610 57.070 ;
        RECT 53.920 56.890 54.090 57.070 ;
        RECT 54.400 56.890 54.570 57.070 ;
        RECT 54.880 56.890 55.050 57.070 ;
        RECT 55.360 56.890 55.530 57.070 ;
        RECT 55.840 56.890 56.010 57.070 ;
        RECT 56.320 56.890 56.490 57.070 ;
        RECT 56.800 56.890 56.970 57.070 ;
        RECT 57.280 56.890 57.450 57.070 ;
        RECT 57.760 56.890 57.930 57.070 ;
        RECT 58.240 56.890 58.410 57.070 ;
        RECT 58.720 56.890 58.890 57.070 ;
        RECT 59.200 56.890 59.370 57.070 ;
        RECT 59.680 56.890 59.850 57.070 ;
        RECT 60.160 56.890 60.330 57.070 ;
        RECT 60.640 56.890 60.810 57.070 ;
        RECT 61.120 56.890 61.290 57.070 ;
        RECT 61.600 56.890 61.770 57.070 ;
        RECT 62.080 56.890 62.250 57.070 ;
        RECT 62.560 56.890 62.730 57.070 ;
        RECT 63.040 56.890 63.210 57.070 ;
        RECT 63.520 56.890 63.690 57.070 ;
        RECT 64.000 56.890 64.170 57.070 ;
        RECT 64.480 56.890 64.650 57.070 ;
        RECT 64.960 56.890 65.130 57.070 ;
        RECT 65.440 56.890 65.610 57.070 ;
        RECT 65.920 56.890 66.090 57.070 ;
        RECT 66.400 56.890 66.570 57.070 ;
        RECT 66.880 56.890 67.050 57.070 ;
        RECT 67.360 56.890 67.530 57.070 ;
        RECT 67.840 56.890 68.010 57.070 ;
        RECT 68.320 56.890 68.490 57.070 ;
        RECT 68.800 56.890 68.970 57.070 ;
        RECT 69.280 56.890 69.450 57.070 ;
        RECT 69.760 56.890 69.930 57.070 ;
        RECT 70.240 56.890 70.410 57.070 ;
        RECT 70.720 56.890 70.890 57.070 ;
        RECT 71.200 56.890 71.370 57.070 ;
        RECT 71.680 56.890 71.850 57.070 ;
        RECT 72.160 56.890 72.330 57.070 ;
        RECT 72.640 56.890 72.810 57.070 ;
        RECT 73.120 56.890 73.290 57.070 ;
        RECT 73.600 56.890 73.770 57.070 ;
        RECT 74.080 56.890 74.250 57.070 ;
        RECT 74.560 56.890 74.730 57.070 ;
        RECT 75.040 56.890 75.210 57.070 ;
        RECT 75.520 56.890 75.690 57.070 ;
        RECT 76.000 56.890 76.170 57.070 ;
        RECT 76.480 56.890 76.650 57.070 ;
        RECT 76.960 56.890 77.130 57.070 ;
        RECT 77.440 56.890 77.610 57.070 ;
        RECT 77.920 56.890 78.090 57.070 ;
        RECT 78.400 56.890 78.570 57.070 ;
        RECT 78.880 56.890 79.050 57.070 ;
        RECT 79.360 56.890 79.530 57.070 ;
        RECT 79.840 56.890 80.010 57.070 ;
        RECT 80.320 56.890 80.490 57.070 ;
        RECT 80.800 56.890 80.970 57.070 ;
        RECT 81.280 56.890 81.450 57.070 ;
        RECT 81.760 56.890 81.930 57.070 ;
        RECT 82.240 56.890 82.410 57.070 ;
        RECT 82.720 56.890 82.890 57.070 ;
        RECT 83.200 56.890 83.370 57.070 ;
        RECT 83.680 56.890 83.850 57.070 ;
        RECT 84.160 56.890 84.330 57.070 ;
        RECT 84.640 56.890 84.810 57.070 ;
        RECT 85.120 56.890 85.290 57.070 ;
        RECT 85.600 56.890 85.770 57.070 ;
        RECT 86.080 56.890 86.250 57.070 ;
        RECT 86.560 56.890 86.730 57.070 ;
        RECT 87.040 56.890 87.210 57.070 ;
        RECT 87.520 56.890 87.690 57.070 ;
        RECT 88.000 56.890 88.170 57.070 ;
        RECT 88.480 56.890 88.650 57.070 ;
        RECT 88.960 56.890 89.130 57.070 ;
        RECT 89.440 56.890 89.610 57.070 ;
        RECT 89.920 56.890 90.090 57.070 ;
        RECT 90.400 56.890 90.570 57.070 ;
        RECT 90.880 56.890 91.050 57.070 ;
        RECT 91.360 56.890 91.530 57.070 ;
        RECT 91.840 56.890 92.010 57.070 ;
        RECT 92.320 56.890 92.490 57.070 ;
        RECT 92.800 56.890 92.970 57.070 ;
        RECT 93.280 56.890 93.450 57.070 ;
        RECT 93.760 56.890 93.930 57.070 ;
        RECT 94.240 56.890 94.410 57.070 ;
        RECT 94.720 56.890 94.890 57.070 ;
        RECT 95.200 56.890 95.370 57.070 ;
        RECT 95.680 56.890 95.850 57.070 ;
        RECT 96.160 56.890 96.330 57.070 ;
        RECT 96.640 56.890 96.810 57.070 ;
        RECT 97.120 56.890 97.290 57.070 ;
        RECT 97.600 56.890 97.770 57.070 ;
        RECT 98.080 56.890 98.250 57.070 ;
        RECT 98.560 56.890 98.730 57.070 ;
        RECT 99.040 56.890 99.210 57.070 ;
        RECT 99.520 56.890 99.690 57.070 ;
        RECT 100.000 56.890 100.170 57.070 ;
        RECT 100.480 56.890 100.650 57.070 ;
        RECT 100.960 56.890 101.130 57.070 ;
        RECT 101.440 56.890 101.610 57.070 ;
      LAYER li1 ;
        RECT 101.760 57.060 102.240 57.070 ;
      LAYER li1 ;
        RECT 101.920 56.890 102.090 57.060 ;
        RECT 102.400 56.890 102.570 57.070 ;
        RECT 102.880 56.890 103.050 57.070 ;
        RECT 103.360 56.890 103.530 57.070 ;
        RECT 103.840 56.890 104.010 57.070 ;
        RECT 104.320 56.890 104.490 57.070 ;
        RECT 104.800 56.890 104.970 57.070 ;
        RECT 105.280 56.890 105.450 57.070 ;
        RECT 105.760 56.890 105.930 57.070 ;
        RECT 106.240 56.890 106.410 57.070 ;
        RECT 106.720 56.890 106.890 57.070 ;
        RECT 107.200 56.890 107.370 57.070 ;
        RECT 107.680 56.890 107.850 57.070 ;
        RECT 108.160 56.890 108.330 57.070 ;
        RECT 108.640 56.890 108.810 57.070 ;
        RECT 109.120 56.890 109.290 57.070 ;
        RECT 109.600 56.890 109.770 57.070 ;
        RECT 110.080 56.890 110.250 57.070 ;
        RECT 110.560 56.890 110.730 57.070 ;
        RECT 111.040 56.890 111.210 57.070 ;
        RECT 111.520 56.890 111.690 57.070 ;
        RECT 112.000 56.890 112.170 57.070 ;
        RECT 112.480 56.890 112.650 57.070 ;
        RECT 112.960 56.890 113.130 57.070 ;
        RECT 113.440 56.890 113.610 57.070 ;
        RECT 113.920 56.890 114.090 57.070 ;
        RECT 114.400 56.890 114.570 57.070 ;
        RECT 114.880 56.890 115.050 57.070 ;
        RECT 115.360 56.890 115.530 57.070 ;
      LAYER li1 ;
        RECT 115.680 57.060 116.160 57.070 ;
      LAYER li1 ;
        RECT 115.840 56.890 116.010 57.060 ;
        RECT 116.320 56.890 116.490 57.070 ;
        RECT 116.800 56.890 116.970 57.070 ;
        RECT 117.280 56.890 117.450 57.070 ;
        RECT 117.760 56.890 117.930 57.070 ;
        RECT 118.240 56.890 118.410 57.070 ;
        RECT 118.720 56.890 118.890 57.070 ;
        RECT 119.200 56.890 119.370 57.070 ;
        RECT 119.680 56.890 119.850 57.070 ;
        RECT 120.160 56.890 120.330 57.070 ;
        RECT 120.640 56.890 120.810 57.070 ;
        RECT 121.120 56.890 121.290 57.070 ;
        RECT 121.600 56.890 121.770 57.070 ;
        RECT 122.080 56.890 122.250 57.070 ;
        RECT 122.560 56.890 122.730 57.070 ;
        RECT 123.040 56.890 123.210 57.070 ;
        RECT 123.520 56.890 123.690 57.070 ;
        RECT 124.000 56.890 124.170 57.070 ;
        RECT 124.480 56.890 124.650 57.070 ;
        RECT 124.960 56.890 125.130 57.070 ;
        RECT 125.440 56.890 125.610 57.070 ;
        RECT 125.920 56.890 126.090 57.070 ;
        RECT 126.400 56.890 126.570 57.070 ;
        RECT 126.880 56.890 127.050 57.070 ;
        RECT 127.360 56.890 127.530 57.070 ;
        RECT 127.840 56.890 128.010 57.070 ;
        RECT 128.320 56.890 128.490 57.070 ;
        RECT 128.800 56.890 128.970 57.070 ;
        RECT 129.280 56.890 129.450 57.070 ;
        RECT 129.760 56.890 129.930 57.070 ;
        RECT 130.240 56.890 130.410 57.070 ;
        RECT 130.720 56.890 130.890 57.070 ;
        RECT 131.200 56.890 131.370 57.070 ;
        RECT 131.680 56.890 131.850 57.070 ;
        RECT 132.160 56.890 132.330 57.070 ;
        RECT 132.640 56.890 132.810 57.070 ;
        RECT 133.120 56.890 133.290 57.070 ;
        RECT 133.600 56.890 133.770 57.070 ;
        RECT 134.080 56.890 134.250 57.070 ;
        RECT 134.560 56.890 134.730 57.070 ;
        RECT 135.040 56.890 135.210 57.070 ;
        RECT 135.520 56.890 135.690 57.070 ;
        RECT 136.000 56.890 136.170 57.070 ;
        RECT 136.480 56.890 136.650 57.070 ;
        RECT 136.960 56.890 137.130 57.070 ;
        RECT 137.440 56.890 137.610 57.070 ;
        RECT 137.920 56.890 138.090 57.070 ;
        RECT 138.400 56.890 138.570 57.070 ;
        RECT 138.880 56.890 139.050 57.070 ;
        RECT 139.360 56.890 139.530 57.070 ;
        RECT 139.840 56.890 140.010 57.070 ;
        RECT 140.320 56.890 140.490 57.070 ;
        RECT 140.800 56.890 140.970 57.070 ;
        RECT 141.280 56.890 141.450 57.070 ;
        RECT 141.760 57.060 141.930 57.070 ;
      LAYER li1 ;
        RECT 141.600 56.890 142.080 57.060 ;
      LAYER li1 ;
        RECT 5.880 56.420 6.050 56.590 ;
        RECT 6.240 56.420 6.410 56.590 ;
        RECT 7.700 56.470 7.870 56.640 ;
        RECT 8.060 56.470 8.230 56.640 ;
        RECT 8.500 56.470 8.670 56.640 ;
        RECT 9.240 56.420 9.410 56.590 ;
        RECT 9.600 56.420 9.770 56.590 ;
        RECT 11.060 56.470 11.230 56.640 ;
        RECT 11.420 56.470 11.590 56.640 ;
        RECT 11.860 56.470 12.030 56.640 ;
        RECT 13.220 56.420 13.390 56.590 ;
        RECT 13.580 56.420 13.750 56.590 ;
        RECT 15.380 56.470 15.550 56.640 ;
        RECT 15.740 56.470 15.910 56.640 ;
        RECT 16.180 56.470 16.350 56.640 ;
        RECT 16.920 56.420 17.090 56.590 ;
        RECT 17.280 56.420 17.450 56.590 ;
        RECT 17.640 56.420 17.810 56.590 ;
        RECT 18.000 56.420 18.170 56.590 ;
        RECT 18.360 56.420 18.530 56.590 ;
        RECT 20.660 56.470 20.830 56.640 ;
        RECT 21.020 56.470 21.190 56.640 ;
        RECT 21.460 56.470 21.630 56.640 ;
        RECT 22.180 56.420 22.350 56.590 ;
        RECT 22.540 56.420 22.710 56.590 ;
        RECT 22.900 56.420 23.070 56.590 ;
        RECT 23.260 56.420 23.430 56.590 ;
        RECT 24.420 56.420 24.590 56.590 ;
        RECT 24.780 56.420 24.950 56.590 ;
        RECT 25.140 56.420 25.310 56.590 ;
        RECT 25.500 56.420 25.670 56.590 ;
        RECT 26.420 56.470 26.590 56.640 ;
        RECT 26.780 56.470 26.950 56.640 ;
        RECT 27.220 56.470 27.390 56.640 ;
        RECT 27.960 56.420 28.130 56.590 ;
        RECT 28.320 56.420 28.490 56.590 ;
        RECT 28.680 56.420 28.850 56.590 ;
        RECT 29.520 56.420 29.690 56.590 ;
        RECT 29.880 56.420 30.050 56.590 ;
        RECT 30.240 56.420 30.410 56.590 ;
        RECT 31.160 56.420 31.330 56.590 ;
        RECT 31.520 56.420 31.690 56.590 ;
        RECT 31.880 56.420 32.050 56.590 ;
        RECT 33.140 56.470 33.310 56.640 ;
        RECT 33.500 56.470 33.670 56.640 ;
        RECT 33.940 56.470 34.110 56.640 ;
        RECT 34.680 56.420 34.850 56.590 ;
        RECT 35.040 56.420 35.210 56.590 ;
        RECT 35.400 56.420 35.570 56.590 ;
        RECT 36.240 56.420 36.410 56.590 ;
        RECT 36.600 56.420 36.770 56.590 ;
        RECT 36.960 56.420 37.130 56.590 ;
        RECT 37.880 56.420 38.050 56.590 ;
        RECT 38.240 56.420 38.410 56.590 ;
        RECT 38.600 56.420 38.770 56.590 ;
        RECT 39.860 56.470 40.030 56.640 ;
        RECT 40.220 56.470 40.390 56.640 ;
        RECT 40.660 56.470 40.830 56.640 ;
        RECT 41.400 56.420 41.570 56.590 ;
        RECT 41.760 56.420 41.930 56.590 ;
        RECT 42.120 56.420 42.290 56.590 ;
        RECT 42.960 56.420 43.130 56.590 ;
        RECT 43.320 56.420 43.490 56.590 ;
        RECT 43.680 56.420 43.850 56.590 ;
        RECT 44.600 56.420 44.770 56.590 ;
        RECT 44.960 56.420 45.130 56.590 ;
        RECT 45.320 56.420 45.490 56.590 ;
        RECT 46.580 56.470 46.750 56.640 ;
        RECT 46.940 56.470 47.110 56.640 ;
        RECT 47.380 56.470 47.550 56.640 ;
        RECT 48.120 56.420 48.290 56.590 ;
        RECT 48.480 56.420 48.650 56.590 ;
        RECT 48.840 56.420 49.010 56.590 ;
        RECT 49.680 56.420 49.850 56.590 ;
        RECT 50.040 56.420 50.210 56.590 ;
        RECT 50.400 56.420 50.570 56.590 ;
        RECT 51.320 56.420 51.490 56.590 ;
        RECT 51.680 56.420 51.850 56.590 ;
        RECT 52.040 56.420 52.210 56.590 ;
        RECT 53.300 56.470 53.470 56.640 ;
        RECT 53.660 56.470 53.830 56.640 ;
        RECT 54.100 56.470 54.270 56.640 ;
        RECT 54.840 56.420 55.010 56.590 ;
        RECT 55.200 56.420 55.370 56.590 ;
        RECT 55.560 56.420 55.730 56.590 ;
        RECT 56.400 56.420 56.570 56.590 ;
        RECT 56.760 56.420 56.930 56.590 ;
        RECT 57.120 56.420 57.290 56.590 ;
        RECT 58.040 56.420 58.210 56.590 ;
        RECT 58.400 56.420 58.570 56.590 ;
        RECT 58.760 56.420 58.930 56.590 ;
        RECT 60.020 56.470 60.190 56.640 ;
        RECT 60.380 56.470 60.550 56.640 ;
        RECT 60.820 56.470 60.990 56.640 ;
        RECT 61.560 56.420 61.730 56.590 ;
        RECT 61.920 56.420 62.090 56.590 ;
        RECT 62.280 56.420 62.450 56.590 ;
        RECT 63.120 56.420 63.290 56.590 ;
        RECT 63.480 56.420 63.650 56.590 ;
        RECT 63.840 56.420 64.010 56.590 ;
        RECT 64.760 56.420 64.930 56.590 ;
        RECT 65.120 56.420 65.290 56.590 ;
        RECT 65.480 56.420 65.650 56.590 ;
        RECT 66.740 56.470 66.910 56.640 ;
        RECT 67.100 56.470 67.270 56.640 ;
        RECT 67.540 56.470 67.710 56.640 ;
        RECT 68.280 56.420 68.450 56.590 ;
        RECT 68.640 56.420 68.810 56.590 ;
        RECT 69.000 56.420 69.170 56.590 ;
        RECT 69.840 56.420 70.010 56.590 ;
        RECT 70.200 56.420 70.370 56.590 ;
        RECT 70.560 56.420 70.730 56.590 ;
        RECT 71.480 56.420 71.650 56.590 ;
        RECT 71.840 56.420 72.010 56.590 ;
        RECT 72.200 56.420 72.370 56.590 ;
        RECT 73.460 56.470 73.630 56.640 ;
        RECT 73.820 56.470 73.990 56.640 ;
        RECT 74.260 56.470 74.430 56.640 ;
        RECT 75.000 56.420 75.170 56.590 ;
        RECT 75.360 56.420 75.530 56.590 ;
        RECT 75.720 56.420 75.890 56.590 ;
        RECT 76.560 56.420 76.730 56.590 ;
        RECT 76.920 56.420 77.090 56.590 ;
        RECT 77.280 56.420 77.450 56.590 ;
        RECT 78.200 56.420 78.370 56.590 ;
        RECT 78.560 56.420 78.730 56.590 ;
        RECT 78.920 56.420 79.090 56.590 ;
        RECT 80.180 56.470 80.350 56.640 ;
        RECT 80.540 56.470 80.710 56.640 ;
        RECT 80.980 56.470 81.150 56.640 ;
        RECT 82.680 56.420 82.850 56.590 ;
        RECT 83.040 56.420 83.210 56.590 ;
        RECT 83.400 56.420 83.570 56.590 ;
        RECT 84.240 56.420 84.410 56.590 ;
        RECT 84.600 56.420 84.770 56.590 ;
        RECT 84.960 56.420 85.130 56.590 ;
        RECT 85.880 56.420 86.050 56.590 ;
        RECT 86.240 56.420 86.410 56.590 ;
        RECT 86.600 56.420 86.770 56.590 ;
        RECT 87.860 56.470 88.030 56.640 ;
        RECT 88.220 56.470 88.390 56.640 ;
        RECT 88.660 56.470 88.830 56.640 ;
        RECT 89.380 56.420 89.550 56.590 ;
        RECT 89.740 56.420 89.910 56.590 ;
        RECT 90.100 56.420 90.270 56.590 ;
        RECT 90.460 56.420 90.630 56.590 ;
        RECT 91.620 56.420 91.790 56.590 ;
        RECT 91.980 56.420 92.150 56.590 ;
        RECT 92.340 56.420 92.510 56.590 ;
        RECT 92.700 56.420 92.870 56.590 ;
        RECT 93.620 56.470 93.790 56.640 ;
        RECT 93.980 56.470 94.150 56.640 ;
        RECT 94.420 56.470 94.590 56.640 ;
        RECT 97.210 56.420 97.380 56.590 ;
        RECT 97.570 56.420 97.740 56.590 ;
        RECT 97.930 56.420 98.100 56.590 ;
        RECT 99.380 56.470 99.550 56.640 ;
        RECT 99.740 56.470 99.910 56.640 ;
        RECT 100.180 56.470 100.350 56.640 ;
        RECT 102.360 56.420 102.530 56.590 ;
        RECT 102.720 56.420 102.890 56.590 ;
        RECT 103.080 56.420 103.250 56.590 ;
        RECT 103.920 56.420 104.090 56.590 ;
        RECT 104.280 56.420 104.450 56.590 ;
        RECT 104.640 56.420 104.810 56.590 ;
        RECT 105.560 56.420 105.730 56.590 ;
        RECT 105.920 56.420 106.090 56.590 ;
        RECT 106.280 56.420 106.450 56.590 ;
        RECT 107.540 56.470 107.710 56.640 ;
        RECT 107.900 56.470 108.070 56.640 ;
        RECT 108.340 56.470 108.510 56.640 ;
        RECT 109.080 56.420 109.250 56.590 ;
        RECT 109.440 56.420 109.610 56.590 ;
        RECT 109.800 56.420 109.970 56.590 ;
        RECT 110.640 56.420 110.810 56.590 ;
        RECT 111.000 56.420 111.170 56.590 ;
        RECT 111.360 56.420 111.530 56.590 ;
        RECT 112.280 56.420 112.450 56.590 ;
        RECT 112.640 56.420 112.810 56.590 ;
        RECT 113.000 56.420 113.170 56.590 ;
        RECT 114.260 56.470 114.430 56.640 ;
        RECT 114.620 56.470 114.790 56.640 ;
        RECT 115.060 56.470 115.230 56.640 ;
        RECT 116.280 56.420 116.450 56.590 ;
        RECT 116.640 56.420 116.810 56.590 ;
        RECT 117.000 56.420 117.170 56.590 ;
        RECT 117.840 56.420 118.010 56.590 ;
        RECT 118.200 56.420 118.370 56.590 ;
        RECT 118.560 56.420 118.730 56.590 ;
        RECT 119.480 56.420 119.650 56.590 ;
        RECT 119.840 56.420 120.010 56.590 ;
        RECT 120.200 56.420 120.370 56.590 ;
        RECT 121.460 56.470 121.630 56.640 ;
        RECT 121.820 56.470 121.990 56.640 ;
        RECT 122.260 56.470 122.430 56.640 ;
        RECT 123.000 56.420 123.170 56.590 ;
        RECT 123.360 56.420 123.530 56.590 ;
        RECT 123.720 56.420 123.890 56.590 ;
        RECT 124.560 56.420 124.730 56.590 ;
        RECT 124.920 56.420 125.090 56.590 ;
        RECT 125.280 56.420 125.450 56.590 ;
        RECT 126.200 56.420 126.370 56.590 ;
        RECT 126.560 56.420 126.730 56.590 ;
        RECT 126.920 56.420 127.090 56.590 ;
        RECT 128.180 56.470 128.350 56.640 ;
        RECT 128.540 56.470 128.710 56.640 ;
        RECT 128.980 56.470 129.150 56.640 ;
        RECT 129.720 56.420 129.890 56.590 ;
        RECT 130.080 56.420 130.250 56.590 ;
        RECT 130.440 56.420 130.610 56.590 ;
        RECT 131.280 56.420 131.450 56.590 ;
        RECT 131.640 56.420 131.810 56.590 ;
        RECT 132.000 56.420 132.170 56.590 ;
        RECT 132.920 56.420 133.090 56.590 ;
        RECT 133.280 56.420 133.450 56.590 ;
        RECT 133.640 56.420 133.810 56.590 ;
        RECT 134.900 56.470 135.070 56.640 ;
        RECT 135.260 56.470 135.430 56.640 ;
        RECT 135.700 56.470 135.870 56.640 ;
        RECT 136.420 56.420 136.590 56.590 ;
        RECT 136.780 56.420 136.950 56.590 ;
        RECT 137.140 56.420 137.310 56.590 ;
        RECT 137.500 56.420 137.670 56.590 ;
        RECT 138.660 56.420 138.830 56.590 ;
        RECT 139.020 56.420 139.190 56.590 ;
        RECT 139.380 56.420 139.550 56.590 ;
        RECT 139.740 56.420 139.910 56.590 ;
        RECT 140.660 56.470 140.830 56.640 ;
        RECT 141.020 56.470 141.190 56.640 ;
        RECT 141.460 56.470 141.630 56.640 ;
        RECT 6.260 49.180 6.430 49.350 ;
        RECT 6.620 49.180 6.790 49.350 ;
        RECT 7.060 49.180 7.230 49.350 ;
        RECT 8.280 49.230 8.450 49.400 ;
        RECT 8.640 49.230 8.810 49.400 ;
        RECT 10.100 49.180 10.270 49.350 ;
        RECT 10.460 49.180 10.630 49.350 ;
        RECT 10.900 49.180 11.070 49.350 ;
        RECT 12.260 49.230 12.430 49.400 ;
        RECT 12.620 49.230 12.790 49.400 ;
        RECT 14.420 49.180 14.590 49.350 ;
        RECT 14.780 49.180 14.950 49.350 ;
        RECT 15.220 49.180 15.390 49.350 ;
        RECT 15.960 49.230 16.130 49.400 ;
        RECT 16.320 49.230 16.490 49.400 ;
        RECT 16.680 49.230 16.850 49.400 ;
        RECT 17.530 49.230 17.700 49.400 ;
        RECT 17.890 49.230 18.060 49.400 ;
        RECT 18.740 49.180 18.910 49.350 ;
        RECT 19.100 49.180 19.270 49.350 ;
        RECT 19.540 49.180 19.710 49.350 ;
        RECT 22.330 49.230 22.500 49.400 ;
        RECT 22.690 49.230 22.860 49.400 ;
        RECT 23.050 49.230 23.220 49.400 ;
        RECT 24.500 49.180 24.670 49.350 ;
        RECT 24.860 49.180 25.030 49.350 ;
        RECT 25.300 49.180 25.470 49.350 ;
        RECT 26.700 49.230 26.870 49.400 ;
        RECT 27.060 49.230 27.230 49.400 ;
        RECT 27.420 49.230 27.590 49.400 ;
        RECT 27.780 49.230 27.950 49.400 ;
        RECT 28.890 49.230 29.060 49.400 ;
        RECT 29.250 49.230 29.420 49.400 ;
        RECT 29.610 49.230 29.780 49.400 ;
        RECT 29.970 49.230 30.140 49.400 ;
        RECT 30.740 49.180 30.910 49.350 ;
        RECT 31.100 49.180 31.270 49.350 ;
        RECT 31.540 49.180 31.710 49.350 ;
        RECT 32.280 49.230 32.450 49.400 ;
        RECT 32.640 49.230 32.810 49.400 ;
        RECT 33.000 49.230 33.170 49.400 ;
        RECT 33.840 49.230 34.010 49.400 ;
        RECT 34.200 49.230 34.370 49.400 ;
        RECT 34.560 49.230 34.730 49.400 ;
        RECT 35.480 49.230 35.650 49.400 ;
        RECT 35.840 49.230 36.010 49.400 ;
        RECT 36.200 49.230 36.370 49.400 ;
        RECT 37.460 49.180 37.630 49.350 ;
        RECT 37.820 49.180 37.990 49.350 ;
        RECT 38.260 49.180 38.430 49.350 ;
        RECT 39.000 49.230 39.170 49.400 ;
        RECT 39.360 49.230 39.530 49.400 ;
        RECT 39.720 49.230 39.890 49.400 ;
        RECT 40.560 49.230 40.730 49.400 ;
        RECT 40.920 49.230 41.090 49.400 ;
        RECT 41.280 49.230 41.450 49.400 ;
        RECT 42.200 49.230 42.370 49.400 ;
        RECT 42.560 49.230 42.730 49.400 ;
        RECT 42.920 49.230 43.090 49.400 ;
        RECT 44.390 49.180 44.560 49.350 ;
        RECT 44.830 49.180 45.000 49.350 ;
        RECT 45.240 49.180 45.410 49.350 ;
        RECT 45.670 49.180 45.840 49.350 ;
        RECT 46.110 49.180 46.280 49.350 ;
        RECT 46.520 49.180 46.690 49.350 ;
        RECT 48.120 49.230 48.290 49.400 ;
        RECT 48.480 49.230 48.650 49.400 ;
        RECT 48.840 49.230 49.010 49.400 ;
        RECT 49.680 49.230 49.850 49.400 ;
        RECT 50.040 49.230 50.210 49.400 ;
        RECT 50.400 49.230 50.570 49.400 ;
        RECT 51.320 49.230 51.490 49.400 ;
        RECT 51.680 49.230 51.850 49.400 ;
        RECT 52.040 49.230 52.210 49.400 ;
        RECT 53.510 49.180 53.680 49.350 ;
        RECT 53.950 49.180 54.120 49.350 ;
        RECT 54.360 49.180 54.530 49.350 ;
        RECT 54.790 49.180 54.960 49.350 ;
        RECT 55.230 49.180 55.400 49.350 ;
        RECT 55.640 49.180 55.810 49.350 ;
        RECT 57.720 49.230 57.890 49.400 ;
        RECT 58.080 49.230 58.250 49.400 ;
        RECT 58.440 49.230 58.610 49.400 ;
        RECT 59.280 49.230 59.450 49.400 ;
        RECT 59.640 49.230 59.810 49.400 ;
        RECT 60.000 49.230 60.170 49.400 ;
        RECT 60.920 49.230 61.090 49.400 ;
        RECT 61.280 49.230 61.450 49.400 ;
        RECT 61.640 49.230 61.810 49.400 ;
        RECT 62.900 49.180 63.070 49.350 ;
        RECT 63.260 49.180 63.430 49.350 ;
        RECT 63.700 49.180 63.870 49.350 ;
        RECT 64.440 49.230 64.610 49.400 ;
        RECT 64.800 49.230 64.970 49.400 ;
        RECT 65.160 49.230 65.330 49.400 ;
        RECT 66.000 49.230 66.170 49.400 ;
        RECT 66.360 49.230 66.530 49.400 ;
        RECT 66.720 49.230 66.890 49.400 ;
        RECT 67.640 49.230 67.810 49.400 ;
        RECT 68.000 49.230 68.170 49.400 ;
        RECT 68.360 49.230 68.530 49.400 ;
        RECT 69.620 49.180 69.790 49.350 ;
        RECT 69.980 49.180 70.150 49.350 ;
        RECT 70.420 49.180 70.590 49.350 ;
        RECT 71.160 49.230 71.330 49.400 ;
        RECT 71.520 49.230 71.690 49.400 ;
        RECT 71.880 49.230 72.050 49.400 ;
        RECT 72.720 49.230 72.890 49.400 ;
        RECT 73.080 49.230 73.250 49.400 ;
        RECT 73.440 49.230 73.610 49.400 ;
        RECT 74.360 49.230 74.530 49.400 ;
        RECT 74.720 49.230 74.890 49.400 ;
        RECT 75.080 49.230 75.250 49.400 ;
        RECT 76.340 49.180 76.510 49.350 ;
        RECT 76.700 49.180 76.870 49.350 ;
        RECT 77.140 49.180 77.310 49.350 ;
        RECT 77.880 49.230 78.050 49.400 ;
        RECT 78.240 49.230 78.410 49.400 ;
        RECT 79.700 49.180 79.870 49.350 ;
        RECT 80.060 49.180 80.230 49.350 ;
        RECT 80.500 49.180 80.670 49.350 ;
        RECT 81.720 49.230 81.890 49.400 ;
        RECT 82.080 49.230 82.250 49.400 ;
        RECT 82.440 49.230 82.610 49.400 ;
        RECT 83.280 49.230 83.450 49.400 ;
        RECT 83.640 49.230 83.810 49.400 ;
        RECT 84.000 49.230 84.170 49.400 ;
        RECT 84.920 49.230 85.090 49.400 ;
        RECT 85.280 49.230 85.450 49.400 ;
        RECT 85.640 49.230 85.810 49.400 ;
        RECT 86.900 49.180 87.070 49.350 ;
        RECT 87.260 49.180 87.430 49.350 ;
        RECT 87.700 49.180 87.870 49.350 ;
        RECT 88.440 49.230 88.610 49.400 ;
        RECT 88.800 49.230 88.970 49.400 ;
        RECT 89.160 49.230 89.330 49.400 ;
        RECT 90.000 49.230 90.170 49.400 ;
        RECT 90.360 49.230 90.530 49.400 ;
        RECT 90.720 49.230 90.890 49.400 ;
        RECT 91.640 49.230 91.810 49.400 ;
        RECT 92.000 49.230 92.170 49.400 ;
        RECT 92.360 49.230 92.530 49.400 ;
        RECT 93.620 49.180 93.790 49.350 ;
        RECT 93.980 49.180 94.150 49.350 ;
        RECT 94.420 49.180 94.590 49.350 ;
        RECT 95.160 49.230 95.330 49.400 ;
        RECT 95.520 49.230 95.690 49.400 ;
        RECT 96.980 49.180 97.150 49.350 ;
        RECT 97.340 49.180 97.510 49.350 ;
        RECT 97.780 49.180 97.950 49.350 ;
        RECT 98.520 49.230 98.690 49.400 ;
        RECT 98.880 49.230 99.050 49.400 ;
        RECT 99.240 49.230 99.410 49.400 ;
        RECT 100.080 49.230 100.250 49.400 ;
        RECT 100.440 49.230 100.610 49.400 ;
        RECT 100.800 49.230 100.970 49.400 ;
        RECT 101.720 49.230 101.890 49.400 ;
        RECT 102.080 49.230 102.250 49.400 ;
        RECT 102.440 49.230 102.610 49.400 ;
        RECT 103.910 49.180 104.080 49.350 ;
        RECT 104.350 49.180 104.520 49.350 ;
        RECT 104.760 49.180 104.930 49.350 ;
        RECT 105.190 49.180 105.360 49.350 ;
        RECT 105.630 49.180 105.800 49.350 ;
        RECT 106.040 49.180 106.210 49.350 ;
        RECT 107.640 49.230 107.810 49.400 ;
        RECT 108.000 49.230 108.170 49.400 ;
        RECT 108.360 49.230 108.530 49.400 ;
        RECT 109.200 49.230 109.370 49.400 ;
        RECT 109.560 49.230 109.730 49.400 ;
        RECT 109.920 49.230 110.090 49.400 ;
        RECT 110.840 49.230 111.010 49.400 ;
        RECT 111.200 49.230 111.370 49.400 ;
        RECT 111.560 49.230 111.730 49.400 ;
        RECT 112.820 49.180 112.990 49.350 ;
        RECT 113.180 49.180 113.350 49.350 ;
        RECT 113.620 49.180 113.790 49.350 ;
        RECT 114.360 49.230 114.530 49.400 ;
        RECT 114.720 49.230 114.890 49.400 ;
        RECT 115.080 49.230 115.250 49.400 ;
        RECT 115.920 49.230 116.090 49.400 ;
        RECT 116.280 49.230 116.450 49.400 ;
        RECT 116.640 49.230 116.810 49.400 ;
        RECT 117.560 49.230 117.730 49.400 ;
        RECT 117.920 49.230 118.090 49.400 ;
        RECT 118.280 49.230 118.450 49.400 ;
        RECT 119.750 49.180 119.920 49.350 ;
        RECT 120.190 49.180 120.360 49.350 ;
        RECT 120.600 49.180 120.770 49.350 ;
        RECT 121.030 49.180 121.200 49.350 ;
        RECT 121.470 49.180 121.640 49.350 ;
        RECT 121.880 49.180 122.050 49.350 ;
        RECT 123.460 49.230 123.630 49.400 ;
        RECT 123.820 49.230 123.990 49.400 ;
        RECT 124.180 49.230 124.350 49.400 ;
        RECT 124.880 49.230 125.050 49.400 ;
        RECT 125.240 49.230 125.410 49.400 ;
        RECT 125.600 49.230 125.770 49.400 ;
        RECT 125.960 49.230 126.130 49.400 ;
        RECT 126.320 49.230 126.490 49.400 ;
        RECT 126.680 49.230 126.850 49.400 ;
        RECT 127.040 49.230 127.210 49.400 ;
        RECT 127.860 49.230 128.030 49.400 ;
        RECT 128.220 49.230 128.390 49.400 ;
        RECT 129.140 49.180 129.310 49.350 ;
        RECT 129.500 49.180 129.670 49.350 ;
        RECT 129.940 49.180 130.110 49.350 ;
        RECT 130.680 49.230 130.850 49.400 ;
        RECT 131.040 49.230 131.210 49.400 ;
        RECT 131.400 49.230 131.570 49.400 ;
        RECT 132.240 49.230 132.410 49.400 ;
        RECT 132.600 49.230 132.770 49.400 ;
        RECT 132.960 49.230 133.130 49.400 ;
        RECT 133.880 49.230 134.050 49.400 ;
        RECT 134.240 49.230 134.410 49.400 ;
        RECT 134.600 49.230 134.770 49.400 ;
        RECT 135.860 49.180 136.030 49.350 ;
        RECT 136.220 49.180 136.390 49.350 ;
        RECT 136.660 49.180 136.830 49.350 ;
        RECT 137.400 49.230 137.570 49.400 ;
        RECT 137.760 49.230 137.930 49.400 ;
        RECT 138.120 49.230 138.290 49.400 ;
        RECT 138.480 49.230 138.650 49.400 ;
        RECT 138.840 49.230 139.010 49.400 ;
        RECT 140.180 49.180 140.350 49.350 ;
        RECT 140.540 49.180 140.710 49.350 ;
        RECT 140.980 49.180 141.150 49.350 ;
        RECT 5.920 48.750 6.090 48.930 ;
        RECT 6.400 48.750 6.570 48.930 ;
        RECT 6.880 48.750 7.050 48.930 ;
        RECT 7.360 48.750 7.530 48.930 ;
        RECT 7.840 48.920 8.010 48.930 ;
      LAYER li1 ;
        RECT 7.680 48.750 8.160 48.920 ;
      LAYER li1 ;
        RECT 8.320 48.750 8.490 48.930 ;
        RECT 8.800 48.750 8.970 48.930 ;
        RECT 9.280 48.750 9.450 48.930 ;
        RECT 9.760 48.750 9.930 48.930 ;
        RECT 10.240 48.750 10.410 48.930 ;
        RECT 10.720 48.750 10.890 48.930 ;
        RECT 11.200 48.750 11.370 48.930 ;
        RECT 11.680 48.750 11.850 48.930 ;
        RECT 12.160 48.750 12.330 48.930 ;
        RECT 12.640 48.750 12.810 48.930 ;
        RECT 13.120 48.750 13.290 48.930 ;
        RECT 13.600 48.750 13.770 48.930 ;
        RECT 14.080 48.750 14.250 48.930 ;
        RECT 14.560 48.750 14.730 48.930 ;
        RECT 15.040 48.750 15.210 48.930 ;
        RECT 15.520 48.750 15.690 48.930 ;
        RECT 16.000 48.750 16.170 48.930 ;
        RECT 16.480 48.750 16.650 48.930 ;
        RECT 16.960 48.750 17.130 48.930 ;
        RECT 17.440 48.750 17.610 48.930 ;
        RECT 17.920 48.750 18.090 48.930 ;
        RECT 18.400 48.750 18.570 48.930 ;
        RECT 18.880 48.750 19.050 48.930 ;
        RECT 19.360 48.750 19.530 48.930 ;
        RECT 19.840 48.750 20.010 48.930 ;
        RECT 20.320 48.750 20.490 48.930 ;
        RECT 20.800 48.750 20.970 48.930 ;
        RECT 21.280 48.750 21.450 48.930 ;
        RECT 21.760 48.750 21.930 48.930 ;
        RECT 22.240 48.750 22.410 48.930 ;
        RECT 22.720 48.750 22.890 48.930 ;
        RECT 23.200 48.750 23.370 48.930 ;
        RECT 23.680 48.750 23.850 48.930 ;
        RECT 24.160 48.750 24.330 48.930 ;
        RECT 24.640 48.750 24.810 48.930 ;
        RECT 25.120 48.750 25.290 48.930 ;
        RECT 25.600 48.750 25.770 48.930 ;
        RECT 26.080 48.750 26.250 48.930 ;
        RECT 26.560 48.750 26.730 48.930 ;
        RECT 27.040 48.750 27.210 48.930 ;
        RECT 27.520 48.750 27.690 48.930 ;
        RECT 28.000 48.750 28.170 48.930 ;
        RECT 28.480 48.750 28.650 48.930 ;
        RECT 28.960 48.750 29.130 48.930 ;
        RECT 29.440 48.750 29.610 48.930 ;
        RECT 29.920 48.750 30.090 48.930 ;
        RECT 30.400 48.750 30.570 48.930 ;
        RECT 30.880 48.750 31.050 48.930 ;
        RECT 31.360 48.750 31.530 48.930 ;
        RECT 31.840 48.750 32.010 48.930 ;
        RECT 32.320 48.750 32.490 48.930 ;
        RECT 32.800 48.750 32.970 48.930 ;
        RECT 33.280 48.750 33.450 48.930 ;
        RECT 33.760 48.750 33.930 48.930 ;
        RECT 34.240 48.750 34.410 48.930 ;
        RECT 34.720 48.750 34.890 48.930 ;
        RECT 35.200 48.750 35.370 48.930 ;
        RECT 35.680 48.750 35.850 48.930 ;
        RECT 36.160 48.750 36.330 48.930 ;
        RECT 36.640 48.750 36.810 48.930 ;
        RECT 37.120 48.750 37.290 48.930 ;
        RECT 37.600 48.750 37.770 48.930 ;
        RECT 38.080 48.750 38.250 48.930 ;
        RECT 38.560 48.750 38.730 48.930 ;
        RECT 39.040 48.750 39.210 48.930 ;
        RECT 39.520 48.750 39.690 48.930 ;
        RECT 40.000 48.750 40.170 48.930 ;
        RECT 40.480 48.750 40.650 48.930 ;
        RECT 40.960 48.750 41.130 48.930 ;
        RECT 41.440 48.750 41.610 48.930 ;
        RECT 41.920 48.750 42.090 48.930 ;
        RECT 42.400 48.750 42.570 48.930 ;
        RECT 42.880 48.750 43.050 48.930 ;
        RECT 43.360 48.750 43.530 48.930 ;
        RECT 43.840 48.750 44.010 48.930 ;
        RECT 44.320 48.750 44.490 48.930 ;
        RECT 44.800 48.750 44.970 48.930 ;
        RECT 45.280 48.750 45.450 48.930 ;
        RECT 45.760 48.750 45.930 48.930 ;
        RECT 46.240 48.750 46.410 48.930 ;
        RECT 46.720 48.750 46.890 48.930 ;
        RECT 47.200 48.750 47.370 48.930 ;
        RECT 47.680 48.920 47.850 48.930 ;
      LAYER li1 ;
        RECT 47.520 48.750 48.000 48.920 ;
      LAYER li1 ;
        RECT 48.160 48.750 48.330 48.930 ;
        RECT 48.640 48.750 48.810 48.930 ;
        RECT 49.120 48.750 49.290 48.930 ;
        RECT 49.600 48.750 49.770 48.930 ;
        RECT 50.080 48.750 50.250 48.930 ;
      LAYER li1 ;
        RECT 50.400 48.920 50.880 48.930 ;
      LAYER li1 ;
        RECT 50.560 48.750 50.730 48.920 ;
        RECT 51.040 48.750 51.210 48.930 ;
        RECT 51.520 48.750 51.690 48.930 ;
        RECT 52.000 48.750 52.170 48.930 ;
        RECT 52.480 48.750 52.650 48.930 ;
        RECT 52.960 48.750 53.130 48.930 ;
        RECT 53.440 48.750 53.610 48.930 ;
        RECT 53.920 48.750 54.090 48.930 ;
        RECT 54.400 48.750 54.570 48.930 ;
        RECT 54.880 48.750 55.050 48.930 ;
        RECT 55.360 48.750 55.530 48.930 ;
        RECT 55.840 48.750 56.010 48.930 ;
        RECT 56.320 48.750 56.490 48.930 ;
        RECT 56.800 48.750 56.970 48.930 ;
        RECT 57.280 48.750 57.450 48.930 ;
        RECT 57.760 48.750 57.930 48.930 ;
        RECT 58.240 48.750 58.410 48.930 ;
        RECT 58.720 48.750 58.890 48.930 ;
        RECT 59.200 48.750 59.370 48.930 ;
        RECT 59.680 48.750 59.850 48.930 ;
        RECT 60.160 48.750 60.330 48.930 ;
        RECT 60.640 48.750 60.810 48.930 ;
        RECT 61.120 48.750 61.290 48.930 ;
        RECT 61.600 48.750 61.770 48.930 ;
        RECT 62.080 48.750 62.250 48.930 ;
        RECT 62.560 48.750 62.730 48.930 ;
        RECT 63.040 48.750 63.210 48.930 ;
        RECT 63.520 48.750 63.690 48.930 ;
        RECT 64.000 48.750 64.170 48.930 ;
        RECT 64.480 48.750 64.650 48.930 ;
        RECT 64.960 48.750 65.130 48.930 ;
        RECT 65.440 48.750 65.610 48.930 ;
        RECT 65.920 48.750 66.090 48.930 ;
        RECT 66.400 48.750 66.570 48.930 ;
        RECT 66.880 48.750 67.050 48.930 ;
        RECT 67.360 48.750 67.530 48.930 ;
        RECT 67.840 48.750 68.010 48.930 ;
        RECT 68.320 48.750 68.490 48.930 ;
        RECT 68.800 48.750 68.970 48.930 ;
        RECT 69.280 48.750 69.450 48.930 ;
        RECT 69.760 48.750 69.930 48.930 ;
        RECT 70.240 48.750 70.410 48.930 ;
        RECT 70.720 48.750 70.890 48.930 ;
        RECT 71.200 48.750 71.370 48.930 ;
        RECT 71.680 48.750 71.850 48.930 ;
        RECT 72.160 48.750 72.330 48.930 ;
        RECT 72.640 48.750 72.810 48.930 ;
        RECT 73.120 48.750 73.290 48.930 ;
        RECT 73.600 48.750 73.770 48.930 ;
        RECT 74.080 48.750 74.250 48.930 ;
        RECT 74.560 48.750 74.730 48.930 ;
        RECT 75.040 48.750 75.210 48.930 ;
        RECT 75.520 48.750 75.690 48.930 ;
        RECT 76.000 48.750 76.170 48.930 ;
        RECT 76.480 48.750 76.650 48.930 ;
        RECT 76.960 48.750 77.130 48.930 ;
        RECT 77.440 48.750 77.610 48.930 ;
        RECT 77.920 48.750 78.090 48.930 ;
        RECT 78.400 48.750 78.570 48.930 ;
        RECT 78.880 48.750 79.050 48.930 ;
        RECT 79.360 48.750 79.530 48.930 ;
        RECT 79.840 48.750 80.010 48.930 ;
        RECT 80.320 48.750 80.490 48.930 ;
        RECT 80.800 48.750 80.970 48.930 ;
        RECT 81.280 48.920 81.450 48.930 ;
      LAYER li1 ;
        RECT 81.120 48.750 81.600 48.920 ;
      LAYER li1 ;
        RECT 81.760 48.750 81.930 48.930 ;
        RECT 82.240 48.750 82.410 48.930 ;
        RECT 82.720 48.750 82.890 48.930 ;
        RECT 83.200 48.750 83.370 48.930 ;
        RECT 83.680 48.750 83.850 48.930 ;
        RECT 84.160 48.750 84.330 48.930 ;
        RECT 84.640 48.750 84.810 48.930 ;
        RECT 85.120 48.750 85.290 48.930 ;
        RECT 85.600 48.750 85.770 48.930 ;
        RECT 86.080 48.750 86.250 48.930 ;
        RECT 86.560 48.750 86.730 48.930 ;
        RECT 87.040 48.750 87.210 48.930 ;
        RECT 87.520 48.750 87.690 48.930 ;
        RECT 88.000 48.750 88.170 48.930 ;
        RECT 88.480 48.750 88.650 48.930 ;
        RECT 88.960 48.750 89.130 48.930 ;
        RECT 89.440 48.750 89.610 48.930 ;
        RECT 89.920 48.750 90.090 48.930 ;
        RECT 90.400 48.750 90.570 48.930 ;
        RECT 90.880 48.750 91.050 48.930 ;
        RECT 91.360 48.750 91.530 48.930 ;
        RECT 91.840 48.750 92.010 48.930 ;
        RECT 92.320 48.750 92.490 48.930 ;
        RECT 92.800 48.750 92.970 48.930 ;
        RECT 93.280 48.750 93.450 48.930 ;
        RECT 93.760 48.750 93.930 48.930 ;
        RECT 94.240 48.750 94.410 48.930 ;
      LAYER li1 ;
        RECT 94.560 48.920 95.040 48.930 ;
      LAYER li1 ;
        RECT 94.720 48.750 94.890 48.920 ;
        RECT 95.200 48.750 95.370 48.930 ;
        RECT 95.680 48.750 95.850 48.930 ;
        RECT 96.160 48.750 96.330 48.930 ;
        RECT 96.640 48.750 96.810 48.930 ;
        RECT 97.120 48.750 97.290 48.930 ;
        RECT 97.600 48.750 97.770 48.930 ;
        RECT 98.080 48.750 98.250 48.930 ;
        RECT 98.560 48.750 98.730 48.930 ;
        RECT 99.040 48.750 99.210 48.930 ;
        RECT 99.520 48.750 99.690 48.930 ;
        RECT 100.000 48.750 100.170 48.930 ;
        RECT 100.480 48.750 100.650 48.930 ;
        RECT 100.960 48.750 101.130 48.930 ;
        RECT 101.440 48.750 101.610 48.930 ;
        RECT 101.920 48.750 102.090 48.930 ;
        RECT 102.400 48.750 102.570 48.930 ;
        RECT 102.880 48.750 103.050 48.930 ;
        RECT 103.360 48.750 103.530 48.930 ;
        RECT 103.840 48.750 104.010 48.930 ;
        RECT 104.320 48.750 104.490 48.930 ;
        RECT 104.800 48.750 104.970 48.930 ;
        RECT 105.280 48.750 105.450 48.930 ;
        RECT 105.760 48.750 105.930 48.930 ;
        RECT 106.240 48.750 106.410 48.930 ;
        RECT 106.720 48.750 106.890 48.930 ;
        RECT 107.200 48.920 107.370 48.930 ;
      LAYER li1 ;
        RECT 107.040 48.750 107.520 48.920 ;
      LAYER li1 ;
        RECT 107.680 48.750 107.850 48.930 ;
      LAYER li1 ;
        RECT 108.000 48.920 108.480 48.930 ;
      LAYER li1 ;
        RECT 108.160 48.750 108.330 48.920 ;
        RECT 108.640 48.750 108.810 48.930 ;
        RECT 109.120 48.750 109.290 48.930 ;
        RECT 109.600 48.750 109.770 48.930 ;
        RECT 110.080 48.750 110.250 48.930 ;
        RECT 110.560 48.750 110.730 48.930 ;
        RECT 111.040 48.750 111.210 48.930 ;
        RECT 111.520 48.750 111.690 48.930 ;
        RECT 112.000 48.750 112.170 48.930 ;
        RECT 112.480 48.750 112.650 48.930 ;
        RECT 112.960 48.750 113.130 48.930 ;
        RECT 113.440 48.750 113.610 48.930 ;
        RECT 113.920 48.750 114.090 48.930 ;
        RECT 114.400 48.750 114.570 48.930 ;
        RECT 114.880 48.750 115.050 48.930 ;
        RECT 115.360 48.750 115.530 48.930 ;
        RECT 115.840 48.750 116.010 48.930 ;
        RECT 116.320 48.750 116.490 48.930 ;
        RECT 116.800 48.750 116.970 48.930 ;
        RECT 117.280 48.750 117.450 48.930 ;
        RECT 117.760 48.750 117.930 48.930 ;
        RECT 118.240 48.750 118.410 48.930 ;
        RECT 118.720 48.750 118.890 48.930 ;
        RECT 119.200 48.750 119.370 48.930 ;
        RECT 119.680 48.750 119.850 48.930 ;
        RECT 120.160 48.750 120.330 48.930 ;
        RECT 120.640 48.750 120.810 48.930 ;
        RECT 121.120 48.750 121.290 48.930 ;
        RECT 121.600 48.750 121.770 48.930 ;
        RECT 122.080 48.750 122.250 48.930 ;
        RECT 122.560 48.750 122.730 48.930 ;
        RECT 123.040 48.920 123.210 48.930 ;
      LAYER li1 ;
        RECT 122.880 48.750 123.360 48.920 ;
      LAYER li1 ;
        RECT 123.520 48.750 123.690 48.930 ;
        RECT 124.000 48.750 124.170 48.930 ;
        RECT 124.480 48.750 124.650 48.930 ;
        RECT 124.960 48.750 125.130 48.930 ;
        RECT 125.440 48.750 125.610 48.930 ;
        RECT 125.920 48.750 126.090 48.930 ;
        RECT 126.400 48.750 126.570 48.930 ;
        RECT 126.880 48.750 127.050 48.930 ;
        RECT 127.360 48.750 127.530 48.930 ;
        RECT 127.840 48.750 128.010 48.930 ;
        RECT 128.320 48.750 128.490 48.930 ;
        RECT 128.800 48.750 128.970 48.930 ;
        RECT 129.280 48.750 129.450 48.930 ;
        RECT 129.760 48.750 129.930 48.930 ;
        RECT 130.240 48.750 130.410 48.930 ;
        RECT 130.720 48.750 130.890 48.930 ;
        RECT 131.200 48.750 131.370 48.930 ;
        RECT 131.680 48.750 131.850 48.930 ;
        RECT 132.160 48.750 132.330 48.930 ;
        RECT 132.640 48.750 132.810 48.930 ;
        RECT 133.120 48.750 133.290 48.930 ;
        RECT 133.600 48.750 133.770 48.930 ;
        RECT 134.080 48.750 134.250 48.930 ;
        RECT 134.560 48.750 134.730 48.930 ;
        RECT 135.040 48.750 135.210 48.930 ;
        RECT 135.520 48.750 135.690 48.930 ;
        RECT 136.000 48.750 136.170 48.930 ;
        RECT 136.480 48.750 136.650 48.930 ;
        RECT 136.960 48.750 137.130 48.930 ;
        RECT 137.440 48.750 137.610 48.930 ;
        RECT 137.920 48.750 138.090 48.930 ;
        RECT 138.400 48.750 138.570 48.930 ;
        RECT 138.880 48.750 139.050 48.930 ;
        RECT 139.360 48.750 139.530 48.930 ;
        RECT 139.840 48.750 140.010 48.930 ;
        RECT 140.320 48.750 140.490 48.930 ;
        RECT 140.800 48.750 140.970 48.930 ;
        RECT 141.280 48.750 141.450 48.930 ;
        RECT 141.760 48.920 141.930 48.930 ;
      LAYER li1 ;
        RECT 141.600 48.750 142.080 48.920 ;
      LAYER li1 ;
        RECT 6.470 48.330 6.640 48.500 ;
        RECT 6.910 48.330 7.080 48.500 ;
        RECT 7.320 48.330 7.490 48.500 ;
        RECT 7.750 48.330 7.920 48.500 ;
        RECT 8.190 48.330 8.360 48.500 ;
        RECT 8.600 48.330 8.770 48.500 ;
        RECT 10.260 48.280 10.430 48.450 ;
        RECT 10.620 48.280 10.790 48.450 ;
        RECT 12.650 48.280 12.820 48.450 ;
        RECT 15.080 48.280 15.250 48.450 ;
        RECT 15.440 48.280 15.610 48.450 ;
        RECT 15.800 48.280 15.970 48.450 ;
        RECT 17.420 48.280 17.590 48.450 ;
        RECT 17.780 48.280 17.950 48.450 ;
        RECT 18.140 48.280 18.310 48.450 ;
        RECT 20.120 48.280 20.290 48.450 ;
        RECT 20.480 48.280 20.650 48.450 ;
        RECT 20.840 48.280 21.010 48.450 ;
        RECT 21.870 48.280 22.040 48.450 ;
        RECT 22.230 48.280 22.400 48.450 ;
        RECT 22.590 48.280 22.760 48.450 ;
        RECT 23.400 48.280 23.570 48.450 ;
        RECT 23.760 48.280 23.930 48.450 ;
        RECT 24.120 48.280 24.290 48.450 ;
        RECT 25.460 48.330 25.630 48.500 ;
        RECT 25.820 48.330 25.990 48.500 ;
        RECT 26.260 48.330 26.430 48.500 ;
        RECT 27.440 48.280 27.610 48.450 ;
        RECT 27.800 48.280 27.970 48.450 ;
        RECT 28.160 48.280 28.330 48.450 ;
        RECT 28.520 48.280 28.690 48.450 ;
        RECT 28.880 48.280 29.050 48.450 ;
        RECT 29.240 48.280 29.410 48.450 ;
        RECT 29.600 48.280 29.770 48.450 ;
        RECT 29.960 48.280 30.130 48.450 ;
        RECT 30.770 48.280 30.940 48.450 ;
        RECT 31.130 48.280 31.300 48.450 ;
        RECT 31.490 48.280 31.660 48.450 ;
        RECT 31.850 48.280 32.020 48.450 ;
        RECT 32.660 48.330 32.830 48.500 ;
        RECT 33.020 48.330 33.190 48.500 ;
        RECT 33.460 48.330 33.630 48.500 ;
        RECT 34.200 48.280 34.370 48.450 ;
        RECT 34.560 48.280 34.730 48.450 ;
        RECT 34.920 48.280 35.090 48.450 ;
        RECT 35.280 48.280 35.450 48.450 ;
        RECT 35.640 48.280 35.810 48.450 ;
        RECT 37.940 48.330 38.110 48.500 ;
        RECT 38.300 48.330 38.470 48.500 ;
        RECT 38.740 48.330 38.910 48.500 ;
        RECT 39.480 48.280 39.650 48.450 ;
        RECT 39.840 48.280 40.010 48.450 ;
        RECT 40.200 48.280 40.370 48.450 ;
        RECT 41.040 48.280 41.210 48.450 ;
        RECT 41.400 48.280 41.570 48.450 ;
        RECT 41.760 48.280 41.930 48.450 ;
        RECT 42.680 48.280 42.850 48.450 ;
        RECT 43.040 48.280 43.210 48.450 ;
        RECT 43.400 48.280 43.570 48.450 ;
        RECT 44.660 48.330 44.830 48.500 ;
        RECT 45.020 48.330 45.190 48.500 ;
        RECT 45.460 48.330 45.630 48.500 ;
        RECT 46.200 48.280 46.370 48.450 ;
        RECT 46.560 48.280 46.730 48.450 ;
        RECT 46.920 48.280 47.090 48.450 ;
        RECT 47.770 48.280 47.940 48.450 ;
        RECT 48.130 48.280 48.300 48.450 ;
        RECT 48.980 48.330 49.150 48.500 ;
        RECT 49.340 48.330 49.510 48.500 ;
        RECT 49.780 48.330 49.950 48.500 ;
        RECT 51.000 48.280 51.170 48.450 ;
        RECT 51.360 48.280 51.530 48.450 ;
        RECT 51.720 48.280 51.890 48.450 ;
        RECT 52.560 48.280 52.730 48.450 ;
        RECT 52.920 48.280 53.090 48.450 ;
        RECT 53.280 48.280 53.450 48.450 ;
        RECT 54.200 48.280 54.370 48.450 ;
        RECT 54.560 48.280 54.730 48.450 ;
        RECT 54.920 48.280 55.090 48.450 ;
        RECT 56.180 48.330 56.350 48.500 ;
        RECT 56.540 48.330 56.710 48.500 ;
        RECT 56.980 48.330 57.150 48.500 ;
        RECT 57.720 48.280 57.890 48.450 ;
        RECT 58.080 48.280 58.250 48.450 ;
        RECT 58.440 48.280 58.610 48.450 ;
        RECT 59.280 48.280 59.450 48.450 ;
        RECT 59.640 48.280 59.810 48.450 ;
        RECT 60.000 48.280 60.170 48.450 ;
        RECT 60.920 48.280 61.090 48.450 ;
        RECT 61.280 48.280 61.450 48.450 ;
        RECT 61.640 48.280 61.810 48.450 ;
        RECT 62.900 48.330 63.070 48.500 ;
        RECT 63.260 48.330 63.430 48.500 ;
        RECT 63.700 48.330 63.870 48.500 ;
        RECT 64.440 48.280 64.610 48.450 ;
        RECT 64.800 48.280 64.970 48.450 ;
        RECT 65.160 48.280 65.330 48.450 ;
        RECT 65.520 48.280 65.690 48.450 ;
        RECT 65.880 48.280 66.050 48.450 ;
        RECT 67.220 48.330 67.390 48.500 ;
        RECT 67.580 48.330 67.750 48.500 ;
        RECT 68.020 48.330 68.190 48.500 ;
        RECT 69.300 48.280 69.470 48.450 ;
        RECT 69.660 48.280 69.830 48.450 ;
        RECT 71.690 48.280 71.860 48.450 ;
        RECT 74.120 48.280 74.290 48.450 ;
        RECT 74.480 48.280 74.650 48.450 ;
        RECT 74.840 48.280 75.010 48.450 ;
        RECT 76.460 48.280 76.630 48.450 ;
        RECT 76.820 48.280 76.990 48.450 ;
        RECT 77.180 48.280 77.350 48.450 ;
        RECT 79.160 48.280 79.330 48.450 ;
        RECT 79.520 48.280 79.690 48.450 ;
        RECT 79.880 48.280 80.050 48.450 ;
        RECT 80.910 48.280 81.080 48.450 ;
        RECT 81.270 48.280 81.440 48.450 ;
        RECT 81.630 48.280 81.800 48.450 ;
        RECT 82.440 48.280 82.610 48.450 ;
        RECT 82.800 48.280 82.970 48.450 ;
        RECT 83.160 48.280 83.330 48.450 ;
        RECT 84.500 48.330 84.670 48.500 ;
        RECT 84.860 48.330 85.030 48.500 ;
        RECT 85.300 48.330 85.470 48.500 ;
        RECT 86.040 48.280 86.210 48.450 ;
        RECT 86.400 48.280 86.570 48.450 ;
        RECT 86.760 48.280 86.930 48.450 ;
        RECT 87.600 48.280 87.770 48.450 ;
        RECT 87.960 48.280 88.130 48.450 ;
        RECT 88.320 48.280 88.490 48.450 ;
        RECT 89.240 48.280 89.410 48.450 ;
        RECT 89.600 48.280 89.770 48.450 ;
        RECT 89.960 48.280 90.130 48.450 ;
        RECT 91.430 48.330 91.600 48.500 ;
        RECT 91.870 48.330 92.040 48.500 ;
        RECT 92.280 48.330 92.450 48.500 ;
        RECT 92.710 48.330 92.880 48.500 ;
        RECT 93.150 48.330 93.320 48.500 ;
        RECT 93.560 48.330 93.730 48.500 ;
        RECT 95.600 48.280 95.770 48.450 ;
        RECT 95.960 48.280 96.130 48.450 ;
        RECT 96.320 48.280 96.490 48.450 ;
        RECT 96.680 48.280 96.850 48.450 ;
        RECT 97.040 48.280 97.210 48.450 ;
        RECT 97.400 48.280 97.570 48.450 ;
        RECT 97.760 48.280 97.930 48.450 ;
        RECT 98.120 48.280 98.290 48.450 ;
        RECT 98.930 48.280 99.100 48.450 ;
        RECT 99.290 48.280 99.460 48.450 ;
        RECT 99.650 48.280 99.820 48.450 ;
        RECT 100.010 48.280 100.180 48.450 ;
        RECT 100.820 48.330 100.990 48.500 ;
        RECT 101.180 48.330 101.350 48.500 ;
        RECT 101.620 48.330 101.790 48.500 ;
        RECT 102.340 48.280 102.510 48.450 ;
        RECT 102.700 48.280 102.870 48.450 ;
        RECT 103.060 48.280 103.230 48.450 ;
        RECT 103.420 48.280 103.590 48.450 ;
        RECT 104.580 48.280 104.750 48.450 ;
        RECT 104.940 48.280 105.110 48.450 ;
        RECT 105.300 48.280 105.470 48.450 ;
        RECT 105.660 48.280 105.830 48.450 ;
        RECT 106.580 48.330 106.750 48.500 ;
        RECT 106.940 48.330 107.110 48.500 ;
        RECT 107.380 48.330 107.550 48.500 ;
        RECT 108.600 48.280 108.770 48.450 ;
        RECT 108.960 48.280 109.130 48.450 ;
        RECT 109.320 48.280 109.490 48.450 ;
        RECT 110.160 48.280 110.330 48.450 ;
        RECT 110.520 48.280 110.690 48.450 ;
        RECT 110.880 48.280 111.050 48.450 ;
        RECT 111.800 48.280 111.970 48.450 ;
        RECT 112.160 48.280 112.330 48.450 ;
        RECT 112.520 48.280 112.690 48.450 ;
        RECT 113.780 48.330 113.950 48.500 ;
        RECT 114.140 48.330 114.310 48.500 ;
        RECT 114.580 48.330 114.750 48.500 ;
        RECT 116.280 48.280 116.450 48.450 ;
        RECT 116.640 48.280 116.810 48.450 ;
        RECT 117.000 48.280 117.170 48.450 ;
        RECT 117.840 48.280 118.010 48.450 ;
        RECT 118.200 48.280 118.370 48.450 ;
        RECT 118.560 48.280 118.730 48.450 ;
        RECT 119.480 48.280 119.650 48.450 ;
        RECT 119.840 48.280 120.010 48.450 ;
        RECT 120.200 48.280 120.370 48.450 ;
        RECT 121.670 48.330 121.840 48.500 ;
        RECT 122.110 48.330 122.280 48.500 ;
        RECT 122.520 48.330 122.690 48.500 ;
        RECT 122.950 48.330 123.120 48.500 ;
        RECT 123.390 48.330 123.560 48.500 ;
        RECT 123.800 48.330 123.970 48.500 ;
        RECT 125.460 48.280 125.630 48.450 ;
        RECT 125.820 48.280 125.990 48.450 ;
        RECT 127.850 48.280 128.020 48.450 ;
        RECT 130.280 48.280 130.450 48.450 ;
        RECT 130.640 48.280 130.810 48.450 ;
        RECT 131.000 48.280 131.170 48.450 ;
        RECT 132.620 48.280 132.790 48.450 ;
        RECT 132.980 48.280 133.150 48.450 ;
        RECT 133.340 48.280 133.510 48.450 ;
        RECT 135.320 48.280 135.490 48.450 ;
        RECT 135.680 48.280 135.850 48.450 ;
        RECT 136.040 48.280 136.210 48.450 ;
        RECT 137.070 48.280 137.240 48.450 ;
        RECT 137.430 48.280 137.600 48.450 ;
        RECT 137.790 48.280 137.960 48.450 ;
        RECT 138.600 48.280 138.770 48.450 ;
        RECT 138.960 48.280 139.130 48.450 ;
        RECT 139.320 48.280 139.490 48.450 ;
        RECT 140.660 48.330 140.830 48.500 ;
        RECT 141.020 48.330 141.190 48.500 ;
        RECT 141.460 48.330 141.630 48.500 ;
        RECT 6.470 41.040 6.640 41.210 ;
        RECT 6.910 41.040 7.080 41.210 ;
        RECT 7.320 41.040 7.490 41.210 ;
        RECT 7.750 41.040 7.920 41.210 ;
        RECT 8.190 41.040 8.360 41.210 ;
        RECT 8.600 41.040 8.770 41.210 ;
        RECT 10.100 41.040 10.270 41.210 ;
        RECT 10.460 41.040 10.630 41.210 ;
        RECT 10.900 41.040 11.070 41.210 ;
        RECT 12.600 41.090 12.770 41.260 ;
        RECT 12.960 41.090 13.130 41.260 ;
        RECT 14.420 41.040 14.590 41.210 ;
        RECT 14.780 41.040 14.950 41.210 ;
        RECT 15.220 41.040 15.390 41.210 ;
        RECT 16.580 41.090 16.750 41.260 ;
        RECT 16.940 41.090 17.110 41.260 ;
        RECT 18.740 41.040 18.910 41.210 ;
        RECT 19.100 41.040 19.270 41.210 ;
        RECT 19.540 41.040 19.710 41.210 ;
        RECT 20.280 41.090 20.450 41.260 ;
        RECT 20.640 41.090 20.810 41.260 ;
        RECT 21.000 41.090 21.170 41.260 ;
        RECT 22.410 41.090 22.580 41.260 ;
        RECT 22.770 41.090 22.940 41.260 ;
        RECT 23.130 41.090 23.300 41.260 ;
        RECT 24.020 41.040 24.190 41.210 ;
        RECT 24.380 41.040 24.550 41.210 ;
        RECT 24.820 41.040 24.990 41.210 ;
        RECT 25.560 41.090 25.730 41.260 ;
        RECT 25.920 41.090 26.090 41.260 ;
        RECT 26.280 41.090 26.450 41.260 ;
        RECT 27.690 41.090 27.860 41.260 ;
        RECT 28.050 41.090 28.220 41.260 ;
        RECT 28.410 41.090 28.580 41.260 ;
        RECT 29.300 41.040 29.470 41.210 ;
        RECT 29.660 41.040 29.830 41.210 ;
        RECT 30.100 41.040 30.270 41.210 ;
        RECT 30.840 41.090 31.010 41.260 ;
        RECT 31.200 41.090 31.370 41.260 ;
        RECT 31.560 41.090 31.730 41.260 ;
        RECT 32.400 41.090 32.570 41.260 ;
        RECT 32.760 41.090 32.930 41.260 ;
        RECT 33.120 41.090 33.290 41.260 ;
        RECT 34.040 41.090 34.210 41.260 ;
        RECT 34.400 41.090 34.570 41.260 ;
        RECT 34.760 41.090 34.930 41.260 ;
        RECT 36.020 41.040 36.190 41.210 ;
        RECT 36.380 41.040 36.550 41.210 ;
        RECT 36.820 41.040 36.990 41.210 ;
        RECT 37.560 41.090 37.730 41.260 ;
        RECT 37.920 41.090 38.090 41.260 ;
        RECT 39.380 41.040 39.550 41.210 ;
        RECT 39.740 41.040 39.910 41.210 ;
        RECT 40.180 41.040 40.350 41.210 ;
        RECT 40.920 41.090 41.090 41.260 ;
        RECT 41.280 41.090 41.450 41.260 ;
        RECT 41.640 41.090 41.810 41.260 ;
        RECT 42.480 41.090 42.650 41.260 ;
        RECT 42.840 41.090 43.010 41.260 ;
        RECT 43.200 41.090 43.370 41.260 ;
        RECT 44.120 41.090 44.290 41.260 ;
        RECT 44.480 41.090 44.650 41.260 ;
        RECT 44.840 41.090 45.010 41.260 ;
        RECT 46.100 41.040 46.270 41.210 ;
        RECT 46.460 41.040 46.630 41.210 ;
        RECT 46.900 41.040 47.070 41.210 ;
        RECT 47.640 41.090 47.810 41.260 ;
        RECT 48.000 41.090 48.170 41.260 ;
        RECT 48.360 41.090 48.530 41.260 ;
        RECT 49.200 41.090 49.370 41.260 ;
        RECT 49.560 41.090 49.730 41.260 ;
        RECT 49.920 41.090 50.090 41.260 ;
        RECT 50.840 41.090 51.010 41.260 ;
        RECT 51.200 41.090 51.370 41.260 ;
        RECT 51.560 41.090 51.730 41.260 ;
        RECT 52.820 41.040 52.990 41.210 ;
        RECT 53.180 41.040 53.350 41.210 ;
        RECT 53.620 41.040 53.790 41.210 ;
        RECT 54.360 41.090 54.530 41.260 ;
        RECT 54.720 41.090 54.890 41.260 ;
        RECT 55.080 41.090 55.250 41.260 ;
        RECT 55.920 41.090 56.090 41.260 ;
        RECT 56.280 41.090 56.450 41.260 ;
        RECT 56.640 41.090 56.810 41.260 ;
        RECT 57.560 41.090 57.730 41.260 ;
        RECT 57.920 41.090 58.090 41.260 ;
        RECT 58.280 41.090 58.450 41.260 ;
        RECT 59.540 41.040 59.710 41.210 ;
        RECT 59.900 41.040 60.070 41.210 ;
        RECT 60.340 41.040 60.510 41.210 ;
        RECT 61.080 41.090 61.250 41.260 ;
        RECT 61.440 41.090 61.610 41.260 ;
        RECT 61.800 41.090 61.970 41.260 ;
        RECT 62.640 41.090 62.810 41.260 ;
        RECT 63.000 41.090 63.170 41.260 ;
        RECT 63.360 41.090 63.530 41.260 ;
        RECT 64.280 41.090 64.450 41.260 ;
        RECT 64.640 41.090 64.810 41.260 ;
        RECT 65.000 41.090 65.170 41.260 ;
        RECT 66.260 41.040 66.430 41.210 ;
        RECT 66.620 41.040 66.790 41.210 ;
        RECT 67.060 41.040 67.230 41.210 ;
        RECT 67.800 41.090 67.970 41.260 ;
        RECT 68.160 41.090 68.330 41.260 ;
        RECT 68.520 41.090 68.690 41.260 ;
        RECT 69.360 41.090 69.530 41.260 ;
        RECT 69.720 41.090 69.890 41.260 ;
        RECT 70.080 41.090 70.250 41.260 ;
        RECT 71.000 41.090 71.170 41.260 ;
        RECT 71.360 41.090 71.530 41.260 ;
        RECT 71.720 41.090 71.890 41.260 ;
        RECT 72.980 41.040 73.150 41.210 ;
        RECT 73.340 41.040 73.510 41.210 ;
        RECT 73.780 41.040 73.950 41.210 ;
        RECT 74.520 41.090 74.690 41.260 ;
        RECT 74.880 41.090 75.050 41.260 ;
        RECT 75.240 41.090 75.410 41.260 ;
        RECT 76.080 41.090 76.250 41.260 ;
        RECT 76.440 41.090 76.610 41.260 ;
        RECT 76.800 41.090 76.970 41.260 ;
        RECT 77.720 41.090 77.890 41.260 ;
        RECT 78.080 41.090 78.250 41.260 ;
        RECT 78.440 41.090 78.610 41.260 ;
        RECT 79.700 41.040 79.870 41.210 ;
        RECT 80.060 41.040 80.230 41.210 ;
        RECT 80.500 41.040 80.670 41.210 ;
        RECT 81.240 41.090 81.410 41.260 ;
        RECT 81.600 41.090 81.770 41.260 ;
        RECT 81.960 41.090 82.130 41.260 ;
        RECT 82.800 41.090 82.970 41.260 ;
        RECT 83.160 41.090 83.330 41.260 ;
        RECT 83.520 41.090 83.690 41.260 ;
        RECT 84.440 41.090 84.610 41.260 ;
        RECT 84.800 41.090 84.970 41.260 ;
        RECT 85.160 41.090 85.330 41.260 ;
        RECT 86.420 41.040 86.590 41.210 ;
        RECT 86.780 41.040 86.950 41.210 ;
        RECT 87.220 41.040 87.390 41.210 ;
        RECT 87.960 41.090 88.130 41.260 ;
        RECT 88.320 41.090 88.490 41.260 ;
        RECT 88.680 41.090 88.850 41.260 ;
        RECT 89.520 41.090 89.690 41.260 ;
        RECT 89.880 41.090 90.050 41.260 ;
        RECT 90.240 41.090 90.410 41.260 ;
        RECT 91.160 41.090 91.330 41.260 ;
        RECT 91.520 41.090 91.690 41.260 ;
        RECT 91.880 41.090 92.050 41.260 ;
        RECT 93.140 41.040 93.310 41.210 ;
        RECT 93.500 41.040 93.670 41.210 ;
        RECT 93.940 41.040 94.110 41.210 ;
        RECT 94.660 41.090 94.830 41.260 ;
        RECT 95.020 41.090 95.190 41.260 ;
        RECT 95.380 41.090 95.550 41.260 ;
        RECT 95.740 41.090 95.910 41.260 ;
        RECT 96.900 41.090 97.070 41.260 ;
        RECT 97.260 41.090 97.430 41.260 ;
        RECT 97.620 41.090 97.790 41.260 ;
        RECT 97.980 41.090 98.150 41.260 ;
        RECT 98.900 41.040 99.070 41.210 ;
        RECT 99.260 41.040 99.430 41.210 ;
        RECT 99.700 41.040 99.870 41.210 ;
        RECT 101.400 41.090 101.570 41.260 ;
        RECT 101.760 41.090 101.930 41.260 ;
        RECT 102.120 41.090 102.290 41.260 ;
        RECT 102.960 41.090 103.130 41.260 ;
        RECT 103.320 41.090 103.490 41.260 ;
        RECT 103.680 41.090 103.850 41.260 ;
        RECT 104.600 41.090 104.770 41.260 ;
        RECT 104.960 41.090 105.130 41.260 ;
        RECT 105.320 41.090 105.490 41.260 ;
        RECT 106.580 41.040 106.750 41.210 ;
        RECT 106.940 41.040 107.110 41.210 ;
        RECT 107.380 41.040 107.550 41.210 ;
        RECT 108.120 41.090 108.290 41.260 ;
        RECT 108.480 41.090 108.650 41.260 ;
        RECT 108.840 41.090 109.010 41.260 ;
        RECT 109.680 41.090 109.850 41.260 ;
        RECT 110.040 41.090 110.210 41.260 ;
        RECT 110.400 41.090 110.570 41.260 ;
        RECT 111.320 41.090 111.490 41.260 ;
        RECT 111.680 41.090 111.850 41.260 ;
        RECT 112.040 41.090 112.210 41.260 ;
        RECT 113.300 41.040 113.470 41.210 ;
        RECT 113.660 41.040 113.830 41.210 ;
        RECT 114.100 41.040 114.270 41.210 ;
        RECT 116.280 41.090 116.450 41.260 ;
        RECT 116.640 41.090 116.810 41.260 ;
        RECT 117.000 41.090 117.170 41.260 ;
        RECT 117.840 41.090 118.010 41.260 ;
        RECT 118.200 41.090 118.370 41.260 ;
        RECT 118.560 41.090 118.730 41.260 ;
        RECT 119.480 41.090 119.650 41.260 ;
        RECT 119.840 41.090 120.010 41.260 ;
        RECT 120.200 41.090 120.370 41.260 ;
        RECT 121.460 41.040 121.630 41.210 ;
        RECT 121.820 41.040 121.990 41.210 ;
        RECT 122.260 41.040 122.430 41.210 ;
        RECT 123.000 41.090 123.170 41.260 ;
        RECT 123.360 41.090 123.530 41.260 ;
        RECT 123.720 41.090 123.890 41.260 ;
        RECT 124.560 41.090 124.730 41.260 ;
        RECT 124.920 41.090 125.090 41.260 ;
        RECT 125.280 41.090 125.450 41.260 ;
        RECT 126.200 41.090 126.370 41.260 ;
        RECT 126.560 41.090 126.730 41.260 ;
        RECT 126.920 41.090 127.090 41.260 ;
        RECT 128.180 41.040 128.350 41.210 ;
        RECT 128.540 41.040 128.710 41.210 ;
        RECT 128.980 41.040 129.150 41.210 ;
        RECT 129.720 41.090 129.890 41.260 ;
        RECT 130.080 41.090 130.250 41.260 ;
        RECT 130.440 41.090 130.610 41.260 ;
        RECT 131.280 41.090 131.450 41.260 ;
        RECT 131.640 41.090 131.810 41.260 ;
        RECT 132.000 41.090 132.170 41.260 ;
        RECT 132.920 41.090 133.090 41.260 ;
        RECT 133.280 41.090 133.450 41.260 ;
        RECT 133.640 41.090 133.810 41.260 ;
        RECT 134.900 41.040 135.070 41.210 ;
        RECT 135.260 41.040 135.430 41.210 ;
        RECT 135.700 41.040 135.870 41.210 ;
        RECT 137.010 41.090 137.180 41.260 ;
        RECT 137.370 41.090 137.540 41.260 ;
        RECT 137.730 41.090 137.900 41.260 ;
        RECT 138.090 41.090 138.260 41.260 ;
        RECT 140.180 41.040 140.350 41.210 ;
        RECT 140.540 41.040 140.710 41.210 ;
        RECT 140.980 41.040 141.150 41.210 ;
        RECT 5.920 40.610 6.090 40.790 ;
        RECT 6.400 40.610 6.570 40.790 ;
        RECT 6.880 40.610 7.050 40.790 ;
        RECT 7.360 40.610 7.530 40.790 ;
        RECT 7.840 40.610 8.010 40.790 ;
        RECT 8.320 40.610 8.490 40.790 ;
        RECT 8.800 40.610 8.970 40.790 ;
        RECT 9.280 40.610 9.450 40.790 ;
        RECT 9.760 40.610 9.930 40.790 ;
        RECT 10.240 40.610 10.410 40.790 ;
        RECT 10.720 40.610 10.890 40.790 ;
        RECT 11.200 40.610 11.370 40.790 ;
        RECT 11.680 40.610 11.850 40.790 ;
        RECT 12.160 40.610 12.330 40.790 ;
        RECT 12.640 40.610 12.810 40.790 ;
        RECT 13.120 40.610 13.290 40.790 ;
        RECT 13.600 40.610 13.770 40.790 ;
        RECT 14.080 40.610 14.250 40.790 ;
      LAYER li1 ;
        RECT 14.400 40.780 14.880 40.790 ;
      LAYER li1 ;
        RECT 14.560 40.610 14.730 40.780 ;
        RECT 15.040 40.610 15.210 40.790 ;
        RECT 15.520 40.610 15.690 40.790 ;
        RECT 16.000 40.610 16.170 40.790 ;
        RECT 16.480 40.610 16.650 40.790 ;
        RECT 16.960 40.610 17.130 40.790 ;
        RECT 17.440 40.610 17.610 40.790 ;
        RECT 17.920 40.610 18.090 40.790 ;
        RECT 18.400 40.610 18.570 40.790 ;
        RECT 18.880 40.610 19.050 40.790 ;
        RECT 19.360 40.610 19.530 40.790 ;
        RECT 19.840 40.610 20.010 40.790 ;
        RECT 20.320 40.610 20.490 40.790 ;
        RECT 20.800 40.610 20.970 40.790 ;
        RECT 21.280 40.610 21.450 40.790 ;
        RECT 21.760 40.610 21.930 40.790 ;
        RECT 22.240 40.610 22.410 40.790 ;
        RECT 22.720 40.610 22.890 40.790 ;
        RECT 23.200 40.610 23.370 40.790 ;
        RECT 23.680 40.610 23.850 40.790 ;
        RECT 24.160 40.610 24.330 40.790 ;
        RECT 24.640 40.610 24.810 40.790 ;
        RECT 25.120 40.610 25.290 40.790 ;
        RECT 25.600 40.610 25.770 40.790 ;
        RECT 26.080 40.610 26.250 40.790 ;
        RECT 26.560 40.610 26.730 40.790 ;
        RECT 27.040 40.610 27.210 40.790 ;
        RECT 27.520 40.610 27.690 40.790 ;
        RECT 28.000 40.610 28.170 40.790 ;
        RECT 28.480 40.610 28.650 40.790 ;
        RECT 28.960 40.610 29.130 40.790 ;
        RECT 29.440 40.610 29.610 40.790 ;
        RECT 29.920 40.610 30.090 40.790 ;
        RECT 30.400 40.610 30.570 40.790 ;
        RECT 30.880 40.610 31.050 40.790 ;
        RECT 31.360 40.610 31.530 40.790 ;
        RECT 31.840 40.610 32.010 40.790 ;
        RECT 32.320 40.610 32.490 40.790 ;
        RECT 32.800 40.610 32.970 40.790 ;
        RECT 33.280 40.610 33.450 40.790 ;
        RECT 33.760 40.610 33.930 40.790 ;
        RECT 34.240 40.610 34.410 40.790 ;
        RECT 34.720 40.610 34.890 40.790 ;
        RECT 35.200 40.610 35.370 40.790 ;
        RECT 35.680 40.610 35.850 40.790 ;
        RECT 36.160 40.610 36.330 40.790 ;
        RECT 36.640 40.610 36.810 40.790 ;
        RECT 37.120 40.610 37.290 40.790 ;
        RECT 37.600 40.610 37.770 40.790 ;
        RECT 38.080 40.610 38.250 40.790 ;
        RECT 38.560 40.610 38.730 40.790 ;
        RECT 39.040 40.610 39.210 40.790 ;
        RECT 39.520 40.610 39.690 40.790 ;
        RECT 40.000 40.610 40.170 40.790 ;
        RECT 40.480 40.610 40.650 40.790 ;
        RECT 40.960 40.610 41.130 40.790 ;
        RECT 41.440 40.610 41.610 40.790 ;
        RECT 41.920 40.610 42.090 40.790 ;
        RECT 42.400 40.610 42.570 40.790 ;
        RECT 42.880 40.610 43.050 40.790 ;
        RECT 43.360 40.610 43.530 40.790 ;
        RECT 43.840 40.610 44.010 40.790 ;
        RECT 44.320 40.610 44.490 40.790 ;
        RECT 44.800 40.610 44.970 40.790 ;
        RECT 45.280 40.610 45.450 40.790 ;
        RECT 45.760 40.610 45.930 40.790 ;
        RECT 46.240 40.610 46.410 40.790 ;
        RECT 46.720 40.610 46.890 40.790 ;
        RECT 47.200 40.610 47.370 40.790 ;
        RECT 47.680 40.610 47.850 40.790 ;
        RECT 48.160 40.610 48.330 40.790 ;
        RECT 48.640 40.610 48.810 40.790 ;
        RECT 49.120 40.610 49.290 40.790 ;
        RECT 49.600 40.610 49.770 40.790 ;
        RECT 50.080 40.610 50.250 40.790 ;
        RECT 50.560 40.610 50.730 40.790 ;
        RECT 51.040 40.610 51.210 40.790 ;
        RECT 51.520 40.610 51.690 40.790 ;
        RECT 52.000 40.610 52.170 40.790 ;
        RECT 52.480 40.610 52.650 40.790 ;
        RECT 52.960 40.610 53.130 40.790 ;
        RECT 53.440 40.610 53.610 40.790 ;
        RECT 53.920 40.610 54.090 40.790 ;
        RECT 54.400 40.610 54.570 40.790 ;
        RECT 54.880 40.610 55.050 40.790 ;
        RECT 55.360 40.610 55.530 40.790 ;
        RECT 55.840 40.610 56.010 40.790 ;
        RECT 56.320 40.610 56.490 40.790 ;
        RECT 56.800 40.610 56.970 40.790 ;
        RECT 57.280 40.610 57.450 40.790 ;
        RECT 57.760 40.610 57.930 40.790 ;
        RECT 58.240 40.610 58.410 40.790 ;
        RECT 58.720 40.610 58.890 40.790 ;
        RECT 59.200 40.610 59.370 40.790 ;
        RECT 59.680 40.610 59.850 40.790 ;
        RECT 60.160 40.610 60.330 40.790 ;
        RECT 60.640 40.610 60.810 40.790 ;
        RECT 61.120 40.610 61.290 40.790 ;
        RECT 61.600 40.610 61.770 40.790 ;
        RECT 62.080 40.610 62.250 40.790 ;
        RECT 62.560 40.610 62.730 40.790 ;
        RECT 63.040 40.610 63.210 40.790 ;
        RECT 63.520 40.610 63.690 40.790 ;
        RECT 64.000 40.610 64.170 40.790 ;
        RECT 64.480 40.610 64.650 40.790 ;
        RECT 64.960 40.610 65.130 40.790 ;
        RECT 65.440 40.610 65.610 40.790 ;
        RECT 65.920 40.610 66.090 40.790 ;
        RECT 66.400 40.610 66.570 40.790 ;
        RECT 66.880 40.610 67.050 40.790 ;
        RECT 67.360 40.610 67.530 40.790 ;
        RECT 67.840 40.610 68.010 40.790 ;
        RECT 68.320 40.610 68.490 40.790 ;
        RECT 68.800 40.610 68.970 40.790 ;
        RECT 69.280 40.610 69.450 40.790 ;
        RECT 69.760 40.610 69.930 40.790 ;
        RECT 70.240 40.610 70.410 40.790 ;
        RECT 70.720 40.610 70.890 40.790 ;
        RECT 71.200 40.610 71.370 40.790 ;
        RECT 71.680 40.610 71.850 40.790 ;
        RECT 72.160 40.610 72.330 40.790 ;
        RECT 72.640 40.610 72.810 40.790 ;
        RECT 73.120 40.610 73.290 40.790 ;
        RECT 73.600 40.610 73.770 40.790 ;
        RECT 74.080 40.610 74.250 40.790 ;
        RECT 74.560 40.610 74.730 40.790 ;
        RECT 75.040 40.610 75.210 40.790 ;
        RECT 75.520 40.610 75.690 40.790 ;
        RECT 76.000 40.610 76.170 40.790 ;
        RECT 76.480 40.610 76.650 40.790 ;
        RECT 76.960 40.610 77.130 40.790 ;
        RECT 77.440 40.610 77.610 40.790 ;
      LAYER li1 ;
        RECT 77.760 40.780 78.240 40.790 ;
      LAYER li1 ;
        RECT 77.920 40.610 78.090 40.780 ;
        RECT 78.400 40.610 78.570 40.790 ;
        RECT 78.880 40.610 79.050 40.790 ;
        RECT 79.360 40.610 79.530 40.790 ;
        RECT 79.840 40.610 80.010 40.790 ;
        RECT 80.320 40.610 80.490 40.790 ;
        RECT 80.800 40.610 80.970 40.790 ;
        RECT 81.280 40.610 81.450 40.790 ;
        RECT 81.760 40.610 81.930 40.790 ;
        RECT 82.240 40.610 82.410 40.790 ;
        RECT 82.720 40.610 82.890 40.790 ;
        RECT 83.200 40.610 83.370 40.790 ;
        RECT 83.680 40.610 83.850 40.790 ;
        RECT 84.160 40.610 84.330 40.790 ;
        RECT 84.640 40.610 84.810 40.790 ;
        RECT 85.120 40.610 85.290 40.790 ;
        RECT 85.600 40.610 85.770 40.790 ;
        RECT 86.080 40.610 86.250 40.790 ;
        RECT 86.560 40.610 86.730 40.790 ;
        RECT 87.040 40.610 87.210 40.790 ;
        RECT 87.520 40.610 87.690 40.790 ;
        RECT 88.000 40.610 88.170 40.790 ;
        RECT 88.480 40.610 88.650 40.790 ;
        RECT 88.960 40.610 89.130 40.790 ;
        RECT 89.440 40.610 89.610 40.790 ;
        RECT 89.920 40.610 90.090 40.790 ;
        RECT 90.400 40.610 90.570 40.790 ;
        RECT 90.880 40.610 91.050 40.790 ;
        RECT 91.360 40.610 91.530 40.790 ;
        RECT 91.840 40.610 92.010 40.790 ;
        RECT 92.320 40.610 92.490 40.790 ;
        RECT 92.800 40.610 92.970 40.790 ;
        RECT 93.280 40.610 93.450 40.790 ;
        RECT 93.760 40.610 93.930 40.790 ;
        RECT 94.240 40.610 94.410 40.790 ;
        RECT 94.720 40.610 94.890 40.790 ;
        RECT 95.200 40.610 95.370 40.790 ;
        RECT 95.680 40.610 95.850 40.790 ;
        RECT 96.160 40.610 96.330 40.790 ;
        RECT 96.640 40.610 96.810 40.790 ;
        RECT 97.120 40.610 97.290 40.790 ;
        RECT 97.600 40.610 97.770 40.790 ;
        RECT 98.080 40.610 98.250 40.790 ;
        RECT 98.560 40.610 98.730 40.790 ;
        RECT 99.040 40.610 99.210 40.790 ;
        RECT 99.520 40.610 99.690 40.790 ;
        RECT 100.000 40.610 100.170 40.790 ;
        RECT 100.480 40.610 100.650 40.790 ;
        RECT 100.960 40.610 101.130 40.790 ;
        RECT 101.440 40.610 101.610 40.790 ;
        RECT 101.920 40.610 102.090 40.790 ;
        RECT 102.400 40.610 102.570 40.790 ;
        RECT 102.880 40.610 103.050 40.790 ;
        RECT 103.360 40.610 103.530 40.790 ;
        RECT 103.840 40.610 104.010 40.790 ;
        RECT 104.320 40.610 104.490 40.790 ;
        RECT 104.800 40.610 104.970 40.790 ;
        RECT 105.280 40.610 105.450 40.790 ;
        RECT 105.760 40.610 105.930 40.790 ;
        RECT 106.240 40.610 106.410 40.790 ;
        RECT 106.720 40.610 106.890 40.790 ;
        RECT 107.200 40.610 107.370 40.790 ;
        RECT 107.680 40.610 107.850 40.790 ;
        RECT 108.160 40.610 108.330 40.790 ;
        RECT 108.640 40.610 108.810 40.790 ;
        RECT 109.120 40.610 109.290 40.790 ;
        RECT 109.600 40.610 109.770 40.790 ;
        RECT 110.080 40.610 110.250 40.790 ;
      LAYER li1 ;
        RECT 110.400 40.780 110.880 40.790 ;
      LAYER li1 ;
        RECT 110.560 40.610 110.730 40.780 ;
        RECT 111.040 40.610 111.210 40.790 ;
        RECT 111.520 40.610 111.690 40.790 ;
        RECT 112.000 40.610 112.170 40.790 ;
        RECT 112.480 40.610 112.650 40.790 ;
        RECT 112.960 40.610 113.130 40.790 ;
        RECT 113.440 40.610 113.610 40.790 ;
        RECT 113.920 40.610 114.090 40.790 ;
        RECT 114.400 40.610 114.570 40.790 ;
        RECT 114.880 40.610 115.050 40.790 ;
        RECT 115.360 40.610 115.530 40.790 ;
        RECT 115.840 40.780 116.010 40.790 ;
      LAYER li1 ;
        RECT 115.680 40.610 116.160 40.780 ;
      LAYER li1 ;
        RECT 116.320 40.610 116.490 40.790 ;
        RECT 116.800 40.610 116.970 40.790 ;
        RECT 117.280 40.610 117.450 40.790 ;
        RECT 117.760 40.610 117.930 40.790 ;
        RECT 118.240 40.610 118.410 40.790 ;
        RECT 118.720 40.610 118.890 40.790 ;
        RECT 119.200 40.610 119.370 40.790 ;
        RECT 119.680 40.610 119.850 40.790 ;
        RECT 120.160 40.610 120.330 40.790 ;
        RECT 120.640 40.610 120.810 40.790 ;
        RECT 121.120 40.610 121.290 40.790 ;
        RECT 121.600 40.610 121.770 40.790 ;
        RECT 122.080 40.610 122.250 40.790 ;
        RECT 122.560 40.610 122.730 40.790 ;
        RECT 123.040 40.610 123.210 40.790 ;
        RECT 123.520 40.610 123.690 40.790 ;
        RECT 124.000 40.610 124.170 40.790 ;
        RECT 124.480 40.610 124.650 40.790 ;
        RECT 124.960 40.610 125.130 40.790 ;
        RECT 125.440 40.610 125.610 40.790 ;
        RECT 125.920 40.610 126.090 40.790 ;
        RECT 126.400 40.610 126.570 40.790 ;
        RECT 126.880 40.610 127.050 40.790 ;
        RECT 127.360 40.610 127.530 40.790 ;
        RECT 127.840 40.610 128.010 40.790 ;
        RECT 128.320 40.610 128.490 40.790 ;
        RECT 128.800 40.610 128.970 40.790 ;
        RECT 129.280 40.610 129.450 40.790 ;
        RECT 129.760 40.610 129.930 40.790 ;
        RECT 130.240 40.610 130.410 40.790 ;
        RECT 130.720 40.610 130.890 40.790 ;
        RECT 131.200 40.610 131.370 40.790 ;
        RECT 131.680 40.610 131.850 40.790 ;
        RECT 132.160 40.610 132.330 40.790 ;
        RECT 132.640 40.610 132.810 40.790 ;
        RECT 133.120 40.610 133.290 40.790 ;
        RECT 133.600 40.610 133.770 40.790 ;
        RECT 134.080 40.610 134.250 40.790 ;
        RECT 134.560 40.610 134.730 40.790 ;
        RECT 135.040 40.610 135.210 40.790 ;
        RECT 135.520 40.610 135.690 40.790 ;
        RECT 136.000 40.610 136.170 40.790 ;
        RECT 136.480 40.610 136.650 40.790 ;
        RECT 136.960 40.610 137.130 40.790 ;
        RECT 137.440 40.610 137.610 40.790 ;
        RECT 137.920 40.610 138.090 40.790 ;
        RECT 138.400 40.610 138.570 40.790 ;
        RECT 138.880 40.610 139.050 40.790 ;
        RECT 139.360 40.610 139.530 40.790 ;
        RECT 139.840 40.610 140.010 40.790 ;
        RECT 140.320 40.610 140.490 40.790 ;
        RECT 140.800 40.610 140.970 40.790 ;
        RECT 141.280 40.610 141.450 40.790 ;
        RECT 141.760 40.780 141.930 40.790 ;
      LAYER li1 ;
        RECT 141.600 40.610 142.080 40.780 ;
      LAYER li1 ;
        RECT 6.470 40.190 6.640 40.360 ;
        RECT 6.910 40.190 7.080 40.360 ;
        RECT 7.320 40.190 7.490 40.360 ;
        RECT 7.750 40.190 7.920 40.360 ;
        RECT 8.190 40.190 8.360 40.360 ;
        RECT 8.600 40.190 8.770 40.360 ;
        RECT 10.310 40.190 10.480 40.360 ;
        RECT 10.750 40.190 10.920 40.360 ;
        RECT 11.160 40.190 11.330 40.360 ;
        RECT 11.590 40.190 11.760 40.360 ;
        RECT 12.030 40.190 12.200 40.360 ;
        RECT 12.440 40.190 12.610 40.360 ;
        RECT 15.000 40.140 15.170 40.310 ;
        RECT 15.360 40.140 15.530 40.310 ;
        RECT 16.820 40.190 16.990 40.360 ;
        RECT 17.180 40.190 17.350 40.360 ;
        RECT 17.620 40.190 17.790 40.360 ;
        RECT 18.360 40.140 18.530 40.310 ;
        RECT 18.720 40.140 18.890 40.310 ;
        RECT 19.080 40.140 19.250 40.310 ;
        RECT 19.440 40.140 19.610 40.310 ;
        RECT 19.800 40.140 19.970 40.310 ;
        RECT 21.140 40.190 21.310 40.360 ;
        RECT 21.500 40.190 21.670 40.360 ;
        RECT 21.940 40.190 22.110 40.360 ;
        RECT 22.680 40.140 22.850 40.310 ;
        RECT 23.040 40.140 23.210 40.310 ;
        RECT 23.400 40.140 23.570 40.310 ;
        RECT 23.760 40.140 23.930 40.310 ;
        RECT 24.120 40.140 24.290 40.310 ;
        RECT 25.460 40.190 25.630 40.360 ;
        RECT 25.820 40.190 25.990 40.360 ;
        RECT 26.260 40.190 26.430 40.360 ;
        RECT 27.000 40.140 27.170 40.310 ;
        RECT 27.360 40.140 27.530 40.310 ;
        RECT 27.720 40.140 27.890 40.310 ;
        RECT 28.080 40.140 28.250 40.310 ;
        RECT 28.440 40.140 28.610 40.310 ;
        RECT 30.740 40.190 30.910 40.360 ;
        RECT 31.100 40.190 31.270 40.360 ;
        RECT 31.540 40.190 31.710 40.360 ;
        RECT 32.280 40.140 32.450 40.310 ;
        RECT 32.640 40.140 32.810 40.310 ;
        RECT 33.000 40.140 33.170 40.310 ;
        RECT 33.360 40.140 33.530 40.310 ;
        RECT 33.720 40.140 33.890 40.310 ;
        RECT 36.020 40.190 36.190 40.360 ;
        RECT 36.380 40.190 36.550 40.360 ;
        RECT 36.820 40.190 36.990 40.360 ;
        RECT 37.560 40.140 37.730 40.310 ;
        RECT 37.920 40.140 38.090 40.310 ;
        RECT 38.280 40.140 38.450 40.310 ;
        RECT 39.120 40.140 39.290 40.310 ;
        RECT 39.480 40.140 39.650 40.310 ;
        RECT 39.840 40.140 40.010 40.310 ;
        RECT 40.760 40.140 40.930 40.310 ;
        RECT 41.120 40.140 41.290 40.310 ;
        RECT 41.480 40.140 41.650 40.310 ;
        RECT 42.740 40.190 42.910 40.360 ;
        RECT 43.100 40.190 43.270 40.360 ;
        RECT 43.540 40.190 43.710 40.360 ;
        RECT 44.280 40.140 44.450 40.310 ;
        RECT 44.640 40.140 44.810 40.310 ;
        RECT 45.000 40.140 45.170 40.310 ;
        RECT 45.840 40.140 46.010 40.310 ;
        RECT 46.200 40.140 46.370 40.310 ;
        RECT 46.560 40.140 46.730 40.310 ;
        RECT 47.480 40.140 47.650 40.310 ;
        RECT 47.840 40.140 48.010 40.310 ;
        RECT 48.200 40.140 48.370 40.310 ;
        RECT 49.460 40.190 49.630 40.360 ;
        RECT 49.820 40.190 49.990 40.360 ;
        RECT 50.260 40.190 50.430 40.360 ;
        RECT 51.000 40.140 51.170 40.310 ;
        RECT 51.360 40.140 51.530 40.310 ;
        RECT 51.720 40.140 51.890 40.310 ;
        RECT 52.560 40.140 52.730 40.310 ;
        RECT 52.920 40.140 53.090 40.310 ;
        RECT 53.280 40.140 53.450 40.310 ;
        RECT 54.200 40.140 54.370 40.310 ;
        RECT 54.560 40.140 54.730 40.310 ;
        RECT 54.920 40.140 55.090 40.310 ;
        RECT 56.180 40.190 56.350 40.360 ;
        RECT 56.540 40.190 56.710 40.360 ;
        RECT 56.980 40.190 57.150 40.360 ;
        RECT 57.720 40.140 57.890 40.310 ;
        RECT 58.080 40.140 58.250 40.310 ;
        RECT 58.440 40.140 58.610 40.310 ;
        RECT 59.280 40.140 59.450 40.310 ;
        RECT 59.640 40.140 59.810 40.310 ;
        RECT 60.000 40.140 60.170 40.310 ;
        RECT 60.920 40.140 61.090 40.310 ;
        RECT 61.280 40.140 61.450 40.310 ;
        RECT 61.640 40.140 61.810 40.310 ;
        RECT 62.900 40.190 63.070 40.360 ;
        RECT 63.260 40.190 63.430 40.360 ;
        RECT 63.700 40.190 63.870 40.360 ;
        RECT 64.440 40.140 64.610 40.310 ;
        RECT 64.800 40.140 64.970 40.310 ;
        RECT 65.160 40.140 65.330 40.310 ;
        RECT 66.000 40.140 66.170 40.310 ;
        RECT 66.360 40.140 66.530 40.310 ;
        RECT 66.720 40.140 66.890 40.310 ;
        RECT 67.640 40.140 67.810 40.310 ;
        RECT 68.000 40.140 68.170 40.310 ;
        RECT 68.360 40.140 68.530 40.310 ;
        RECT 69.620 40.190 69.790 40.360 ;
        RECT 69.980 40.190 70.150 40.360 ;
        RECT 70.420 40.190 70.590 40.360 ;
        RECT 71.160 40.140 71.330 40.310 ;
        RECT 71.520 40.140 71.690 40.310 ;
        RECT 71.880 40.140 72.050 40.310 ;
        RECT 72.720 40.140 72.890 40.310 ;
        RECT 73.080 40.140 73.250 40.310 ;
        RECT 73.440 40.140 73.610 40.310 ;
        RECT 74.360 40.140 74.530 40.310 ;
        RECT 74.720 40.140 74.890 40.310 ;
        RECT 75.080 40.140 75.250 40.310 ;
        RECT 76.340 40.190 76.510 40.360 ;
        RECT 76.700 40.190 76.870 40.360 ;
        RECT 77.140 40.190 77.310 40.360 ;
        RECT 78.980 40.140 79.150 40.310 ;
        RECT 79.340 40.140 79.510 40.310 ;
        RECT 81.140 40.190 81.310 40.360 ;
        RECT 81.500 40.190 81.670 40.360 ;
        RECT 81.940 40.190 82.110 40.360 ;
        RECT 82.680 40.140 82.850 40.310 ;
        RECT 83.040 40.140 83.210 40.310 ;
        RECT 83.400 40.140 83.570 40.310 ;
        RECT 84.240 40.140 84.410 40.310 ;
        RECT 84.600 40.140 84.770 40.310 ;
        RECT 84.960 40.140 85.130 40.310 ;
        RECT 85.880 40.140 86.050 40.310 ;
        RECT 86.240 40.140 86.410 40.310 ;
        RECT 86.600 40.140 86.770 40.310 ;
        RECT 87.860 40.190 88.030 40.360 ;
        RECT 88.220 40.190 88.390 40.360 ;
        RECT 88.660 40.190 88.830 40.360 ;
        RECT 89.400 40.140 89.570 40.310 ;
        RECT 89.760 40.140 89.930 40.310 ;
        RECT 90.120 40.140 90.290 40.310 ;
        RECT 90.960 40.140 91.130 40.310 ;
        RECT 91.320 40.140 91.490 40.310 ;
        RECT 91.680 40.140 91.850 40.310 ;
        RECT 92.600 40.140 92.770 40.310 ;
        RECT 92.960 40.140 93.130 40.310 ;
        RECT 93.320 40.140 93.490 40.310 ;
        RECT 94.580 40.190 94.750 40.360 ;
        RECT 94.940 40.190 95.110 40.360 ;
        RECT 95.380 40.190 95.550 40.360 ;
        RECT 96.100 40.140 96.270 40.310 ;
        RECT 96.460 40.140 96.630 40.310 ;
        RECT 96.820 40.140 96.990 40.310 ;
        RECT 97.180 40.140 97.350 40.310 ;
        RECT 98.340 40.140 98.510 40.310 ;
        RECT 98.700 40.140 98.870 40.310 ;
        RECT 99.060 40.140 99.230 40.310 ;
        RECT 99.420 40.140 99.590 40.310 ;
        RECT 100.340 40.190 100.510 40.360 ;
        RECT 100.700 40.190 100.870 40.360 ;
        RECT 101.140 40.190 101.310 40.360 ;
        RECT 101.880 40.140 102.050 40.310 ;
        RECT 102.240 40.140 102.410 40.310 ;
        RECT 102.600 40.140 102.770 40.310 ;
        RECT 102.960 40.140 103.130 40.310 ;
        RECT 103.320 40.140 103.490 40.310 ;
        RECT 105.620 40.190 105.790 40.360 ;
        RECT 105.980 40.190 106.150 40.360 ;
        RECT 106.420 40.190 106.590 40.360 ;
        RECT 107.160 40.140 107.330 40.310 ;
        RECT 107.520 40.140 107.690 40.310 ;
        RECT 108.980 40.190 109.150 40.360 ;
        RECT 109.340 40.190 109.510 40.360 ;
        RECT 109.780 40.190 109.950 40.360 ;
        RECT 111.000 40.140 111.170 40.310 ;
        RECT 111.360 40.140 111.530 40.310 ;
        RECT 111.720 40.140 111.890 40.310 ;
        RECT 112.560 40.140 112.730 40.310 ;
        RECT 112.920 40.140 113.090 40.310 ;
        RECT 113.280 40.140 113.450 40.310 ;
        RECT 114.200 40.140 114.370 40.310 ;
        RECT 114.560 40.140 114.730 40.310 ;
        RECT 114.920 40.140 115.090 40.310 ;
        RECT 116.390 40.190 116.560 40.360 ;
        RECT 116.830 40.190 117.000 40.360 ;
        RECT 117.240 40.190 117.410 40.360 ;
        RECT 117.670 40.190 117.840 40.360 ;
        RECT 118.110 40.190 118.280 40.360 ;
        RECT 118.520 40.190 118.690 40.360 ;
        RECT 120.600 40.140 120.770 40.310 ;
        RECT 120.960 40.140 121.130 40.310 ;
        RECT 121.320 40.140 121.490 40.310 ;
        RECT 122.160 40.140 122.330 40.310 ;
        RECT 122.520 40.140 122.690 40.310 ;
        RECT 122.880 40.140 123.050 40.310 ;
        RECT 123.800 40.140 123.970 40.310 ;
        RECT 124.160 40.140 124.330 40.310 ;
        RECT 124.520 40.140 124.690 40.310 ;
        RECT 125.780 40.190 125.950 40.360 ;
        RECT 126.140 40.190 126.310 40.360 ;
        RECT 126.580 40.190 126.750 40.360 ;
        RECT 127.980 40.140 128.150 40.310 ;
        RECT 128.340 40.140 128.510 40.310 ;
        RECT 128.700 40.140 128.870 40.310 ;
        RECT 129.060 40.140 129.230 40.310 ;
        RECT 130.170 40.140 130.340 40.310 ;
        RECT 130.530 40.140 130.700 40.310 ;
        RECT 130.890 40.140 131.060 40.310 ;
        RECT 131.250 40.140 131.420 40.310 ;
        RECT 132.020 40.190 132.190 40.360 ;
        RECT 132.380 40.190 132.550 40.360 ;
        RECT 132.820 40.190 132.990 40.360 ;
        RECT 134.180 40.140 134.350 40.310 ;
        RECT 134.540 40.140 134.710 40.310 ;
        RECT 136.340 40.190 136.510 40.360 ;
        RECT 136.700 40.190 136.870 40.360 ;
        RECT 137.140 40.190 137.310 40.360 ;
        RECT 138.040 40.140 138.210 40.310 ;
        RECT 138.400 40.140 138.570 40.310 ;
        RECT 140.660 40.190 140.830 40.360 ;
        RECT 141.020 40.190 141.190 40.360 ;
        RECT 141.460 40.190 141.630 40.360 ;
        RECT 6.470 32.900 6.640 33.070 ;
        RECT 6.910 32.900 7.080 33.070 ;
        RECT 7.320 32.900 7.490 33.070 ;
        RECT 7.750 32.900 7.920 33.070 ;
        RECT 8.190 32.900 8.360 33.070 ;
        RECT 8.600 32.900 8.770 33.070 ;
        RECT 10.680 32.950 10.850 33.120 ;
        RECT 11.040 32.950 11.210 33.120 ;
        RECT 12.500 32.900 12.670 33.070 ;
        RECT 12.860 32.900 13.030 33.070 ;
        RECT 13.300 32.900 13.470 33.070 ;
        RECT 14.660 32.950 14.830 33.120 ;
        RECT 15.020 32.950 15.190 33.120 ;
        RECT 17.030 32.900 17.200 33.070 ;
        RECT 17.470 32.900 17.640 33.070 ;
        RECT 17.880 32.900 18.050 33.070 ;
        RECT 18.310 32.900 18.480 33.070 ;
        RECT 18.750 32.900 18.920 33.070 ;
        RECT 19.160 32.900 19.330 33.070 ;
        RECT 21.240 32.950 21.410 33.120 ;
        RECT 21.600 32.950 21.770 33.120 ;
        RECT 21.960 32.950 22.130 33.120 ;
        RECT 22.810 32.950 22.980 33.120 ;
        RECT 23.170 32.950 23.340 33.120 ;
        RECT 24.020 32.900 24.190 33.070 ;
        RECT 24.380 32.900 24.550 33.070 ;
        RECT 24.820 32.900 24.990 33.070 ;
        RECT 25.540 32.950 25.710 33.120 ;
        RECT 25.900 32.950 26.070 33.120 ;
        RECT 26.260 32.950 26.430 33.120 ;
        RECT 26.620 32.950 26.790 33.120 ;
        RECT 27.780 32.950 27.950 33.120 ;
        RECT 28.140 32.950 28.310 33.120 ;
        RECT 28.500 32.950 28.670 33.120 ;
        RECT 28.860 32.950 29.030 33.120 ;
        RECT 29.780 32.900 29.950 33.070 ;
        RECT 30.140 32.900 30.310 33.070 ;
        RECT 30.580 32.900 30.750 33.070 ;
        RECT 31.760 32.950 31.930 33.120 ;
        RECT 32.120 32.950 32.290 33.120 ;
        RECT 32.480 32.950 32.650 33.120 ;
        RECT 32.840 32.950 33.010 33.120 ;
        RECT 33.200 32.950 33.370 33.120 ;
        RECT 33.560 32.950 33.730 33.120 ;
        RECT 33.920 32.950 34.090 33.120 ;
        RECT 34.280 32.950 34.450 33.120 ;
        RECT 35.090 32.950 35.260 33.120 ;
        RECT 35.450 32.950 35.620 33.120 ;
        RECT 35.810 32.950 35.980 33.120 ;
        RECT 36.170 32.950 36.340 33.120 ;
        RECT 37.190 32.900 37.360 33.070 ;
        RECT 37.630 32.900 37.800 33.070 ;
        RECT 38.040 32.900 38.210 33.070 ;
        RECT 38.470 32.900 38.640 33.070 ;
        RECT 38.910 32.900 39.080 33.070 ;
        RECT 39.320 32.900 39.490 33.070 ;
        RECT 40.920 32.950 41.090 33.120 ;
        RECT 41.280 32.950 41.450 33.120 ;
        RECT 41.640 32.950 41.810 33.120 ;
        RECT 42.480 32.950 42.650 33.120 ;
        RECT 42.840 32.950 43.010 33.120 ;
        RECT 43.200 32.950 43.370 33.120 ;
        RECT 44.120 32.950 44.290 33.120 ;
        RECT 44.480 32.950 44.650 33.120 ;
        RECT 44.840 32.950 45.010 33.120 ;
        RECT 46.100 32.900 46.270 33.070 ;
        RECT 46.460 32.900 46.630 33.070 ;
        RECT 46.900 32.900 47.070 33.070 ;
        RECT 47.640 32.950 47.810 33.120 ;
        RECT 48.000 32.950 48.170 33.120 ;
        RECT 48.360 32.950 48.530 33.120 ;
        RECT 49.200 32.950 49.370 33.120 ;
        RECT 49.560 32.950 49.730 33.120 ;
        RECT 49.920 32.950 50.090 33.120 ;
        RECT 50.840 32.950 51.010 33.120 ;
        RECT 51.200 32.950 51.370 33.120 ;
        RECT 51.560 32.950 51.730 33.120 ;
        RECT 52.820 32.900 52.990 33.070 ;
        RECT 53.180 32.900 53.350 33.070 ;
        RECT 53.620 32.900 53.790 33.070 ;
        RECT 54.360 32.950 54.530 33.120 ;
        RECT 54.720 32.950 54.890 33.120 ;
        RECT 55.080 32.950 55.250 33.120 ;
        RECT 55.920 32.950 56.090 33.120 ;
        RECT 56.280 32.950 56.450 33.120 ;
        RECT 56.640 32.950 56.810 33.120 ;
        RECT 57.560 32.950 57.730 33.120 ;
        RECT 57.920 32.950 58.090 33.120 ;
        RECT 58.280 32.950 58.450 33.120 ;
        RECT 59.540 32.900 59.710 33.070 ;
        RECT 59.900 32.900 60.070 33.070 ;
        RECT 60.340 32.900 60.510 33.070 ;
        RECT 61.620 32.950 61.790 33.120 ;
        RECT 61.980 32.950 62.150 33.120 ;
        RECT 64.010 32.950 64.180 33.120 ;
        RECT 66.440 32.950 66.610 33.120 ;
        RECT 66.800 32.950 66.970 33.120 ;
        RECT 67.160 32.950 67.330 33.120 ;
        RECT 68.780 32.950 68.950 33.120 ;
        RECT 69.140 32.950 69.310 33.120 ;
        RECT 69.500 32.950 69.670 33.120 ;
        RECT 71.480 32.950 71.650 33.120 ;
        RECT 71.840 32.950 72.010 33.120 ;
        RECT 72.200 32.950 72.370 33.120 ;
        RECT 73.230 32.950 73.400 33.120 ;
        RECT 73.590 32.950 73.760 33.120 ;
        RECT 73.950 32.950 74.120 33.120 ;
        RECT 74.760 32.950 74.930 33.120 ;
        RECT 75.120 32.950 75.290 33.120 ;
        RECT 75.480 32.950 75.650 33.120 ;
        RECT 76.820 32.900 76.990 33.070 ;
        RECT 77.180 32.900 77.350 33.070 ;
        RECT 77.620 32.900 77.790 33.070 ;
        RECT 78.360 32.950 78.530 33.120 ;
        RECT 78.720 32.950 78.890 33.120 ;
        RECT 80.180 32.900 80.350 33.070 ;
        RECT 80.540 32.900 80.710 33.070 ;
        RECT 80.980 32.900 81.150 33.070 ;
        RECT 81.720 32.950 81.890 33.120 ;
        RECT 82.080 32.950 82.250 33.120 ;
        RECT 82.440 32.950 82.610 33.120 ;
        RECT 83.280 32.950 83.450 33.120 ;
        RECT 83.640 32.950 83.810 33.120 ;
        RECT 84.000 32.950 84.170 33.120 ;
        RECT 84.920 32.950 85.090 33.120 ;
        RECT 85.280 32.950 85.450 33.120 ;
        RECT 85.640 32.950 85.810 33.120 ;
        RECT 86.900 32.900 87.070 33.070 ;
        RECT 87.260 32.900 87.430 33.070 ;
        RECT 87.700 32.900 87.870 33.070 ;
        RECT 89.400 32.950 89.570 33.120 ;
        RECT 89.760 32.950 89.930 33.120 ;
        RECT 90.120 32.950 90.290 33.120 ;
        RECT 90.960 32.950 91.130 33.120 ;
        RECT 91.320 32.950 91.490 33.120 ;
        RECT 91.680 32.950 91.850 33.120 ;
        RECT 92.600 32.950 92.770 33.120 ;
        RECT 92.960 32.950 93.130 33.120 ;
        RECT 93.320 32.950 93.490 33.120 ;
        RECT 94.580 32.900 94.750 33.070 ;
        RECT 94.940 32.900 95.110 33.070 ;
        RECT 95.380 32.900 95.550 33.070 ;
        RECT 96.100 32.950 96.270 33.120 ;
        RECT 96.460 32.950 96.630 33.120 ;
        RECT 96.820 32.950 96.990 33.120 ;
        RECT 97.180 32.950 97.350 33.120 ;
        RECT 98.340 32.950 98.510 33.120 ;
        RECT 98.700 32.950 98.870 33.120 ;
        RECT 99.060 32.950 99.230 33.120 ;
        RECT 99.420 32.950 99.590 33.120 ;
        RECT 100.550 32.900 100.720 33.070 ;
        RECT 100.990 32.900 101.160 33.070 ;
        RECT 101.400 32.900 101.570 33.070 ;
        RECT 101.830 32.900 102.000 33.070 ;
        RECT 102.270 32.900 102.440 33.070 ;
        RECT 102.680 32.900 102.850 33.070 ;
        RECT 105.470 32.950 105.640 33.120 ;
        RECT 105.830 32.950 106.000 33.120 ;
        RECT 106.190 32.950 106.360 33.120 ;
        RECT 106.550 32.950 106.720 33.120 ;
        RECT 106.910 32.950 107.080 33.120 ;
        RECT 107.270 32.950 107.440 33.120 ;
        RECT 108.500 32.900 108.670 33.070 ;
        RECT 108.860 32.900 109.030 33.070 ;
        RECT 109.300 32.900 109.470 33.070 ;
        RECT 110.040 32.950 110.210 33.120 ;
        RECT 110.400 32.950 110.570 33.120 ;
        RECT 110.760 32.950 110.930 33.120 ;
        RECT 111.120 32.950 111.290 33.120 ;
        RECT 111.480 32.950 111.650 33.120 ;
        RECT 113.780 32.900 113.950 33.070 ;
        RECT 114.140 32.900 114.310 33.070 ;
        RECT 114.580 32.900 114.750 33.070 ;
        RECT 116.280 32.950 116.450 33.120 ;
        RECT 116.640 32.950 116.810 33.120 ;
        RECT 117.000 32.950 117.170 33.120 ;
        RECT 117.840 32.950 118.010 33.120 ;
        RECT 118.200 32.950 118.370 33.120 ;
        RECT 118.560 32.950 118.730 33.120 ;
        RECT 119.480 32.950 119.650 33.120 ;
        RECT 119.840 32.950 120.010 33.120 ;
        RECT 120.200 32.950 120.370 33.120 ;
        RECT 121.460 32.900 121.630 33.070 ;
        RECT 121.820 32.900 121.990 33.070 ;
        RECT 122.260 32.900 122.430 33.070 ;
        RECT 124.550 32.950 124.720 33.120 ;
        RECT 124.910 32.950 125.080 33.120 ;
        RECT 125.270 32.950 125.440 33.120 ;
        RECT 125.630 32.950 125.800 33.120 ;
        RECT 125.990 32.950 126.160 33.120 ;
        RECT 127.220 32.900 127.390 33.070 ;
        RECT 127.580 32.900 127.750 33.070 ;
        RECT 128.020 32.900 128.190 33.070 ;
        RECT 128.760 32.950 128.930 33.120 ;
        RECT 129.120 32.950 129.290 33.120 ;
        RECT 129.480 32.950 129.650 33.120 ;
        RECT 129.840 32.950 130.010 33.120 ;
        RECT 130.200 32.950 130.370 33.120 ;
        RECT 131.750 32.900 131.920 33.070 ;
        RECT 132.190 32.900 132.360 33.070 ;
        RECT 132.600 32.900 132.770 33.070 ;
        RECT 133.030 32.900 133.200 33.070 ;
        RECT 133.470 32.900 133.640 33.070 ;
        RECT 133.880 32.900 134.050 33.070 ;
        RECT 135.000 32.950 135.170 33.120 ;
        RECT 135.360 32.950 135.530 33.120 ;
        RECT 136.820 32.900 136.990 33.070 ;
        RECT 137.180 32.900 137.350 33.070 ;
        RECT 137.620 32.900 137.790 33.070 ;
        RECT 138.360 32.950 138.530 33.120 ;
        RECT 138.720 32.950 138.890 33.120 ;
        RECT 140.180 32.900 140.350 33.070 ;
        RECT 140.540 32.900 140.710 33.070 ;
        RECT 140.980 32.900 141.150 33.070 ;
        RECT 5.920 32.470 6.090 32.650 ;
        RECT 6.400 32.470 6.570 32.650 ;
        RECT 6.880 32.470 7.050 32.650 ;
        RECT 7.360 32.470 7.530 32.650 ;
        RECT 7.840 32.470 8.010 32.650 ;
        RECT 8.320 32.470 8.490 32.650 ;
        RECT 8.800 32.470 8.970 32.650 ;
        RECT 9.280 32.470 9.450 32.650 ;
        RECT 9.760 32.470 9.930 32.650 ;
        RECT 10.240 32.470 10.410 32.650 ;
        RECT 10.720 32.470 10.890 32.650 ;
        RECT 11.200 32.470 11.370 32.650 ;
        RECT 11.680 32.470 11.850 32.650 ;
        RECT 12.160 32.470 12.330 32.650 ;
        RECT 12.640 32.470 12.810 32.650 ;
        RECT 13.120 32.470 13.290 32.650 ;
        RECT 13.600 32.470 13.770 32.650 ;
        RECT 14.080 32.470 14.250 32.650 ;
        RECT 14.560 32.470 14.730 32.650 ;
        RECT 15.040 32.470 15.210 32.650 ;
        RECT 15.520 32.470 15.690 32.650 ;
        RECT 16.000 32.470 16.170 32.650 ;
        RECT 16.480 32.470 16.650 32.650 ;
        RECT 16.960 32.470 17.130 32.650 ;
        RECT 17.440 32.470 17.610 32.650 ;
        RECT 17.920 32.470 18.090 32.650 ;
        RECT 18.400 32.470 18.570 32.650 ;
        RECT 18.880 32.470 19.050 32.650 ;
        RECT 19.360 32.470 19.530 32.650 ;
        RECT 19.840 32.470 20.010 32.650 ;
        RECT 20.320 32.470 20.490 32.650 ;
        RECT 20.800 32.470 20.970 32.650 ;
        RECT 21.280 32.470 21.450 32.650 ;
        RECT 21.760 32.470 21.930 32.650 ;
        RECT 22.240 32.470 22.410 32.650 ;
        RECT 22.720 32.470 22.890 32.650 ;
        RECT 23.200 32.470 23.370 32.650 ;
        RECT 23.680 32.470 23.850 32.650 ;
        RECT 24.160 32.470 24.330 32.650 ;
        RECT 24.640 32.470 24.810 32.650 ;
        RECT 25.120 32.470 25.290 32.650 ;
        RECT 25.600 32.470 25.770 32.650 ;
        RECT 26.080 32.470 26.250 32.650 ;
        RECT 26.560 32.470 26.730 32.650 ;
        RECT 27.040 32.470 27.210 32.650 ;
        RECT 27.520 32.470 27.690 32.650 ;
        RECT 28.000 32.470 28.170 32.650 ;
        RECT 28.480 32.470 28.650 32.650 ;
        RECT 28.960 32.470 29.130 32.650 ;
        RECT 29.440 32.470 29.610 32.650 ;
        RECT 29.920 32.470 30.090 32.650 ;
        RECT 30.400 32.470 30.570 32.650 ;
        RECT 30.880 32.470 31.050 32.650 ;
        RECT 31.360 32.470 31.530 32.650 ;
        RECT 31.840 32.470 32.010 32.650 ;
        RECT 32.320 32.470 32.490 32.650 ;
        RECT 32.800 32.470 32.970 32.650 ;
        RECT 33.280 32.470 33.450 32.650 ;
        RECT 33.760 32.470 33.930 32.650 ;
        RECT 34.240 32.470 34.410 32.650 ;
        RECT 34.720 32.470 34.890 32.650 ;
        RECT 35.200 32.470 35.370 32.650 ;
        RECT 35.680 32.470 35.850 32.650 ;
        RECT 36.160 32.470 36.330 32.650 ;
        RECT 36.640 32.470 36.810 32.650 ;
        RECT 37.120 32.470 37.290 32.650 ;
        RECT 37.600 32.470 37.770 32.650 ;
        RECT 38.080 32.470 38.250 32.650 ;
        RECT 38.560 32.470 38.730 32.650 ;
        RECT 39.040 32.470 39.210 32.650 ;
        RECT 39.520 32.470 39.690 32.650 ;
        RECT 40.000 32.470 40.170 32.650 ;
        RECT 40.480 32.640 40.650 32.650 ;
      LAYER li1 ;
        RECT 40.320 32.470 40.800 32.640 ;
      LAYER li1 ;
        RECT 40.960 32.470 41.130 32.650 ;
        RECT 41.440 32.470 41.610 32.650 ;
        RECT 41.920 32.470 42.090 32.650 ;
        RECT 42.400 32.470 42.570 32.650 ;
        RECT 42.880 32.470 43.050 32.650 ;
        RECT 43.360 32.470 43.530 32.650 ;
        RECT 43.840 32.470 44.010 32.650 ;
        RECT 44.320 32.470 44.490 32.650 ;
        RECT 44.800 32.470 44.970 32.650 ;
        RECT 45.280 32.470 45.450 32.650 ;
        RECT 45.760 32.470 45.930 32.650 ;
        RECT 46.240 32.470 46.410 32.650 ;
        RECT 46.720 32.470 46.890 32.650 ;
        RECT 47.200 32.470 47.370 32.650 ;
        RECT 47.680 32.470 47.850 32.650 ;
        RECT 48.160 32.470 48.330 32.650 ;
        RECT 48.640 32.470 48.810 32.650 ;
        RECT 49.120 32.470 49.290 32.650 ;
        RECT 49.600 32.470 49.770 32.650 ;
        RECT 50.080 32.470 50.250 32.650 ;
        RECT 50.560 32.470 50.730 32.650 ;
        RECT 51.040 32.470 51.210 32.650 ;
        RECT 51.520 32.470 51.690 32.650 ;
        RECT 52.000 32.470 52.170 32.650 ;
        RECT 52.480 32.470 52.650 32.650 ;
        RECT 52.960 32.470 53.130 32.650 ;
        RECT 53.440 32.470 53.610 32.650 ;
        RECT 53.920 32.470 54.090 32.650 ;
        RECT 54.400 32.470 54.570 32.650 ;
        RECT 54.880 32.470 55.050 32.650 ;
        RECT 55.360 32.470 55.530 32.650 ;
        RECT 55.840 32.470 56.010 32.650 ;
        RECT 56.320 32.470 56.490 32.650 ;
        RECT 56.800 32.470 56.970 32.650 ;
        RECT 57.280 32.470 57.450 32.650 ;
        RECT 57.760 32.470 57.930 32.650 ;
        RECT 58.240 32.470 58.410 32.650 ;
        RECT 58.720 32.470 58.890 32.650 ;
        RECT 59.200 32.470 59.370 32.650 ;
        RECT 59.680 32.470 59.850 32.650 ;
        RECT 60.160 32.470 60.330 32.650 ;
        RECT 60.640 32.470 60.810 32.650 ;
        RECT 61.120 32.470 61.290 32.650 ;
        RECT 61.600 32.470 61.770 32.650 ;
        RECT 62.080 32.470 62.250 32.650 ;
        RECT 62.560 32.470 62.730 32.650 ;
        RECT 63.040 32.470 63.210 32.650 ;
        RECT 63.520 32.470 63.690 32.650 ;
        RECT 64.000 32.470 64.170 32.650 ;
        RECT 64.480 32.470 64.650 32.650 ;
        RECT 64.960 32.470 65.130 32.650 ;
        RECT 65.440 32.470 65.610 32.650 ;
        RECT 65.920 32.470 66.090 32.650 ;
        RECT 66.400 32.470 66.570 32.650 ;
        RECT 66.880 32.470 67.050 32.650 ;
        RECT 67.360 32.470 67.530 32.650 ;
        RECT 67.840 32.470 68.010 32.650 ;
        RECT 68.320 32.470 68.490 32.650 ;
        RECT 68.800 32.470 68.970 32.650 ;
        RECT 69.280 32.470 69.450 32.650 ;
        RECT 69.760 32.470 69.930 32.650 ;
        RECT 70.240 32.470 70.410 32.650 ;
        RECT 70.720 32.470 70.890 32.650 ;
        RECT 71.200 32.470 71.370 32.650 ;
        RECT 71.680 32.470 71.850 32.650 ;
        RECT 72.160 32.470 72.330 32.650 ;
        RECT 72.640 32.470 72.810 32.650 ;
        RECT 73.120 32.470 73.290 32.650 ;
        RECT 73.600 32.470 73.770 32.650 ;
        RECT 74.080 32.470 74.250 32.650 ;
        RECT 74.560 32.470 74.730 32.650 ;
        RECT 75.040 32.470 75.210 32.650 ;
        RECT 75.520 32.470 75.690 32.650 ;
        RECT 76.000 32.470 76.170 32.650 ;
        RECT 76.480 32.470 76.650 32.650 ;
        RECT 76.960 32.470 77.130 32.650 ;
        RECT 77.440 32.470 77.610 32.650 ;
        RECT 77.920 32.470 78.090 32.650 ;
        RECT 78.400 32.470 78.570 32.650 ;
        RECT 78.880 32.470 79.050 32.650 ;
        RECT 79.360 32.470 79.530 32.650 ;
        RECT 79.840 32.470 80.010 32.650 ;
        RECT 80.320 32.470 80.490 32.650 ;
        RECT 80.800 32.470 80.970 32.650 ;
        RECT 81.280 32.470 81.450 32.650 ;
        RECT 81.760 32.470 81.930 32.650 ;
        RECT 82.240 32.470 82.410 32.650 ;
        RECT 82.720 32.470 82.890 32.650 ;
        RECT 83.200 32.470 83.370 32.650 ;
        RECT 83.680 32.470 83.850 32.650 ;
        RECT 84.160 32.470 84.330 32.650 ;
        RECT 84.640 32.470 84.810 32.650 ;
        RECT 85.120 32.470 85.290 32.650 ;
        RECT 85.600 32.470 85.770 32.650 ;
        RECT 86.080 32.470 86.250 32.650 ;
        RECT 86.560 32.470 86.730 32.650 ;
        RECT 87.040 32.470 87.210 32.650 ;
        RECT 87.520 32.470 87.690 32.650 ;
        RECT 88.000 32.470 88.170 32.650 ;
        RECT 88.480 32.470 88.650 32.650 ;
        RECT 88.960 32.470 89.130 32.650 ;
        RECT 89.440 32.470 89.610 32.650 ;
        RECT 89.920 32.470 90.090 32.650 ;
        RECT 90.400 32.470 90.570 32.650 ;
        RECT 90.880 32.470 91.050 32.650 ;
        RECT 91.360 32.470 91.530 32.650 ;
        RECT 91.840 32.470 92.010 32.650 ;
        RECT 92.320 32.470 92.490 32.650 ;
        RECT 92.800 32.470 92.970 32.650 ;
        RECT 93.280 32.470 93.450 32.650 ;
        RECT 93.760 32.470 93.930 32.650 ;
        RECT 94.240 32.470 94.410 32.650 ;
        RECT 94.720 32.470 94.890 32.650 ;
        RECT 95.200 32.470 95.370 32.650 ;
        RECT 95.680 32.470 95.850 32.650 ;
        RECT 96.160 32.470 96.330 32.650 ;
        RECT 96.640 32.470 96.810 32.650 ;
        RECT 97.120 32.470 97.290 32.650 ;
        RECT 97.600 32.470 97.770 32.650 ;
        RECT 98.080 32.470 98.250 32.650 ;
        RECT 98.560 32.470 98.730 32.650 ;
        RECT 99.040 32.470 99.210 32.650 ;
        RECT 99.520 32.470 99.690 32.650 ;
        RECT 100.000 32.470 100.170 32.650 ;
        RECT 100.480 32.470 100.650 32.650 ;
        RECT 100.960 32.470 101.130 32.650 ;
        RECT 101.440 32.470 101.610 32.650 ;
        RECT 101.920 32.470 102.090 32.650 ;
        RECT 102.400 32.470 102.570 32.650 ;
        RECT 102.880 32.470 103.050 32.650 ;
        RECT 103.360 32.470 103.530 32.650 ;
        RECT 103.840 32.470 104.010 32.650 ;
      LAYER li1 ;
        RECT 104.160 32.640 104.640 32.650 ;
      LAYER li1 ;
        RECT 104.320 32.470 104.490 32.640 ;
        RECT 104.800 32.470 104.970 32.650 ;
        RECT 105.280 32.470 105.450 32.650 ;
        RECT 105.760 32.470 105.930 32.650 ;
        RECT 106.240 32.470 106.410 32.650 ;
        RECT 106.720 32.470 106.890 32.650 ;
        RECT 107.200 32.470 107.370 32.650 ;
        RECT 107.680 32.470 107.850 32.650 ;
        RECT 108.160 32.470 108.330 32.650 ;
        RECT 108.640 32.470 108.810 32.650 ;
        RECT 109.120 32.470 109.290 32.650 ;
        RECT 109.600 32.470 109.770 32.650 ;
        RECT 110.080 32.470 110.250 32.650 ;
        RECT 110.560 32.470 110.730 32.650 ;
        RECT 111.040 32.470 111.210 32.650 ;
        RECT 111.520 32.470 111.690 32.650 ;
        RECT 112.000 32.470 112.170 32.650 ;
        RECT 112.480 32.470 112.650 32.650 ;
        RECT 112.960 32.470 113.130 32.650 ;
        RECT 113.440 32.470 113.610 32.650 ;
        RECT 113.920 32.470 114.090 32.650 ;
        RECT 114.400 32.470 114.570 32.650 ;
        RECT 114.880 32.470 115.050 32.650 ;
        RECT 115.360 32.470 115.530 32.650 ;
        RECT 115.840 32.470 116.010 32.650 ;
        RECT 116.320 32.470 116.490 32.650 ;
        RECT 116.800 32.470 116.970 32.650 ;
        RECT 117.280 32.470 117.450 32.650 ;
        RECT 117.760 32.470 117.930 32.650 ;
        RECT 118.240 32.470 118.410 32.650 ;
        RECT 118.720 32.470 118.890 32.650 ;
        RECT 119.200 32.470 119.370 32.650 ;
      LAYER li1 ;
        RECT 119.520 32.640 120.000 32.650 ;
      LAYER li1 ;
        RECT 119.680 32.470 119.850 32.640 ;
        RECT 120.160 32.470 120.330 32.650 ;
        RECT 120.640 32.470 120.810 32.650 ;
        RECT 121.120 32.470 121.290 32.650 ;
        RECT 121.600 32.470 121.770 32.650 ;
        RECT 122.080 32.470 122.250 32.650 ;
        RECT 122.560 32.470 122.730 32.650 ;
        RECT 123.040 32.470 123.210 32.650 ;
        RECT 123.520 32.470 123.690 32.650 ;
        RECT 124.000 32.470 124.170 32.650 ;
        RECT 124.480 32.470 124.650 32.650 ;
        RECT 124.960 32.470 125.130 32.650 ;
        RECT 125.440 32.470 125.610 32.650 ;
        RECT 125.920 32.470 126.090 32.650 ;
        RECT 126.400 32.470 126.570 32.650 ;
        RECT 126.880 32.470 127.050 32.650 ;
        RECT 127.360 32.470 127.530 32.650 ;
        RECT 127.840 32.470 128.010 32.650 ;
        RECT 128.320 32.470 128.490 32.650 ;
        RECT 128.800 32.470 128.970 32.650 ;
        RECT 129.280 32.470 129.450 32.650 ;
        RECT 129.760 32.470 129.930 32.650 ;
        RECT 130.240 32.470 130.410 32.650 ;
        RECT 130.720 32.470 130.890 32.650 ;
        RECT 131.200 32.470 131.370 32.650 ;
        RECT 131.680 32.470 131.850 32.650 ;
      LAYER li1 ;
        RECT 132.000 32.640 132.480 32.650 ;
      LAYER li1 ;
        RECT 132.160 32.470 132.330 32.640 ;
        RECT 132.640 32.470 132.810 32.650 ;
        RECT 133.120 32.470 133.290 32.650 ;
        RECT 133.600 32.470 133.770 32.650 ;
        RECT 134.080 32.470 134.250 32.650 ;
        RECT 134.560 32.470 134.730 32.650 ;
        RECT 135.040 32.470 135.210 32.650 ;
        RECT 135.520 32.470 135.690 32.650 ;
        RECT 136.000 32.470 136.170 32.650 ;
        RECT 136.480 32.470 136.650 32.650 ;
        RECT 136.960 32.470 137.130 32.650 ;
        RECT 137.440 32.470 137.610 32.650 ;
        RECT 137.920 32.470 138.090 32.650 ;
        RECT 138.400 32.470 138.570 32.650 ;
        RECT 138.880 32.470 139.050 32.650 ;
        RECT 139.360 32.470 139.530 32.650 ;
        RECT 139.840 32.470 140.010 32.650 ;
        RECT 140.320 32.470 140.490 32.650 ;
        RECT 140.800 32.470 140.970 32.650 ;
        RECT 141.280 32.470 141.450 32.650 ;
      LAYER li1 ;
        RECT 141.600 32.470 142.080 32.650 ;
      LAYER li1 ;
        RECT 7.380 32.000 7.550 32.170 ;
        RECT 7.740 32.000 7.910 32.170 ;
        RECT 9.770 32.000 9.940 32.170 ;
        RECT 12.200 32.000 12.370 32.170 ;
        RECT 12.560 32.000 12.730 32.170 ;
        RECT 12.920 32.000 13.090 32.170 ;
        RECT 14.540 32.000 14.710 32.170 ;
        RECT 14.900 32.000 15.070 32.170 ;
        RECT 15.260 32.000 15.430 32.170 ;
        RECT 17.240 32.000 17.410 32.170 ;
        RECT 17.600 32.000 17.770 32.170 ;
        RECT 17.960 32.000 18.130 32.170 ;
        RECT 18.990 32.000 19.160 32.170 ;
        RECT 19.350 32.000 19.520 32.170 ;
        RECT 19.710 32.000 19.880 32.170 ;
        RECT 20.520 32.000 20.690 32.170 ;
        RECT 20.880 32.000 21.050 32.170 ;
        RECT 21.240 32.000 21.410 32.170 ;
        RECT 22.580 32.050 22.750 32.220 ;
        RECT 22.940 32.050 23.110 32.220 ;
        RECT 23.380 32.050 23.550 32.220 ;
        RECT 24.120 32.000 24.290 32.170 ;
        RECT 24.480 32.000 24.650 32.170 ;
        RECT 25.940 32.050 26.110 32.220 ;
        RECT 26.300 32.050 26.470 32.220 ;
        RECT 26.740 32.050 26.910 32.220 ;
        RECT 28.050 32.000 28.220 32.170 ;
        RECT 28.410 32.000 28.580 32.170 ;
        RECT 28.770 32.000 28.940 32.170 ;
        RECT 29.130 32.000 29.300 32.170 ;
        RECT 31.220 32.050 31.390 32.220 ;
        RECT 31.580 32.050 31.750 32.220 ;
        RECT 32.020 32.050 32.190 32.220 ;
        RECT 33.330 32.000 33.500 32.170 ;
        RECT 33.690 32.000 33.860 32.170 ;
        RECT 34.050 32.000 34.220 32.170 ;
        RECT 34.410 32.000 34.580 32.170 ;
        RECT 36.500 32.050 36.670 32.220 ;
        RECT 36.860 32.050 37.030 32.220 ;
        RECT 37.300 32.050 37.470 32.220 ;
        RECT 38.980 32.000 39.150 32.170 ;
        RECT 39.340 32.000 39.510 32.170 ;
        RECT 39.700 32.000 39.870 32.170 ;
        RECT 40.060 32.000 40.230 32.170 ;
        RECT 41.220 32.000 41.390 32.170 ;
        RECT 41.580 32.000 41.750 32.170 ;
        RECT 41.940 32.000 42.110 32.170 ;
        RECT 42.300 32.000 42.470 32.170 ;
        RECT 43.220 32.050 43.390 32.220 ;
        RECT 43.580 32.050 43.750 32.220 ;
        RECT 44.020 32.050 44.190 32.220 ;
        RECT 44.760 32.000 44.930 32.170 ;
        RECT 45.120 32.000 45.290 32.170 ;
        RECT 45.480 32.000 45.650 32.170 ;
        RECT 46.320 32.000 46.490 32.170 ;
        RECT 46.680 32.000 46.850 32.170 ;
        RECT 47.040 32.000 47.210 32.170 ;
        RECT 47.960 32.000 48.130 32.170 ;
        RECT 48.320 32.000 48.490 32.170 ;
        RECT 48.680 32.000 48.850 32.170 ;
        RECT 49.940 32.050 50.110 32.220 ;
        RECT 50.300 32.050 50.470 32.220 ;
        RECT 50.740 32.050 50.910 32.220 ;
        RECT 51.480 32.000 51.650 32.170 ;
        RECT 51.840 32.000 52.010 32.170 ;
        RECT 52.200 32.000 52.370 32.170 ;
        RECT 53.040 32.000 53.210 32.170 ;
        RECT 53.400 32.000 53.570 32.170 ;
        RECT 53.760 32.000 53.930 32.170 ;
        RECT 54.680 32.000 54.850 32.170 ;
        RECT 55.040 32.000 55.210 32.170 ;
        RECT 55.400 32.000 55.570 32.170 ;
        RECT 56.870 32.050 57.040 32.220 ;
        RECT 57.310 32.050 57.480 32.220 ;
        RECT 57.720 32.050 57.890 32.220 ;
        RECT 58.150 32.050 58.320 32.220 ;
        RECT 58.590 32.050 58.760 32.220 ;
        RECT 59.000 32.050 59.170 32.220 ;
        RECT 60.120 32.000 60.290 32.170 ;
        RECT 60.480 32.000 60.650 32.170 ;
        RECT 60.840 32.000 61.010 32.170 ;
        RECT 61.680 32.000 61.850 32.170 ;
        RECT 62.040 32.000 62.210 32.170 ;
        RECT 62.400 32.000 62.570 32.170 ;
        RECT 63.320 32.000 63.490 32.170 ;
        RECT 63.680 32.000 63.850 32.170 ;
        RECT 64.040 32.000 64.210 32.170 ;
        RECT 65.300 32.050 65.470 32.220 ;
        RECT 65.660 32.050 65.830 32.220 ;
        RECT 66.100 32.050 66.270 32.220 ;
        RECT 66.840 32.000 67.010 32.170 ;
        RECT 67.200 32.000 67.370 32.170 ;
        RECT 67.560 32.000 67.730 32.170 ;
        RECT 68.400 32.000 68.570 32.170 ;
        RECT 68.760 32.000 68.930 32.170 ;
        RECT 69.120 32.000 69.290 32.170 ;
        RECT 70.040 32.000 70.210 32.170 ;
        RECT 70.400 32.000 70.570 32.170 ;
        RECT 70.760 32.000 70.930 32.170 ;
        RECT 72.020 32.050 72.190 32.220 ;
        RECT 72.380 32.050 72.550 32.220 ;
        RECT 72.820 32.050 72.990 32.220 ;
        RECT 73.560 32.000 73.730 32.170 ;
        RECT 73.920 32.000 74.090 32.170 ;
        RECT 74.280 32.000 74.450 32.170 ;
        RECT 75.120 32.000 75.290 32.170 ;
        RECT 75.480 32.000 75.650 32.170 ;
        RECT 75.840 32.000 76.010 32.170 ;
        RECT 76.760 32.000 76.930 32.170 ;
        RECT 77.120 32.000 77.290 32.170 ;
        RECT 77.480 32.000 77.650 32.170 ;
        RECT 78.740 32.050 78.910 32.220 ;
        RECT 79.100 32.050 79.270 32.220 ;
        RECT 79.540 32.050 79.710 32.220 ;
        RECT 80.260 32.000 80.430 32.170 ;
        RECT 80.620 32.000 80.790 32.170 ;
        RECT 80.980 32.000 81.150 32.170 ;
        RECT 81.340 32.000 81.510 32.170 ;
        RECT 82.500 32.000 82.670 32.170 ;
        RECT 82.860 32.000 83.030 32.170 ;
        RECT 83.220 32.000 83.390 32.170 ;
        RECT 83.580 32.000 83.750 32.170 ;
        RECT 84.500 32.050 84.670 32.220 ;
        RECT 84.860 32.050 85.030 32.220 ;
        RECT 85.300 32.050 85.470 32.220 ;
        RECT 86.020 32.000 86.190 32.170 ;
        RECT 86.380 32.000 86.550 32.170 ;
        RECT 86.740 32.000 86.910 32.170 ;
        RECT 87.100 32.000 87.270 32.170 ;
        RECT 88.260 32.000 88.430 32.170 ;
        RECT 88.620 32.000 88.790 32.170 ;
        RECT 88.980 32.000 89.150 32.170 ;
        RECT 89.340 32.000 89.510 32.170 ;
        RECT 90.260 32.050 90.430 32.220 ;
        RECT 90.620 32.050 90.790 32.220 ;
        RECT 91.060 32.050 91.230 32.220 ;
        RECT 92.240 32.000 92.410 32.170 ;
        RECT 92.600 32.000 92.770 32.170 ;
        RECT 92.960 32.000 93.130 32.170 ;
        RECT 93.320 32.000 93.490 32.170 ;
        RECT 93.680 32.000 93.850 32.170 ;
        RECT 94.040 32.000 94.210 32.170 ;
        RECT 94.400 32.000 94.570 32.170 ;
        RECT 94.760 32.000 94.930 32.170 ;
        RECT 95.570 32.000 95.740 32.170 ;
        RECT 95.930 32.000 96.100 32.170 ;
        RECT 96.290 32.000 96.460 32.170 ;
        RECT 96.650 32.000 96.820 32.170 ;
        RECT 97.460 32.050 97.630 32.220 ;
        RECT 97.820 32.050 97.990 32.220 ;
        RECT 98.260 32.050 98.430 32.220 ;
        RECT 99.710 32.000 99.880 32.170 ;
        RECT 100.070 32.000 100.240 32.170 ;
        RECT 100.430 32.000 100.600 32.170 ;
        RECT 100.790 32.000 100.960 32.170 ;
        RECT 101.150 32.000 101.320 32.170 ;
        RECT 101.510 32.000 101.680 32.170 ;
        RECT 102.740 32.050 102.910 32.220 ;
        RECT 103.100 32.050 103.270 32.220 ;
        RECT 103.540 32.050 103.710 32.220 ;
        RECT 104.740 32.000 104.910 32.170 ;
        RECT 105.100 32.000 105.270 32.170 ;
        RECT 105.460 32.000 105.630 32.170 ;
        RECT 105.820 32.000 105.990 32.170 ;
        RECT 106.980 32.000 107.150 32.170 ;
        RECT 107.340 32.000 107.510 32.170 ;
        RECT 107.700 32.000 107.870 32.170 ;
        RECT 108.060 32.000 108.230 32.170 ;
        RECT 108.980 32.050 109.150 32.220 ;
        RECT 109.340 32.050 109.510 32.220 ;
        RECT 109.780 32.050 109.950 32.220 ;
        RECT 110.960 32.000 111.130 32.170 ;
        RECT 111.320 32.000 111.490 32.170 ;
        RECT 111.680 32.000 111.850 32.170 ;
        RECT 112.040 32.000 112.210 32.170 ;
        RECT 112.400 32.000 112.570 32.170 ;
        RECT 112.760 32.000 112.930 32.170 ;
        RECT 113.120 32.000 113.290 32.170 ;
        RECT 113.480 32.000 113.650 32.170 ;
        RECT 114.290 32.000 114.460 32.170 ;
        RECT 114.650 32.000 114.820 32.170 ;
        RECT 115.010 32.000 115.180 32.170 ;
        RECT 115.370 32.000 115.540 32.170 ;
        RECT 116.390 32.050 116.560 32.220 ;
        RECT 116.830 32.050 117.000 32.220 ;
        RECT 117.240 32.050 117.410 32.220 ;
        RECT 117.670 32.050 117.840 32.220 ;
        RECT 118.110 32.050 118.280 32.220 ;
        RECT 118.520 32.050 118.690 32.220 ;
        RECT 120.100 32.000 120.270 32.170 ;
        RECT 120.460 32.000 120.630 32.170 ;
        RECT 120.820 32.000 120.990 32.170 ;
        RECT 121.180 32.000 121.350 32.170 ;
        RECT 122.340 32.000 122.510 32.170 ;
        RECT 122.700 32.000 122.870 32.170 ;
        RECT 123.060 32.000 123.230 32.170 ;
        RECT 123.420 32.000 123.590 32.170 ;
        RECT 124.340 32.050 124.510 32.220 ;
        RECT 124.700 32.050 124.870 32.220 ;
        RECT 125.140 32.050 125.310 32.220 ;
        RECT 125.880 32.000 126.050 32.170 ;
        RECT 126.240 32.000 126.410 32.170 ;
        RECT 126.600 32.000 126.770 32.170 ;
        RECT 127.450 32.000 127.620 32.170 ;
        RECT 127.810 32.000 127.980 32.170 ;
        RECT 128.870 32.050 129.040 32.220 ;
        RECT 129.310 32.050 129.480 32.220 ;
        RECT 129.720 32.050 129.890 32.220 ;
        RECT 130.150 32.050 130.320 32.220 ;
        RECT 130.590 32.050 130.760 32.220 ;
        RECT 131.000 32.050 131.170 32.220 ;
        RECT 132.600 32.000 132.770 32.170 ;
        RECT 132.960 32.000 133.130 32.170 ;
        RECT 134.630 32.050 134.800 32.220 ;
        RECT 135.070 32.050 135.240 32.220 ;
        RECT 135.480 32.050 135.650 32.220 ;
        RECT 135.910 32.050 136.080 32.220 ;
        RECT 136.350 32.050 136.520 32.220 ;
        RECT 136.760 32.050 136.930 32.220 ;
        RECT 138.470 32.050 138.640 32.220 ;
        RECT 138.910 32.050 139.080 32.220 ;
        RECT 139.320 32.050 139.490 32.220 ;
        RECT 139.750 32.050 139.920 32.220 ;
        RECT 140.190 32.050 140.360 32.220 ;
        RECT 140.600 32.050 140.770 32.220 ;
        RECT 6.470 24.760 6.640 24.930 ;
        RECT 6.910 24.760 7.080 24.930 ;
        RECT 7.320 24.760 7.490 24.930 ;
        RECT 7.750 24.760 7.920 24.930 ;
        RECT 8.190 24.760 8.360 24.930 ;
        RECT 8.600 24.760 8.770 24.930 ;
        RECT 10.310 24.760 10.480 24.930 ;
        RECT 10.750 24.760 10.920 24.930 ;
        RECT 11.160 24.760 11.330 24.930 ;
        RECT 11.590 24.760 11.760 24.930 ;
        RECT 12.030 24.760 12.200 24.930 ;
        RECT 12.440 24.760 12.610 24.930 ;
        RECT 15.000 24.810 15.170 24.980 ;
        RECT 15.360 24.810 15.530 24.980 ;
        RECT 16.820 24.760 16.990 24.930 ;
        RECT 17.180 24.760 17.350 24.930 ;
        RECT 17.620 24.760 17.790 24.930 ;
        RECT 18.360 24.810 18.530 24.980 ;
        RECT 18.720 24.810 18.890 24.980 ;
        RECT 19.080 24.810 19.250 24.980 ;
        RECT 19.440 24.810 19.610 24.980 ;
        RECT 19.800 24.810 19.970 24.980 ;
        RECT 21.140 24.760 21.310 24.930 ;
        RECT 21.500 24.760 21.670 24.930 ;
        RECT 21.940 24.760 22.110 24.930 ;
        RECT 23.300 24.810 23.470 24.980 ;
        RECT 23.660 24.810 23.830 24.980 ;
        RECT 25.460 24.760 25.630 24.930 ;
        RECT 25.820 24.760 25.990 24.930 ;
        RECT 26.260 24.760 26.430 24.930 ;
        RECT 27.000 24.810 27.170 24.980 ;
        RECT 27.360 24.810 27.530 24.980 ;
        RECT 27.720 24.810 27.890 24.980 ;
        RECT 28.080 24.810 28.250 24.980 ;
        RECT 28.440 24.810 28.610 24.980 ;
        RECT 29.780 24.760 29.950 24.930 ;
        RECT 30.140 24.760 30.310 24.930 ;
        RECT 30.580 24.760 30.750 24.930 ;
        RECT 31.310 24.810 31.480 24.980 ;
        RECT 31.670 24.810 31.840 24.980 ;
        RECT 32.030 24.810 32.200 24.980 ;
        RECT 32.750 24.810 32.920 24.980 ;
        RECT 33.110 24.810 33.280 24.980 ;
        RECT 33.470 24.810 33.640 24.980 ;
        RECT 33.830 24.810 34.000 24.980 ;
        RECT 35.270 24.760 35.440 24.930 ;
        RECT 35.710 24.760 35.880 24.930 ;
        RECT 36.120 24.760 36.290 24.930 ;
        RECT 36.550 24.760 36.720 24.930 ;
        RECT 36.990 24.760 37.160 24.930 ;
        RECT 37.400 24.760 37.570 24.930 ;
        RECT 39.480 24.810 39.650 24.980 ;
        RECT 39.840 24.810 40.010 24.980 ;
        RECT 40.200 24.810 40.370 24.980 ;
        RECT 40.560 24.810 40.730 24.980 ;
        RECT 40.920 24.810 41.090 24.980 ;
        RECT 43.220 24.760 43.390 24.930 ;
        RECT 43.580 24.760 43.750 24.930 ;
        RECT 44.020 24.760 44.190 24.930 ;
        RECT 46.310 24.810 46.480 24.980 ;
        RECT 46.670 24.810 46.840 24.980 ;
        RECT 47.030 24.810 47.200 24.980 ;
        RECT 47.390 24.810 47.560 24.980 ;
        RECT 47.750 24.810 47.920 24.980 ;
        RECT 49.190 24.760 49.360 24.930 ;
        RECT 49.630 24.760 49.800 24.930 ;
        RECT 50.040 24.760 50.210 24.930 ;
        RECT 50.470 24.760 50.640 24.930 ;
        RECT 50.910 24.760 51.080 24.930 ;
        RECT 51.320 24.760 51.490 24.930 ;
        RECT 52.920 24.810 53.090 24.980 ;
        RECT 53.280 24.810 53.450 24.980 ;
        RECT 53.640 24.810 53.810 24.980 ;
        RECT 54.480 24.810 54.650 24.980 ;
        RECT 54.840 24.810 55.010 24.980 ;
        RECT 55.200 24.810 55.370 24.980 ;
        RECT 56.120 24.810 56.290 24.980 ;
        RECT 56.480 24.810 56.650 24.980 ;
        RECT 56.840 24.810 57.010 24.980 ;
        RECT 58.100 24.760 58.270 24.930 ;
        RECT 58.460 24.760 58.630 24.930 ;
        RECT 58.900 24.760 59.070 24.930 ;
        RECT 59.640 24.810 59.810 24.980 ;
        RECT 60.000 24.810 60.170 24.980 ;
        RECT 60.360 24.810 60.530 24.980 ;
        RECT 61.200 24.810 61.370 24.980 ;
        RECT 61.560 24.810 61.730 24.980 ;
        RECT 61.920 24.810 62.090 24.980 ;
        RECT 62.840 24.810 63.010 24.980 ;
        RECT 63.200 24.810 63.370 24.980 ;
        RECT 63.560 24.810 63.730 24.980 ;
        RECT 64.820 24.760 64.990 24.930 ;
        RECT 65.180 24.760 65.350 24.930 ;
        RECT 65.620 24.760 65.790 24.930 ;
        RECT 66.360 24.810 66.530 24.980 ;
        RECT 66.720 24.810 66.890 24.980 ;
        RECT 67.080 24.810 67.250 24.980 ;
        RECT 67.920 24.810 68.090 24.980 ;
        RECT 68.280 24.810 68.450 24.980 ;
        RECT 68.640 24.810 68.810 24.980 ;
        RECT 69.560 24.810 69.730 24.980 ;
        RECT 69.920 24.810 70.090 24.980 ;
        RECT 70.280 24.810 70.450 24.980 ;
        RECT 71.540 24.760 71.710 24.930 ;
        RECT 71.900 24.760 72.070 24.930 ;
        RECT 72.340 24.760 72.510 24.930 ;
        RECT 73.080 24.810 73.250 24.980 ;
        RECT 73.440 24.810 73.610 24.980 ;
        RECT 73.800 24.810 73.970 24.980 ;
        RECT 74.640 24.810 74.810 24.980 ;
        RECT 75.000 24.810 75.170 24.980 ;
        RECT 75.360 24.810 75.530 24.980 ;
        RECT 76.280 24.810 76.450 24.980 ;
        RECT 76.640 24.810 76.810 24.980 ;
        RECT 77.000 24.810 77.170 24.980 ;
        RECT 78.470 24.760 78.640 24.930 ;
        RECT 78.910 24.760 79.080 24.930 ;
        RECT 79.320 24.760 79.490 24.930 ;
        RECT 79.750 24.760 79.920 24.930 ;
        RECT 80.190 24.760 80.360 24.930 ;
        RECT 80.600 24.760 80.770 24.930 ;
        RECT 82.820 24.810 82.990 24.980 ;
        RECT 83.180 24.810 83.350 24.980 ;
        RECT 85.190 24.760 85.360 24.930 ;
        RECT 85.630 24.760 85.800 24.930 ;
        RECT 86.040 24.760 86.210 24.930 ;
        RECT 86.470 24.760 86.640 24.930 ;
        RECT 86.910 24.760 87.080 24.930 ;
        RECT 87.320 24.760 87.490 24.930 ;
        RECT 88.920 24.810 89.090 24.980 ;
        RECT 89.280 24.810 89.450 24.980 ;
        RECT 89.640 24.810 89.810 24.980 ;
        RECT 90.000 24.810 90.170 24.980 ;
        RECT 90.360 24.810 90.530 24.980 ;
        RECT 91.700 24.760 91.870 24.930 ;
        RECT 92.060 24.760 92.230 24.930 ;
        RECT 92.500 24.760 92.670 24.930 ;
        RECT 94.680 24.810 94.850 24.980 ;
        RECT 95.040 24.810 95.210 24.980 ;
        RECT 95.400 24.810 95.570 24.980 ;
        RECT 96.250 24.810 96.420 24.980 ;
        RECT 96.610 24.810 96.780 24.980 ;
        RECT 97.460 24.760 97.630 24.930 ;
        RECT 97.820 24.760 97.990 24.930 ;
        RECT 98.260 24.760 98.430 24.930 ;
        RECT 99.000 24.810 99.170 24.980 ;
        RECT 99.360 24.810 99.530 24.980 ;
        RECT 100.820 24.760 100.990 24.930 ;
        RECT 101.180 24.760 101.350 24.930 ;
        RECT 101.620 24.760 101.790 24.930 ;
        RECT 102.980 24.810 103.150 24.980 ;
        RECT 103.340 24.810 103.510 24.980 ;
        RECT 105.140 24.760 105.310 24.930 ;
        RECT 105.500 24.760 105.670 24.930 ;
        RECT 105.940 24.760 106.110 24.930 ;
        RECT 107.300 24.810 107.470 24.980 ;
        RECT 107.660 24.810 107.830 24.980 ;
        RECT 109.460 24.760 109.630 24.930 ;
        RECT 109.820 24.760 109.990 24.930 ;
        RECT 110.260 24.760 110.430 24.930 ;
        RECT 111.000 24.810 111.170 24.980 ;
        RECT 111.360 24.810 111.530 24.980 ;
        RECT 111.720 24.810 111.890 24.980 ;
        RECT 112.570 24.810 112.740 24.980 ;
        RECT 112.930 24.810 113.100 24.980 ;
        RECT 113.780 24.760 113.950 24.930 ;
        RECT 114.140 24.760 114.310 24.930 ;
        RECT 114.580 24.760 114.750 24.930 ;
        RECT 115.320 24.810 115.490 24.980 ;
        RECT 115.680 24.810 115.850 24.980 ;
        RECT 116.040 24.810 116.210 24.980 ;
        RECT 116.400 24.810 116.570 24.980 ;
        RECT 116.760 24.810 116.930 24.980 ;
        RECT 119.060 24.760 119.230 24.930 ;
        RECT 119.420 24.760 119.590 24.930 ;
        RECT 119.860 24.760 120.030 24.930 ;
        RECT 121.170 24.810 121.340 24.980 ;
        RECT 121.530 24.810 121.700 24.980 ;
        RECT 121.890 24.810 122.060 24.980 ;
        RECT 122.250 24.810 122.420 24.980 ;
        RECT 124.340 24.760 124.510 24.930 ;
        RECT 124.700 24.760 124.870 24.930 ;
        RECT 125.140 24.760 125.310 24.930 ;
        RECT 125.880 24.810 126.050 24.980 ;
        RECT 126.240 24.810 126.410 24.980 ;
        RECT 127.700 24.760 127.870 24.930 ;
        RECT 128.060 24.760 128.230 24.930 ;
        RECT 128.500 24.760 128.670 24.930 ;
        RECT 129.860 24.810 130.030 24.980 ;
        RECT 130.220 24.810 130.390 24.980 ;
        RECT 132.020 24.760 132.190 24.930 ;
        RECT 132.380 24.760 132.550 24.930 ;
        RECT 132.820 24.760 132.990 24.930 ;
        RECT 134.680 24.810 134.850 24.980 ;
        RECT 135.040 24.810 135.210 24.980 ;
        RECT 137.510 24.760 137.680 24.930 ;
        RECT 137.950 24.760 138.120 24.930 ;
        RECT 138.360 24.760 138.530 24.930 ;
        RECT 138.790 24.760 138.960 24.930 ;
        RECT 139.230 24.760 139.400 24.930 ;
        RECT 139.640 24.760 139.810 24.930 ;
        RECT 5.920 24.330 6.090 24.510 ;
        RECT 6.400 24.330 6.570 24.510 ;
        RECT 6.880 24.330 7.050 24.510 ;
        RECT 7.360 24.330 7.530 24.510 ;
        RECT 7.840 24.330 8.010 24.510 ;
        RECT 8.320 24.330 8.490 24.510 ;
        RECT 8.800 24.330 8.970 24.510 ;
        RECT 9.280 24.330 9.450 24.510 ;
        RECT 9.760 24.330 9.930 24.510 ;
        RECT 10.240 24.330 10.410 24.510 ;
        RECT 10.720 24.330 10.890 24.510 ;
        RECT 11.200 24.330 11.370 24.510 ;
        RECT 11.680 24.330 11.850 24.510 ;
        RECT 12.160 24.330 12.330 24.510 ;
        RECT 12.640 24.330 12.810 24.510 ;
        RECT 13.120 24.330 13.290 24.510 ;
        RECT 13.600 24.330 13.770 24.510 ;
        RECT 14.080 24.330 14.250 24.510 ;
        RECT 14.560 24.500 14.730 24.510 ;
      LAYER li1 ;
        RECT 14.400 24.330 14.880 24.500 ;
      LAYER li1 ;
        RECT 15.040 24.330 15.210 24.510 ;
        RECT 15.520 24.330 15.690 24.510 ;
        RECT 16.000 24.330 16.170 24.510 ;
        RECT 16.480 24.330 16.650 24.510 ;
      LAYER li1 ;
        RECT 16.800 24.500 17.280 24.510 ;
      LAYER li1 ;
        RECT 16.960 24.330 17.130 24.500 ;
        RECT 17.440 24.330 17.610 24.510 ;
        RECT 17.920 24.330 18.090 24.510 ;
        RECT 18.400 24.330 18.570 24.510 ;
        RECT 18.880 24.330 19.050 24.510 ;
        RECT 19.360 24.330 19.530 24.510 ;
        RECT 19.840 24.330 20.010 24.510 ;
        RECT 20.320 24.330 20.490 24.510 ;
        RECT 20.800 24.330 20.970 24.510 ;
        RECT 21.280 24.330 21.450 24.510 ;
        RECT 21.760 24.330 21.930 24.510 ;
        RECT 22.240 24.330 22.410 24.510 ;
        RECT 22.720 24.330 22.890 24.510 ;
        RECT 23.200 24.330 23.370 24.510 ;
        RECT 23.680 24.330 23.850 24.510 ;
        RECT 24.160 24.330 24.330 24.510 ;
        RECT 24.640 24.330 24.810 24.510 ;
        RECT 25.120 24.330 25.290 24.510 ;
        RECT 25.600 24.330 25.770 24.510 ;
        RECT 26.080 24.330 26.250 24.510 ;
        RECT 26.560 24.330 26.730 24.510 ;
        RECT 27.040 24.330 27.210 24.510 ;
        RECT 27.520 24.330 27.690 24.510 ;
        RECT 28.000 24.330 28.170 24.510 ;
        RECT 28.480 24.330 28.650 24.510 ;
        RECT 28.960 24.330 29.130 24.510 ;
        RECT 29.440 24.330 29.610 24.510 ;
        RECT 29.920 24.330 30.090 24.510 ;
        RECT 30.400 24.330 30.570 24.510 ;
        RECT 30.880 24.330 31.050 24.510 ;
        RECT 31.360 24.330 31.530 24.510 ;
        RECT 31.840 24.330 32.010 24.510 ;
        RECT 32.320 24.330 32.490 24.510 ;
        RECT 32.800 24.330 32.970 24.510 ;
        RECT 33.280 24.330 33.450 24.510 ;
        RECT 33.760 24.330 33.930 24.510 ;
        RECT 34.240 24.330 34.410 24.510 ;
        RECT 34.720 24.330 34.890 24.510 ;
        RECT 35.200 24.330 35.370 24.510 ;
        RECT 35.680 24.330 35.850 24.510 ;
        RECT 36.160 24.330 36.330 24.510 ;
        RECT 36.640 24.330 36.810 24.510 ;
        RECT 37.120 24.330 37.290 24.510 ;
        RECT 37.600 24.330 37.770 24.510 ;
        RECT 38.080 24.330 38.250 24.510 ;
        RECT 38.560 24.330 38.730 24.510 ;
        RECT 39.040 24.330 39.210 24.510 ;
        RECT 39.520 24.330 39.690 24.510 ;
        RECT 40.000 24.330 40.170 24.510 ;
        RECT 40.480 24.330 40.650 24.510 ;
        RECT 40.960 24.330 41.130 24.510 ;
        RECT 41.440 24.330 41.610 24.510 ;
        RECT 41.920 24.330 42.090 24.510 ;
        RECT 42.400 24.330 42.570 24.510 ;
        RECT 42.880 24.330 43.050 24.510 ;
        RECT 43.360 24.330 43.530 24.510 ;
        RECT 43.840 24.330 44.010 24.510 ;
        RECT 44.320 24.330 44.490 24.510 ;
        RECT 44.800 24.330 44.970 24.510 ;
        RECT 45.280 24.330 45.450 24.510 ;
        RECT 45.760 24.330 45.930 24.510 ;
        RECT 46.240 24.330 46.410 24.510 ;
        RECT 46.720 24.330 46.890 24.510 ;
        RECT 47.200 24.330 47.370 24.510 ;
        RECT 47.680 24.330 47.850 24.510 ;
        RECT 48.160 24.330 48.330 24.510 ;
        RECT 48.640 24.330 48.810 24.510 ;
        RECT 49.120 24.330 49.290 24.510 ;
        RECT 49.600 24.330 49.770 24.510 ;
        RECT 50.080 24.330 50.250 24.510 ;
        RECT 50.560 24.330 50.730 24.510 ;
        RECT 51.040 24.330 51.210 24.510 ;
        RECT 51.520 24.330 51.690 24.510 ;
        RECT 52.000 24.330 52.170 24.510 ;
        RECT 52.480 24.500 52.650 24.510 ;
      LAYER li1 ;
        RECT 52.320 24.330 52.800 24.500 ;
      LAYER li1 ;
        RECT 52.960 24.330 53.130 24.510 ;
        RECT 53.440 24.330 53.610 24.510 ;
        RECT 53.920 24.330 54.090 24.510 ;
        RECT 54.400 24.330 54.570 24.510 ;
        RECT 54.880 24.330 55.050 24.510 ;
        RECT 55.360 24.330 55.530 24.510 ;
        RECT 55.840 24.330 56.010 24.510 ;
        RECT 56.320 24.330 56.490 24.510 ;
        RECT 56.800 24.330 56.970 24.510 ;
        RECT 57.280 24.330 57.450 24.510 ;
        RECT 57.760 24.330 57.930 24.510 ;
        RECT 58.240 24.330 58.410 24.510 ;
        RECT 58.720 24.330 58.890 24.510 ;
        RECT 59.200 24.330 59.370 24.510 ;
        RECT 59.680 24.330 59.850 24.510 ;
        RECT 60.160 24.330 60.330 24.510 ;
        RECT 60.640 24.330 60.810 24.510 ;
        RECT 61.120 24.330 61.290 24.510 ;
        RECT 61.600 24.330 61.770 24.510 ;
        RECT 62.080 24.330 62.250 24.510 ;
        RECT 62.560 24.330 62.730 24.510 ;
        RECT 63.040 24.330 63.210 24.510 ;
        RECT 63.520 24.330 63.690 24.510 ;
        RECT 64.000 24.330 64.170 24.510 ;
        RECT 64.480 24.330 64.650 24.510 ;
        RECT 64.960 24.330 65.130 24.510 ;
        RECT 65.440 24.330 65.610 24.510 ;
        RECT 65.920 24.330 66.090 24.510 ;
        RECT 66.400 24.330 66.570 24.510 ;
        RECT 66.880 24.330 67.050 24.510 ;
        RECT 67.360 24.330 67.530 24.510 ;
        RECT 67.840 24.330 68.010 24.510 ;
        RECT 68.320 24.330 68.490 24.510 ;
        RECT 68.800 24.330 68.970 24.510 ;
        RECT 69.280 24.330 69.450 24.510 ;
        RECT 69.760 24.330 69.930 24.510 ;
        RECT 70.240 24.330 70.410 24.510 ;
        RECT 70.720 24.330 70.890 24.510 ;
        RECT 71.200 24.330 71.370 24.510 ;
        RECT 71.680 24.330 71.850 24.510 ;
        RECT 72.160 24.330 72.330 24.510 ;
        RECT 72.640 24.330 72.810 24.510 ;
        RECT 73.120 24.330 73.290 24.510 ;
        RECT 73.600 24.330 73.770 24.510 ;
        RECT 74.080 24.330 74.250 24.510 ;
        RECT 74.560 24.330 74.730 24.510 ;
        RECT 75.040 24.330 75.210 24.510 ;
        RECT 75.520 24.330 75.690 24.510 ;
        RECT 76.000 24.330 76.170 24.510 ;
        RECT 76.480 24.330 76.650 24.510 ;
        RECT 76.960 24.330 77.130 24.510 ;
        RECT 77.440 24.330 77.610 24.510 ;
        RECT 77.920 24.330 78.090 24.510 ;
        RECT 78.400 24.330 78.570 24.510 ;
        RECT 78.880 24.330 79.050 24.510 ;
        RECT 79.360 24.330 79.530 24.510 ;
        RECT 79.840 24.330 80.010 24.510 ;
        RECT 80.320 24.330 80.490 24.510 ;
        RECT 80.800 24.330 80.970 24.510 ;
        RECT 81.280 24.330 81.450 24.510 ;
        RECT 81.760 24.500 81.930 24.510 ;
      LAYER li1 ;
        RECT 81.600 24.330 82.080 24.500 ;
      LAYER li1 ;
        RECT 82.240 24.330 82.410 24.510 ;
        RECT 82.720 24.330 82.890 24.510 ;
        RECT 83.200 24.330 83.370 24.510 ;
        RECT 83.680 24.330 83.850 24.510 ;
        RECT 84.160 24.330 84.330 24.510 ;
        RECT 84.640 24.330 84.810 24.510 ;
        RECT 85.120 24.330 85.290 24.510 ;
        RECT 85.600 24.330 85.770 24.510 ;
        RECT 86.080 24.330 86.250 24.510 ;
        RECT 86.560 24.330 86.730 24.510 ;
        RECT 87.040 24.330 87.210 24.510 ;
        RECT 87.520 24.330 87.690 24.510 ;
        RECT 88.000 24.330 88.170 24.510 ;
        RECT 88.480 24.500 88.650 24.510 ;
      LAYER li1 ;
        RECT 88.320 24.330 88.800 24.500 ;
      LAYER li1 ;
        RECT 88.960 24.330 89.130 24.510 ;
        RECT 89.440 24.330 89.610 24.510 ;
        RECT 89.920 24.330 90.090 24.510 ;
        RECT 90.400 24.330 90.570 24.510 ;
        RECT 90.880 24.330 91.050 24.510 ;
        RECT 91.360 24.330 91.530 24.510 ;
        RECT 91.840 24.330 92.010 24.510 ;
        RECT 92.320 24.330 92.490 24.510 ;
        RECT 92.800 24.330 92.970 24.510 ;
        RECT 93.280 24.330 93.450 24.510 ;
        RECT 93.760 24.330 93.930 24.510 ;
        RECT 94.240 24.500 94.410 24.510 ;
      LAYER li1 ;
        RECT 94.080 24.330 94.560 24.500 ;
      LAYER li1 ;
        RECT 94.720 24.330 94.890 24.510 ;
        RECT 95.200 24.330 95.370 24.510 ;
        RECT 95.680 24.330 95.850 24.510 ;
        RECT 96.160 24.330 96.330 24.510 ;
        RECT 96.640 24.330 96.810 24.510 ;
        RECT 97.120 24.330 97.290 24.510 ;
        RECT 97.600 24.330 97.770 24.510 ;
        RECT 98.080 24.330 98.250 24.510 ;
        RECT 98.560 24.330 98.730 24.510 ;
        RECT 99.040 24.330 99.210 24.510 ;
        RECT 99.520 24.330 99.690 24.510 ;
        RECT 100.000 24.330 100.170 24.510 ;
        RECT 100.480 24.330 100.650 24.510 ;
        RECT 100.960 24.330 101.130 24.510 ;
        RECT 101.440 24.330 101.610 24.510 ;
        RECT 101.920 24.330 102.090 24.510 ;
        RECT 102.400 24.330 102.570 24.510 ;
        RECT 102.880 24.330 103.050 24.510 ;
        RECT 103.360 24.330 103.530 24.510 ;
        RECT 103.840 24.330 104.010 24.510 ;
        RECT 104.320 24.330 104.490 24.510 ;
        RECT 104.800 24.330 104.970 24.510 ;
        RECT 105.280 24.330 105.450 24.510 ;
        RECT 105.760 24.330 105.930 24.510 ;
        RECT 106.240 24.330 106.410 24.510 ;
        RECT 106.720 24.330 106.890 24.510 ;
        RECT 107.200 24.330 107.370 24.510 ;
        RECT 107.680 24.330 107.850 24.510 ;
        RECT 108.160 24.330 108.330 24.510 ;
        RECT 108.640 24.330 108.810 24.510 ;
        RECT 109.120 24.330 109.290 24.510 ;
        RECT 109.600 24.330 109.770 24.510 ;
        RECT 110.080 24.330 110.250 24.510 ;
        RECT 110.560 24.330 110.730 24.510 ;
        RECT 111.040 24.330 111.210 24.510 ;
        RECT 111.520 24.330 111.690 24.510 ;
        RECT 112.000 24.330 112.170 24.510 ;
        RECT 112.480 24.330 112.650 24.510 ;
        RECT 112.960 24.330 113.130 24.510 ;
        RECT 113.440 24.330 113.610 24.510 ;
        RECT 113.920 24.330 114.090 24.510 ;
        RECT 114.400 24.330 114.570 24.510 ;
        RECT 114.880 24.330 115.050 24.510 ;
        RECT 115.360 24.330 115.530 24.510 ;
        RECT 115.840 24.330 116.010 24.510 ;
        RECT 116.320 24.330 116.490 24.510 ;
        RECT 116.800 24.330 116.970 24.510 ;
        RECT 117.280 24.330 117.450 24.510 ;
        RECT 117.760 24.330 117.930 24.510 ;
        RECT 118.240 24.330 118.410 24.510 ;
        RECT 118.720 24.330 118.890 24.510 ;
        RECT 119.200 24.330 119.370 24.510 ;
        RECT 119.680 24.330 119.850 24.510 ;
        RECT 120.160 24.330 120.330 24.510 ;
        RECT 120.640 24.330 120.810 24.510 ;
        RECT 121.120 24.330 121.290 24.510 ;
        RECT 121.600 24.330 121.770 24.510 ;
        RECT 122.080 24.330 122.250 24.510 ;
        RECT 122.560 24.330 122.730 24.510 ;
        RECT 123.040 24.330 123.210 24.510 ;
        RECT 123.520 24.330 123.690 24.510 ;
        RECT 124.000 24.330 124.170 24.510 ;
        RECT 124.480 24.330 124.650 24.510 ;
        RECT 124.960 24.330 125.130 24.510 ;
        RECT 125.440 24.330 125.610 24.510 ;
        RECT 125.920 24.330 126.090 24.510 ;
        RECT 126.400 24.330 126.570 24.510 ;
        RECT 126.880 24.330 127.050 24.510 ;
        RECT 127.360 24.330 127.530 24.510 ;
        RECT 127.840 24.330 128.010 24.510 ;
        RECT 128.320 24.330 128.490 24.510 ;
        RECT 128.800 24.330 128.970 24.510 ;
        RECT 129.280 24.330 129.450 24.510 ;
        RECT 129.760 24.330 129.930 24.510 ;
        RECT 130.240 24.330 130.410 24.510 ;
        RECT 130.720 24.330 130.890 24.510 ;
        RECT 131.200 24.330 131.370 24.510 ;
        RECT 131.680 24.330 131.850 24.510 ;
        RECT 132.160 24.330 132.330 24.510 ;
        RECT 132.640 24.330 132.810 24.510 ;
        RECT 133.120 24.330 133.290 24.510 ;
        RECT 133.600 24.330 133.770 24.510 ;
        RECT 134.080 24.330 134.250 24.510 ;
        RECT 134.560 24.330 134.730 24.510 ;
        RECT 135.040 24.330 135.210 24.510 ;
        RECT 135.520 24.330 135.690 24.510 ;
        RECT 136.000 24.330 136.170 24.510 ;
        RECT 136.480 24.330 136.650 24.510 ;
        RECT 136.960 24.330 137.130 24.510 ;
        RECT 137.440 24.330 137.610 24.510 ;
        RECT 137.920 24.330 138.090 24.510 ;
        RECT 138.400 24.330 138.570 24.510 ;
        RECT 138.880 24.330 139.050 24.510 ;
        RECT 139.360 24.330 139.530 24.510 ;
        RECT 139.840 24.330 140.010 24.510 ;
        RECT 140.320 24.330 140.490 24.510 ;
        RECT 140.800 24.330 140.970 24.510 ;
        RECT 141.280 24.330 141.450 24.510 ;
        RECT 141.760 24.500 141.930 24.510 ;
      LAYER li1 ;
        RECT 141.600 24.330 142.080 24.500 ;
      LAYER li1 ;
        RECT 6.470 23.910 6.640 24.080 ;
        RECT 6.910 23.910 7.080 24.080 ;
        RECT 7.320 23.910 7.490 24.080 ;
        RECT 7.750 23.910 7.920 24.080 ;
        RECT 8.190 23.910 8.360 24.080 ;
        RECT 8.600 23.910 8.770 24.080 ;
        RECT 10.840 23.860 11.010 24.030 ;
        RECT 11.200 23.860 11.370 24.030 ;
        RECT 13.670 23.910 13.840 24.080 ;
        RECT 14.110 23.910 14.280 24.080 ;
        RECT 14.520 23.910 14.690 24.080 ;
        RECT 14.950 23.910 15.120 24.080 ;
        RECT 15.390 23.910 15.560 24.080 ;
        RECT 15.800 23.910 15.970 24.080 ;
        RECT 17.560 23.860 17.730 24.030 ;
        RECT 17.920 23.860 18.090 24.030 ;
        RECT 20.180 23.910 20.350 24.080 ;
        RECT 20.540 23.910 20.710 24.080 ;
        RECT 20.980 23.910 21.150 24.080 ;
        RECT 21.880 23.860 22.050 24.030 ;
        RECT 22.240 23.860 22.410 24.030 ;
        RECT 24.500 23.910 24.670 24.080 ;
        RECT 24.860 23.910 25.030 24.080 ;
        RECT 25.300 23.910 25.470 24.080 ;
        RECT 26.580 23.860 26.750 24.030 ;
        RECT 26.940 23.860 27.110 24.030 ;
        RECT 28.970 23.860 29.140 24.030 ;
        RECT 31.400 23.860 31.570 24.030 ;
        RECT 31.760 23.860 31.930 24.030 ;
        RECT 32.120 23.860 32.290 24.030 ;
        RECT 33.740 23.860 33.910 24.030 ;
        RECT 34.100 23.860 34.270 24.030 ;
        RECT 34.460 23.860 34.630 24.030 ;
        RECT 36.440 23.860 36.610 24.030 ;
        RECT 36.800 23.860 36.970 24.030 ;
        RECT 37.160 23.860 37.330 24.030 ;
        RECT 38.190 23.860 38.360 24.030 ;
        RECT 38.550 23.860 38.720 24.030 ;
        RECT 38.910 23.860 39.080 24.030 ;
        RECT 39.720 23.860 39.890 24.030 ;
        RECT 40.080 23.860 40.250 24.030 ;
        RECT 40.440 23.860 40.610 24.030 ;
        RECT 41.990 23.910 42.160 24.080 ;
        RECT 42.430 23.910 42.600 24.080 ;
        RECT 42.840 23.910 43.010 24.080 ;
        RECT 43.270 23.910 43.440 24.080 ;
        RECT 43.710 23.910 43.880 24.080 ;
        RECT 44.120 23.910 44.290 24.080 ;
        RECT 45.700 23.860 45.870 24.030 ;
        RECT 46.060 23.860 46.230 24.030 ;
        RECT 46.420 23.860 46.590 24.030 ;
        RECT 47.390 23.860 47.560 24.030 ;
        RECT 50.760 23.860 50.930 24.030 ;
        RECT 52.230 23.860 52.400 24.030 ;
        RECT 52.590 23.860 52.760 24.030 ;
        RECT 52.950 23.860 53.120 24.030 ;
        RECT 55.160 23.860 55.330 24.030 ;
        RECT 55.520 23.860 55.690 24.030 ;
        RECT 55.880 23.860 56.050 24.030 ;
        RECT 56.880 23.860 57.050 24.030 ;
        RECT 57.240 23.860 57.410 24.030 ;
        RECT 57.600 23.860 57.770 24.030 ;
        RECT 58.440 23.860 58.610 24.030 ;
        RECT 58.800 23.860 58.970 24.030 ;
        RECT 59.160 23.860 59.330 24.030 ;
        RECT 60.710 23.910 60.880 24.080 ;
        RECT 61.150 23.910 61.320 24.080 ;
        RECT 61.560 23.910 61.730 24.080 ;
        RECT 61.990 23.910 62.160 24.080 ;
        RECT 62.430 23.910 62.600 24.080 ;
        RECT 62.840 23.910 63.010 24.080 ;
        RECT 64.500 23.860 64.670 24.030 ;
        RECT 64.860 23.860 65.030 24.030 ;
        RECT 66.890 23.860 67.060 24.030 ;
        RECT 69.320 23.860 69.490 24.030 ;
        RECT 69.680 23.860 69.850 24.030 ;
        RECT 70.040 23.860 70.210 24.030 ;
        RECT 71.660 23.860 71.830 24.030 ;
        RECT 72.020 23.860 72.190 24.030 ;
        RECT 72.380 23.860 72.550 24.030 ;
        RECT 74.360 23.860 74.530 24.030 ;
        RECT 74.720 23.860 74.890 24.030 ;
        RECT 75.080 23.860 75.250 24.030 ;
        RECT 76.110 23.860 76.280 24.030 ;
        RECT 76.470 23.860 76.640 24.030 ;
        RECT 76.830 23.860 77.000 24.030 ;
        RECT 77.640 23.860 77.810 24.030 ;
        RECT 78.000 23.860 78.170 24.030 ;
        RECT 78.360 23.860 78.530 24.030 ;
        RECT 79.700 23.910 79.870 24.080 ;
        RECT 80.060 23.910 80.230 24.080 ;
        RECT 80.500 23.910 80.670 24.080 ;
        RECT 81.860 23.860 82.030 24.030 ;
        RECT 82.220 23.860 82.390 24.030 ;
        RECT 84.020 23.910 84.190 24.080 ;
        RECT 84.380 23.910 84.550 24.080 ;
        RECT 84.820 23.910 84.990 24.080 ;
        RECT 86.180 23.860 86.350 24.030 ;
        RECT 86.540 23.860 86.710 24.030 ;
        RECT 88.340 23.910 88.510 24.080 ;
        RECT 88.700 23.910 88.870 24.080 ;
        RECT 89.140 23.910 89.310 24.080 ;
        RECT 90.840 23.860 91.010 24.030 ;
        RECT 91.200 23.860 91.370 24.030 ;
        RECT 91.560 23.860 91.730 24.030 ;
        RECT 91.920 23.860 92.090 24.030 ;
        RECT 92.280 23.860 92.450 24.030 ;
        RECT 93.620 23.910 93.790 24.080 ;
        RECT 93.980 23.910 94.150 24.080 ;
        RECT 94.420 23.910 94.590 24.080 ;
        RECT 95.780 23.860 95.950 24.030 ;
        RECT 96.140 23.860 96.310 24.030 ;
        RECT 97.940 23.910 98.110 24.080 ;
        RECT 98.300 23.910 98.470 24.080 ;
        RECT 98.740 23.910 98.910 24.080 ;
        RECT 99.480 23.860 99.650 24.030 ;
        RECT 99.840 23.860 100.010 24.030 ;
        RECT 100.200 23.860 100.370 24.030 ;
        RECT 101.050 23.860 101.220 24.030 ;
        RECT 101.410 23.860 101.580 24.030 ;
        RECT 102.260 23.910 102.430 24.080 ;
        RECT 102.620 23.910 102.790 24.080 ;
        RECT 103.060 23.910 103.230 24.080 ;
        RECT 103.800 23.860 103.970 24.030 ;
        RECT 104.160 23.860 104.330 24.030 ;
        RECT 104.520 23.860 104.690 24.030 ;
        RECT 105.370 23.860 105.540 24.030 ;
        RECT 105.730 23.860 105.900 24.030 ;
        RECT 106.580 23.910 106.750 24.080 ;
        RECT 106.940 23.910 107.110 24.080 ;
        RECT 107.380 23.910 107.550 24.080 ;
        RECT 109.700 23.860 109.870 24.030 ;
        RECT 110.060 23.860 110.230 24.030 ;
        RECT 111.860 23.910 112.030 24.080 ;
        RECT 112.220 23.910 112.390 24.080 ;
        RECT 112.660 23.910 112.830 24.080 ;
        RECT 113.400 23.860 113.570 24.030 ;
        RECT 113.760 23.860 113.930 24.030 ;
        RECT 114.120 23.860 114.290 24.030 ;
        RECT 114.480 23.860 114.650 24.030 ;
        RECT 114.840 23.860 115.010 24.030 ;
        RECT 116.180 23.910 116.350 24.080 ;
        RECT 116.540 23.910 116.710 24.080 ;
        RECT 116.980 23.910 117.150 24.080 ;
        RECT 117.720 23.860 117.890 24.030 ;
        RECT 118.080 23.860 118.250 24.030 ;
        RECT 118.440 23.860 118.610 24.030 ;
        RECT 118.800 23.860 118.970 24.030 ;
        RECT 119.160 23.860 119.330 24.030 ;
        RECT 120.500 23.910 120.670 24.080 ;
        RECT 120.860 23.910 121.030 24.080 ;
        RECT 121.300 23.910 121.470 24.080 ;
        RECT 122.580 23.860 122.750 24.030 ;
        RECT 122.940 23.860 123.110 24.030 ;
        RECT 124.970 23.860 125.140 24.030 ;
        RECT 127.400 23.860 127.570 24.030 ;
        RECT 127.760 23.860 127.930 24.030 ;
        RECT 128.120 23.860 128.290 24.030 ;
        RECT 129.740 23.860 129.910 24.030 ;
        RECT 130.100 23.860 130.270 24.030 ;
        RECT 130.460 23.860 130.630 24.030 ;
        RECT 132.440 23.860 132.610 24.030 ;
        RECT 132.800 23.860 132.970 24.030 ;
        RECT 133.160 23.860 133.330 24.030 ;
        RECT 134.190 23.860 134.360 24.030 ;
        RECT 134.550 23.860 134.720 24.030 ;
        RECT 134.910 23.860 135.080 24.030 ;
        RECT 135.720 23.860 135.890 24.030 ;
        RECT 136.080 23.860 136.250 24.030 ;
        RECT 136.440 23.860 136.610 24.030 ;
        RECT 137.990 23.910 138.160 24.080 ;
        RECT 138.430 23.910 138.600 24.080 ;
        RECT 138.840 23.910 139.010 24.080 ;
        RECT 139.270 23.910 139.440 24.080 ;
        RECT 139.710 23.910 139.880 24.080 ;
        RECT 140.120 23.910 140.290 24.080 ;
        RECT 6.470 16.620 6.640 16.790 ;
        RECT 6.910 16.620 7.080 16.790 ;
        RECT 7.320 16.620 7.490 16.790 ;
        RECT 7.750 16.620 7.920 16.790 ;
        RECT 8.190 16.620 8.360 16.790 ;
        RECT 8.600 16.620 8.770 16.790 ;
        RECT 10.100 16.620 10.270 16.790 ;
        RECT 10.460 16.620 10.630 16.790 ;
        RECT 10.900 16.620 11.070 16.790 ;
        RECT 11.800 16.670 11.970 16.840 ;
        RECT 12.160 16.670 12.330 16.840 ;
        RECT 14.420 16.620 14.590 16.790 ;
        RECT 14.780 16.620 14.950 16.790 ;
        RECT 15.220 16.620 15.390 16.790 ;
        RECT 16.120 16.670 16.290 16.840 ;
        RECT 16.480 16.670 16.650 16.840 ;
        RECT 18.740 16.620 18.910 16.790 ;
        RECT 19.100 16.620 19.270 16.790 ;
        RECT 19.540 16.620 19.710 16.790 ;
        RECT 20.440 16.670 20.610 16.840 ;
        RECT 20.800 16.670 20.970 16.840 ;
        RECT 23.060 16.620 23.230 16.790 ;
        RECT 23.420 16.620 23.590 16.790 ;
        RECT 23.860 16.620 24.030 16.790 ;
        RECT 25.220 16.670 25.390 16.840 ;
        RECT 25.580 16.670 25.750 16.840 ;
        RECT 27.380 16.620 27.550 16.790 ;
        RECT 27.740 16.620 27.910 16.790 ;
        RECT 28.180 16.620 28.350 16.790 ;
        RECT 29.540 16.670 29.710 16.840 ;
        RECT 29.900 16.670 30.070 16.840 ;
        RECT 31.700 16.620 31.870 16.790 ;
        RECT 32.060 16.620 32.230 16.790 ;
        RECT 32.500 16.620 32.670 16.790 ;
        RECT 33.860 16.670 34.030 16.840 ;
        RECT 34.220 16.670 34.390 16.840 ;
        RECT 36.020 16.620 36.190 16.790 ;
        RECT 36.380 16.620 36.550 16.790 ;
        RECT 36.820 16.620 36.990 16.790 ;
        RECT 38.040 16.670 38.210 16.840 ;
        RECT 38.400 16.670 38.570 16.840 ;
        RECT 39.860 16.620 40.030 16.790 ;
        RECT 40.220 16.620 40.390 16.790 ;
        RECT 40.660 16.620 40.830 16.790 ;
        RECT 42.020 16.670 42.190 16.840 ;
        RECT 42.380 16.670 42.550 16.840 ;
        RECT 44.180 16.620 44.350 16.790 ;
        RECT 44.540 16.620 44.710 16.790 ;
        RECT 44.980 16.620 45.150 16.790 ;
        RECT 45.720 16.670 45.890 16.840 ;
        RECT 46.080 16.670 46.250 16.840 ;
        RECT 46.440 16.670 46.610 16.840 ;
        RECT 46.800 16.670 46.970 16.840 ;
        RECT 47.160 16.670 47.330 16.840 ;
        RECT 49.460 16.620 49.630 16.790 ;
        RECT 49.820 16.620 49.990 16.790 ;
        RECT 50.260 16.620 50.430 16.790 ;
        RECT 51.000 16.670 51.170 16.840 ;
        RECT 51.360 16.670 51.530 16.840 ;
        RECT 51.720 16.670 51.890 16.840 ;
        RECT 52.080 16.670 52.250 16.840 ;
        RECT 52.440 16.670 52.610 16.840 ;
        RECT 54.740 16.620 54.910 16.790 ;
        RECT 55.100 16.620 55.270 16.790 ;
        RECT 55.540 16.620 55.710 16.790 ;
        RECT 56.280 16.670 56.450 16.840 ;
        RECT 56.640 16.670 56.810 16.840 ;
        RECT 58.100 16.620 58.270 16.790 ;
        RECT 58.460 16.620 58.630 16.790 ;
        RECT 58.900 16.620 59.070 16.790 ;
        RECT 59.640 16.670 59.810 16.840 ;
        RECT 60.000 16.670 60.170 16.840 ;
        RECT 60.360 16.670 60.530 16.840 ;
        RECT 61.200 16.670 61.370 16.840 ;
        RECT 61.560 16.670 61.730 16.840 ;
        RECT 61.920 16.670 62.090 16.840 ;
        RECT 62.840 16.670 63.010 16.840 ;
        RECT 63.200 16.670 63.370 16.840 ;
        RECT 63.560 16.670 63.730 16.840 ;
        RECT 64.820 16.620 64.990 16.790 ;
        RECT 65.180 16.620 65.350 16.790 ;
        RECT 65.620 16.620 65.790 16.790 ;
        RECT 66.340 16.670 66.510 16.840 ;
        RECT 66.700 16.670 66.870 16.840 ;
        RECT 67.060 16.670 67.230 16.840 ;
        RECT 67.420 16.670 67.590 16.840 ;
        RECT 68.580 16.670 68.750 16.840 ;
        RECT 68.940 16.670 69.110 16.840 ;
        RECT 69.300 16.670 69.470 16.840 ;
        RECT 69.660 16.670 69.830 16.840 ;
        RECT 70.580 16.620 70.750 16.790 ;
        RECT 70.940 16.620 71.110 16.790 ;
        RECT 71.380 16.620 71.550 16.790 ;
        RECT 72.740 16.670 72.910 16.840 ;
        RECT 73.100 16.670 73.270 16.840 ;
        RECT 74.900 16.620 75.070 16.790 ;
        RECT 75.260 16.620 75.430 16.790 ;
        RECT 75.700 16.620 75.870 16.790 ;
        RECT 77.060 16.670 77.230 16.840 ;
        RECT 77.420 16.670 77.590 16.840 ;
        RECT 79.430 16.620 79.600 16.790 ;
        RECT 79.870 16.620 80.040 16.790 ;
        RECT 80.280 16.620 80.450 16.790 ;
        RECT 80.710 16.620 80.880 16.790 ;
        RECT 81.150 16.620 81.320 16.790 ;
        RECT 81.560 16.620 81.730 16.790 ;
        RECT 83.220 16.670 83.390 16.840 ;
        RECT 83.580 16.670 83.750 16.840 ;
        RECT 85.610 16.670 85.780 16.840 ;
        RECT 88.040 16.670 88.210 16.840 ;
        RECT 88.400 16.670 88.570 16.840 ;
        RECT 88.760 16.670 88.930 16.840 ;
        RECT 90.380 16.670 90.550 16.840 ;
        RECT 90.740 16.670 90.910 16.840 ;
        RECT 91.100 16.670 91.270 16.840 ;
        RECT 93.080 16.670 93.250 16.840 ;
        RECT 93.440 16.670 93.610 16.840 ;
        RECT 93.800 16.670 93.970 16.840 ;
        RECT 94.830 16.670 95.000 16.840 ;
        RECT 95.190 16.670 95.360 16.840 ;
        RECT 95.550 16.670 95.720 16.840 ;
        RECT 96.360 16.670 96.530 16.840 ;
        RECT 96.720 16.670 96.890 16.840 ;
        RECT 97.080 16.670 97.250 16.840 ;
        RECT 98.630 16.620 98.800 16.790 ;
        RECT 99.070 16.620 99.240 16.790 ;
        RECT 99.480 16.620 99.650 16.790 ;
        RECT 99.910 16.620 100.080 16.790 ;
        RECT 100.350 16.620 100.520 16.790 ;
        RECT 100.760 16.620 100.930 16.790 ;
        RECT 103.380 16.670 103.550 16.840 ;
        RECT 103.740 16.670 103.910 16.840 ;
        RECT 105.770 16.670 105.940 16.840 ;
        RECT 108.200 16.670 108.370 16.840 ;
        RECT 108.560 16.670 108.730 16.840 ;
        RECT 108.920 16.670 109.090 16.840 ;
        RECT 110.540 16.670 110.710 16.840 ;
        RECT 110.900 16.670 111.070 16.840 ;
        RECT 111.260 16.670 111.430 16.840 ;
        RECT 113.240 16.670 113.410 16.840 ;
        RECT 113.600 16.670 113.770 16.840 ;
        RECT 113.960 16.670 114.130 16.840 ;
        RECT 114.990 16.670 115.160 16.840 ;
        RECT 115.350 16.670 115.520 16.840 ;
        RECT 115.710 16.670 115.880 16.840 ;
        RECT 116.520 16.670 116.690 16.840 ;
        RECT 116.880 16.670 117.050 16.840 ;
        RECT 117.240 16.670 117.410 16.840 ;
        RECT 118.580 16.620 118.750 16.790 ;
        RECT 118.940 16.620 119.110 16.790 ;
        RECT 119.380 16.620 119.550 16.790 ;
        RECT 120.280 16.670 120.450 16.840 ;
        RECT 120.640 16.670 120.810 16.840 ;
        RECT 122.900 16.620 123.070 16.790 ;
        RECT 123.260 16.620 123.430 16.790 ;
        RECT 123.700 16.620 123.870 16.790 ;
        RECT 124.600 16.670 124.770 16.840 ;
        RECT 124.960 16.670 125.130 16.840 ;
        RECT 127.430 16.620 127.600 16.790 ;
        RECT 127.870 16.620 128.040 16.790 ;
        RECT 128.280 16.620 128.450 16.790 ;
        RECT 128.710 16.620 128.880 16.790 ;
        RECT 129.150 16.620 129.320 16.790 ;
        RECT 129.560 16.620 129.730 16.790 ;
        RECT 131.270 16.620 131.440 16.790 ;
        RECT 131.710 16.620 131.880 16.790 ;
        RECT 132.120 16.620 132.290 16.790 ;
        RECT 132.550 16.620 132.720 16.790 ;
        RECT 132.990 16.620 133.160 16.790 ;
        RECT 133.400 16.620 133.570 16.790 ;
        RECT 134.680 16.670 134.850 16.840 ;
        RECT 135.040 16.670 135.210 16.840 ;
        RECT 137.510 16.620 137.680 16.790 ;
        RECT 137.950 16.620 138.120 16.790 ;
        RECT 138.360 16.620 138.530 16.790 ;
        RECT 138.790 16.620 138.960 16.790 ;
        RECT 139.230 16.620 139.400 16.790 ;
        RECT 139.640 16.620 139.810 16.790 ;
        RECT 5.920 16.190 6.090 16.360 ;
        RECT 6.400 16.190 6.570 16.360 ;
        RECT 6.880 16.190 7.050 16.360 ;
        RECT 7.360 16.190 7.530 16.360 ;
        RECT 7.840 16.190 8.010 16.360 ;
        RECT 8.320 16.190 8.490 16.360 ;
        RECT 8.800 16.190 8.970 16.360 ;
        RECT 9.280 16.190 9.450 16.360 ;
        RECT 9.760 16.190 9.930 16.360 ;
        RECT 10.240 16.190 10.410 16.360 ;
        RECT 10.720 16.190 10.890 16.360 ;
        RECT 11.200 16.190 11.370 16.360 ;
        RECT 11.680 16.190 11.850 16.360 ;
        RECT 12.160 16.190 12.330 16.360 ;
        RECT 12.640 16.190 12.810 16.360 ;
        RECT 13.120 16.190 13.290 16.360 ;
        RECT 13.600 16.190 13.770 16.360 ;
        RECT 14.080 16.190 14.250 16.360 ;
        RECT 14.560 16.190 14.730 16.360 ;
        RECT 15.040 16.190 15.210 16.360 ;
        RECT 15.520 16.190 15.690 16.360 ;
        RECT 16.000 16.190 16.170 16.360 ;
        RECT 16.480 16.190 16.650 16.360 ;
        RECT 16.960 16.190 17.130 16.360 ;
        RECT 17.440 16.190 17.610 16.360 ;
        RECT 17.920 16.190 18.090 16.360 ;
        RECT 18.400 16.190 18.570 16.360 ;
        RECT 18.880 16.190 19.050 16.360 ;
        RECT 19.360 16.190 19.530 16.360 ;
        RECT 19.840 16.190 20.010 16.360 ;
        RECT 20.320 16.190 20.490 16.360 ;
        RECT 20.800 16.190 20.970 16.360 ;
        RECT 21.280 16.190 21.450 16.360 ;
        RECT 21.760 16.190 21.930 16.360 ;
        RECT 22.240 16.190 22.410 16.360 ;
        RECT 22.720 16.190 22.890 16.360 ;
        RECT 23.200 16.190 23.370 16.360 ;
        RECT 23.680 16.190 23.850 16.360 ;
        RECT 24.160 16.190 24.330 16.360 ;
        RECT 24.640 16.190 24.810 16.360 ;
        RECT 25.120 16.190 25.290 16.360 ;
        RECT 25.600 16.190 25.770 16.360 ;
        RECT 26.080 16.190 26.250 16.360 ;
        RECT 26.560 16.190 26.730 16.360 ;
        RECT 27.040 16.190 27.210 16.360 ;
        RECT 27.520 16.190 27.690 16.360 ;
        RECT 28.000 16.190 28.170 16.360 ;
        RECT 28.480 16.190 28.650 16.360 ;
        RECT 28.960 16.190 29.130 16.360 ;
        RECT 29.440 16.190 29.610 16.360 ;
        RECT 29.920 16.190 30.090 16.360 ;
        RECT 30.400 16.190 30.570 16.360 ;
        RECT 30.880 16.190 31.050 16.360 ;
        RECT 31.360 16.190 31.530 16.360 ;
        RECT 31.840 16.190 32.010 16.360 ;
        RECT 32.320 16.190 32.490 16.360 ;
        RECT 32.800 16.190 32.970 16.360 ;
        RECT 33.280 16.190 33.450 16.360 ;
        RECT 33.760 16.190 33.930 16.360 ;
        RECT 34.240 16.190 34.410 16.360 ;
        RECT 34.720 16.190 34.890 16.360 ;
        RECT 35.200 16.190 35.370 16.360 ;
        RECT 35.680 16.190 35.850 16.360 ;
        RECT 36.160 16.190 36.330 16.360 ;
        RECT 36.640 16.190 36.810 16.360 ;
        RECT 37.120 16.190 37.290 16.360 ;
      LAYER li1 ;
        RECT 37.440 16.190 37.920 16.360 ;
      LAYER li1 ;
        RECT 38.080 16.190 38.250 16.360 ;
        RECT 38.560 16.190 38.730 16.360 ;
        RECT 39.040 16.190 39.210 16.360 ;
        RECT 39.520 16.190 39.690 16.360 ;
        RECT 40.000 16.190 40.170 16.360 ;
        RECT 40.480 16.190 40.650 16.360 ;
        RECT 40.960 16.190 41.130 16.360 ;
        RECT 41.440 16.190 41.610 16.360 ;
        RECT 41.920 16.190 42.090 16.360 ;
        RECT 42.400 16.190 42.570 16.360 ;
        RECT 42.880 16.190 43.050 16.360 ;
        RECT 43.360 16.190 43.530 16.360 ;
        RECT 43.840 16.190 44.010 16.360 ;
        RECT 44.320 16.190 44.490 16.360 ;
        RECT 44.800 16.190 44.970 16.360 ;
        RECT 45.280 16.190 45.450 16.360 ;
        RECT 45.760 16.190 45.930 16.360 ;
        RECT 46.240 16.190 46.410 16.360 ;
        RECT 46.720 16.190 46.890 16.360 ;
        RECT 47.200 16.190 47.370 16.360 ;
        RECT 47.680 16.190 47.850 16.360 ;
        RECT 48.160 16.190 48.330 16.360 ;
        RECT 48.640 16.190 48.810 16.360 ;
        RECT 49.120 16.190 49.290 16.360 ;
        RECT 49.600 16.190 49.770 16.360 ;
        RECT 50.080 16.190 50.250 16.360 ;
        RECT 50.560 16.190 50.730 16.360 ;
        RECT 51.040 16.190 51.210 16.360 ;
        RECT 51.520 16.190 51.690 16.360 ;
        RECT 52.000 16.190 52.170 16.360 ;
        RECT 52.480 16.190 52.650 16.360 ;
        RECT 52.960 16.190 53.130 16.360 ;
        RECT 53.440 16.190 53.610 16.360 ;
        RECT 53.920 16.190 54.090 16.360 ;
        RECT 54.400 16.190 54.570 16.360 ;
        RECT 54.880 16.190 55.050 16.360 ;
        RECT 55.360 16.190 55.530 16.360 ;
        RECT 55.840 16.190 56.010 16.360 ;
        RECT 56.320 16.190 56.490 16.360 ;
        RECT 56.800 16.190 56.970 16.360 ;
        RECT 57.280 16.190 57.450 16.360 ;
        RECT 57.760 16.190 57.930 16.360 ;
        RECT 58.240 16.190 58.410 16.360 ;
        RECT 58.720 16.190 58.890 16.360 ;
        RECT 59.200 16.190 59.370 16.360 ;
        RECT 59.680 16.190 59.850 16.360 ;
        RECT 60.160 16.190 60.330 16.360 ;
        RECT 60.640 16.190 60.810 16.360 ;
        RECT 61.120 16.190 61.290 16.360 ;
        RECT 61.600 16.190 61.770 16.360 ;
        RECT 62.080 16.190 62.250 16.360 ;
        RECT 62.560 16.190 62.730 16.360 ;
        RECT 63.040 16.190 63.210 16.360 ;
        RECT 63.520 16.190 63.690 16.360 ;
        RECT 64.000 16.190 64.170 16.360 ;
        RECT 64.480 16.190 64.650 16.360 ;
        RECT 64.960 16.190 65.130 16.360 ;
        RECT 65.440 16.190 65.610 16.360 ;
        RECT 65.920 16.190 66.090 16.360 ;
        RECT 66.400 16.190 66.570 16.360 ;
        RECT 66.880 16.190 67.050 16.360 ;
        RECT 67.360 16.190 67.530 16.360 ;
        RECT 67.840 16.190 68.010 16.360 ;
        RECT 68.320 16.190 68.490 16.360 ;
        RECT 68.800 16.190 68.970 16.360 ;
        RECT 69.280 16.190 69.450 16.360 ;
        RECT 69.760 16.190 69.930 16.360 ;
        RECT 70.240 16.190 70.410 16.360 ;
        RECT 70.720 16.190 70.890 16.360 ;
        RECT 71.200 16.190 71.370 16.360 ;
        RECT 71.680 16.190 71.850 16.360 ;
        RECT 72.160 16.190 72.330 16.360 ;
        RECT 72.640 16.190 72.810 16.360 ;
        RECT 73.120 16.190 73.290 16.360 ;
        RECT 73.600 16.190 73.770 16.360 ;
        RECT 74.080 16.190 74.250 16.360 ;
        RECT 74.560 16.190 74.730 16.360 ;
        RECT 75.040 16.190 75.210 16.360 ;
        RECT 75.520 16.190 75.690 16.360 ;
        RECT 76.000 16.190 76.170 16.360 ;
        RECT 76.480 16.190 76.650 16.360 ;
        RECT 76.960 16.190 77.130 16.360 ;
        RECT 77.440 16.190 77.610 16.360 ;
        RECT 77.920 16.190 78.090 16.360 ;
        RECT 78.400 16.190 78.570 16.360 ;
        RECT 78.880 16.190 79.050 16.360 ;
        RECT 79.360 16.190 79.530 16.360 ;
        RECT 79.840 16.190 80.010 16.360 ;
        RECT 80.320 16.190 80.490 16.360 ;
        RECT 80.800 16.190 80.970 16.360 ;
        RECT 81.280 16.190 81.450 16.360 ;
        RECT 81.760 16.190 81.930 16.360 ;
        RECT 82.240 16.190 82.410 16.360 ;
        RECT 82.720 16.190 82.890 16.360 ;
        RECT 83.200 16.190 83.370 16.360 ;
        RECT 83.680 16.190 83.850 16.360 ;
        RECT 84.160 16.190 84.330 16.360 ;
        RECT 84.640 16.190 84.810 16.360 ;
        RECT 85.120 16.190 85.290 16.360 ;
        RECT 85.600 16.190 85.770 16.360 ;
        RECT 86.080 16.190 86.250 16.360 ;
        RECT 86.560 16.190 86.730 16.360 ;
        RECT 87.040 16.190 87.210 16.360 ;
        RECT 87.520 16.190 87.690 16.360 ;
        RECT 88.000 16.190 88.170 16.360 ;
        RECT 88.480 16.190 88.650 16.360 ;
        RECT 88.960 16.190 89.130 16.360 ;
        RECT 89.440 16.190 89.610 16.360 ;
        RECT 89.920 16.190 90.090 16.360 ;
        RECT 90.400 16.190 90.570 16.360 ;
        RECT 90.880 16.190 91.050 16.360 ;
        RECT 91.360 16.190 91.530 16.360 ;
        RECT 91.840 16.190 92.010 16.360 ;
        RECT 92.320 16.190 92.490 16.360 ;
        RECT 92.800 16.190 92.970 16.360 ;
        RECT 93.280 16.190 93.450 16.360 ;
        RECT 93.760 16.190 93.930 16.360 ;
        RECT 94.240 16.190 94.410 16.360 ;
        RECT 94.720 16.190 94.890 16.360 ;
        RECT 95.200 16.190 95.370 16.360 ;
        RECT 95.680 16.190 95.850 16.360 ;
        RECT 96.160 16.190 96.330 16.360 ;
        RECT 96.640 16.190 96.810 16.360 ;
        RECT 97.120 16.190 97.290 16.360 ;
        RECT 97.600 16.190 97.770 16.360 ;
        RECT 98.080 16.190 98.250 16.360 ;
        RECT 98.560 16.190 98.730 16.360 ;
        RECT 99.040 16.190 99.210 16.360 ;
        RECT 99.520 16.190 99.690 16.360 ;
        RECT 100.000 16.190 100.170 16.360 ;
        RECT 100.480 16.190 100.650 16.360 ;
        RECT 100.960 16.190 101.130 16.360 ;
        RECT 101.440 16.190 101.610 16.360 ;
        RECT 101.920 16.190 102.090 16.360 ;
        RECT 102.400 16.190 102.570 16.360 ;
        RECT 102.880 16.190 103.050 16.360 ;
        RECT 103.360 16.190 103.530 16.360 ;
        RECT 103.840 16.190 104.010 16.360 ;
        RECT 104.320 16.190 104.490 16.360 ;
        RECT 104.800 16.190 104.970 16.360 ;
        RECT 105.280 16.190 105.450 16.360 ;
        RECT 105.760 16.190 105.930 16.360 ;
        RECT 106.240 16.190 106.410 16.360 ;
        RECT 106.720 16.190 106.890 16.360 ;
        RECT 107.200 16.190 107.370 16.360 ;
        RECT 107.680 16.190 107.850 16.360 ;
        RECT 108.160 16.190 108.330 16.360 ;
        RECT 108.640 16.190 108.810 16.360 ;
        RECT 109.120 16.190 109.290 16.360 ;
        RECT 109.600 16.190 109.770 16.360 ;
        RECT 110.080 16.190 110.250 16.360 ;
        RECT 110.560 16.190 110.730 16.360 ;
        RECT 111.040 16.190 111.210 16.360 ;
        RECT 111.520 16.190 111.690 16.360 ;
        RECT 112.000 16.190 112.170 16.360 ;
        RECT 112.480 16.190 112.650 16.360 ;
        RECT 112.960 16.190 113.130 16.360 ;
        RECT 113.440 16.190 113.610 16.360 ;
        RECT 113.920 16.190 114.090 16.360 ;
        RECT 114.400 16.190 114.570 16.360 ;
        RECT 114.880 16.190 115.050 16.360 ;
        RECT 115.360 16.190 115.530 16.360 ;
        RECT 115.840 16.190 116.010 16.360 ;
        RECT 116.320 16.190 116.490 16.360 ;
        RECT 116.800 16.190 116.970 16.360 ;
        RECT 117.280 16.190 117.450 16.360 ;
        RECT 117.760 16.190 117.930 16.360 ;
        RECT 118.240 16.190 118.410 16.360 ;
        RECT 118.720 16.190 118.890 16.360 ;
        RECT 119.200 16.190 119.370 16.360 ;
        RECT 119.680 16.190 119.850 16.360 ;
        RECT 120.160 16.190 120.330 16.360 ;
        RECT 120.640 16.190 120.810 16.360 ;
        RECT 121.120 16.190 121.290 16.360 ;
        RECT 121.600 16.190 121.770 16.360 ;
        RECT 122.080 16.190 122.250 16.360 ;
        RECT 122.560 16.190 122.730 16.360 ;
        RECT 123.040 16.190 123.210 16.360 ;
        RECT 123.520 16.190 123.690 16.360 ;
        RECT 124.000 16.190 124.170 16.360 ;
        RECT 124.480 16.190 124.650 16.360 ;
        RECT 124.960 16.190 125.130 16.360 ;
        RECT 125.440 16.190 125.610 16.360 ;
        RECT 125.920 16.190 126.090 16.360 ;
        RECT 126.400 16.190 126.570 16.360 ;
        RECT 126.880 16.190 127.050 16.360 ;
        RECT 127.360 16.190 127.530 16.360 ;
        RECT 127.840 16.190 128.010 16.360 ;
        RECT 128.320 16.190 128.490 16.360 ;
        RECT 128.800 16.190 128.970 16.360 ;
        RECT 129.280 16.190 129.450 16.360 ;
        RECT 129.760 16.190 129.930 16.360 ;
        RECT 130.240 16.190 130.410 16.360 ;
        RECT 130.720 16.190 130.890 16.360 ;
        RECT 131.200 16.190 131.370 16.360 ;
        RECT 131.680 16.190 131.850 16.360 ;
        RECT 132.160 16.190 132.330 16.360 ;
        RECT 132.640 16.190 132.810 16.360 ;
        RECT 133.120 16.190 133.290 16.360 ;
        RECT 133.600 16.190 133.770 16.360 ;
        RECT 134.080 16.190 134.250 16.360 ;
        RECT 134.560 16.190 134.730 16.360 ;
        RECT 135.040 16.190 135.210 16.360 ;
        RECT 135.520 16.190 135.690 16.360 ;
        RECT 136.000 16.190 136.170 16.360 ;
        RECT 136.480 16.190 136.650 16.360 ;
        RECT 136.960 16.190 137.130 16.360 ;
        RECT 137.440 16.190 137.610 16.360 ;
        RECT 137.920 16.190 138.090 16.360 ;
        RECT 138.400 16.190 138.570 16.360 ;
        RECT 138.880 16.190 139.050 16.360 ;
        RECT 139.360 16.190 139.530 16.360 ;
        RECT 139.840 16.190 140.010 16.360 ;
        RECT 140.320 16.190 140.490 16.360 ;
        RECT 140.800 16.190 140.970 16.360 ;
        RECT 141.280 16.190 141.450 16.360 ;
      LAYER li1 ;
        RECT 141.600 16.190 142.080 16.360 ;
      LAYER L1M1_PR_C ;
        RECT 17.920 146.600 18.090 146.610 ;
        RECT 36.160 146.600 36.330 146.610 ;
        RECT 43.840 146.600 44.010 146.610 ;
        RECT 85.600 146.600 85.770 146.610 ;
        RECT 141.760 146.430 141.930 146.610 ;
        RECT 30.400 138.460 30.570 138.470 ;
        RECT 29.920 138.290 30.090 138.460 ;
        RECT 62.560 138.460 62.730 138.470 ;
        RECT 75.040 138.460 75.210 138.470 ;
        RECT 98.080 138.460 98.250 138.470 ;
        RECT 109.600 138.460 109.770 138.470 ;
        RECT 141.760 138.460 141.930 138.470 ;
        RECT 31.360 130.150 31.530 130.320 ;
        RECT 34.240 130.320 34.410 130.330 ;
        RECT 43.840 130.320 44.010 130.330 ;
        RECT 73.120 130.150 73.290 130.320 ;
        RECT 74.080 130.320 74.250 130.330 ;
        RECT 110.560 130.150 110.730 130.330 ;
        RECT 118.240 130.320 118.410 130.330 ;
        RECT 141.760 130.150 141.930 130.320 ;
        RECT 7.840 122.010 8.010 122.020 ;
        RECT 10.720 122.180 10.890 122.190 ;
        RECT 28.480 122.020 28.650 122.190 ;
        RECT 43.360 122.020 43.530 122.190 ;
        RECT 43.840 122.010 44.010 122.020 ;
        RECT 50.080 122.020 50.250 122.190 ;
        RECT 67.360 122.180 67.530 122.190 ;
        RECT 100.480 122.020 100.650 122.190 ;
        RECT 141.760 122.180 141.930 122.190 ;
        RECT 13.600 113.870 13.770 114.040 ;
        RECT 24.160 114.040 24.330 114.050 ;
        RECT 37.120 114.040 37.290 114.050 ;
        RECT 71.680 114.040 71.850 114.050 ;
        RECT 88.480 113.870 88.650 114.040 ;
        RECT 116.800 113.870 116.970 114.040 ;
        RECT 40.480 105.900 40.650 105.910 ;
        RECT 61.120 105.900 61.290 105.910 ;
        RECT 73.600 105.730 73.770 105.900 ;
        RECT 116.800 105.730 116.970 105.900 ;
        RECT 121.120 105.900 121.290 105.910 ;
        RECT 141.760 105.730 141.930 105.900 ;
        RECT 21.760 97.590 21.930 97.760 ;
        RECT 28.480 97.590 28.650 97.760 ;
        RECT 32.800 97.760 32.970 97.770 ;
        RECT 72.160 97.590 72.330 97.760 ;
        RECT 74.080 97.760 74.250 97.770 ;
        RECT 98.560 97.760 98.730 97.770 ;
        RECT 121.120 97.760 121.290 97.770 ;
        RECT 141.760 97.590 141.930 97.760 ;
        RECT 12.640 89.450 12.810 89.620 ;
        RECT 20.320 89.460 20.490 89.630 ;
        RECT 56.320 89.450 56.490 89.620 ;
        RECT 68.320 89.460 68.490 89.630 ;
        RECT 101.440 89.460 101.610 89.630 ;
        RECT 117.760 89.620 117.930 89.630 ;
        RECT 134.080 89.460 134.250 89.630 ;
        RECT 141.760 89.450 141.930 89.630 ;
        RECT 14.560 81.480 14.730 81.490 ;
        RECT 64.480 81.310 64.650 81.480 ;
        RECT 71.200 81.480 71.370 81.490 ;
        RECT 80.800 81.480 80.970 81.490 ;
        RECT 104.800 81.310 104.970 81.480 ;
        RECT 141.760 81.310 141.930 81.480 ;
        RECT 47.680 73.340 47.850 73.350 ;
        RECT 47.200 73.170 47.370 73.340 ;
        RECT 59.200 73.340 59.370 73.350 ;
        RECT 76.480 73.340 76.650 73.350 ;
        RECT 78.880 73.170 79.050 73.340 ;
        RECT 134.080 73.170 134.250 73.340 ;
        RECT 141.760 73.170 141.930 73.340 ;
        RECT 8.800 65.030 8.970 65.200 ;
        RECT 47.680 65.030 47.850 65.200 ;
        RECT 91.360 65.030 91.530 65.210 ;
        RECT 105.760 65.200 105.930 65.210 ;
        RECT 130.240 65.030 130.410 65.200 ;
        RECT 141.760 65.200 141.930 65.210 ;
        RECT 49.600 56.890 49.770 57.060 ;
        RECT 101.920 57.060 102.090 57.070 ;
        RECT 115.840 57.060 116.010 57.070 ;
        RECT 141.760 56.890 141.930 57.060 ;
        RECT 7.840 48.750 8.010 48.920 ;
        RECT 47.680 48.750 47.850 48.920 ;
        RECT 50.560 48.920 50.730 48.930 ;
        RECT 81.280 48.750 81.450 48.920 ;
        RECT 94.720 48.920 94.890 48.930 ;
        RECT 107.200 48.750 107.370 48.920 ;
        RECT 108.160 48.920 108.330 48.930 ;
        RECT 123.040 48.750 123.210 48.920 ;
        RECT 141.760 48.750 141.930 48.920 ;
        RECT 14.560 40.780 14.730 40.790 ;
        RECT 77.920 40.780 78.090 40.790 ;
        RECT 110.560 40.780 110.730 40.790 ;
        RECT 115.840 40.610 116.010 40.780 ;
        RECT 141.760 40.610 141.930 40.780 ;
        RECT 40.480 32.470 40.650 32.640 ;
        RECT 104.320 32.640 104.490 32.650 ;
        RECT 119.680 32.640 119.850 32.650 ;
        RECT 132.160 32.640 132.330 32.650 ;
        RECT 141.760 32.470 141.930 32.650 ;
        RECT 14.560 24.330 14.730 24.500 ;
        RECT 16.960 24.500 17.130 24.510 ;
        RECT 52.480 24.330 52.650 24.500 ;
        RECT 81.760 24.330 81.930 24.500 ;
        RECT 88.480 24.330 88.650 24.500 ;
        RECT 94.240 24.330 94.410 24.500 ;
        RECT 141.760 24.330 141.930 24.500 ;
        RECT 37.600 16.190 37.770 16.360 ;
        RECT 141.760 16.190 141.930 16.360 ;
      LAYER met1 ;
        RECT 5.760 145.900 142.080 147.140 ;
        RECT 5.760 137.760 142.080 139.000 ;
        RECT 5.760 129.620 142.080 130.860 ;
        RECT 5.760 121.480 142.080 122.720 ;
        RECT 5.760 113.340 142.080 114.580 ;
        RECT 5.760 105.200 142.080 106.440 ;
        RECT 5.760 97.060 142.080 98.300 ;
        RECT 5.760 88.920 142.080 90.160 ;
        RECT 5.760 80.780 142.080 82.020 ;
        RECT 5.760 72.640 142.080 73.880 ;
        RECT 5.760 64.500 142.080 65.740 ;
        RECT 5.760 56.360 142.080 57.600 ;
        RECT 5.760 48.220 142.080 49.460 ;
        RECT 5.760 40.080 142.080 41.320 ;
        RECT 5.760 31.940 142.080 33.180 ;
        RECT 5.760 23.800 142.080 25.040 ;
        RECT 5.760 16.020 142.080 16.900 ;
      LAYER via ;
        RECT 27.870 146.390 28.130 146.650 ;
        RECT 28.190 146.390 28.450 146.650 ;
        RECT 28.510 146.390 28.770 146.650 ;
        RECT 28.830 146.390 29.090 146.650 ;
        RECT 73.310 146.390 73.570 146.650 ;
        RECT 73.630 146.390 73.890 146.650 ;
        RECT 73.950 146.390 74.210 146.650 ;
        RECT 74.270 146.390 74.530 146.650 ;
        RECT 118.750 146.390 119.010 146.650 ;
        RECT 119.070 146.390 119.330 146.650 ;
        RECT 119.390 146.390 119.650 146.650 ;
        RECT 119.710 146.390 119.970 146.650 ;
        RECT 27.870 138.250 28.130 138.510 ;
        RECT 28.190 138.250 28.450 138.510 ;
        RECT 28.510 138.250 28.770 138.510 ;
        RECT 28.830 138.250 29.090 138.510 ;
        RECT 73.310 138.250 73.570 138.510 ;
        RECT 73.630 138.250 73.890 138.510 ;
        RECT 73.950 138.250 74.210 138.510 ;
        RECT 74.270 138.250 74.530 138.510 ;
        RECT 118.750 138.250 119.010 138.510 ;
        RECT 119.070 138.250 119.330 138.510 ;
        RECT 119.390 138.250 119.650 138.510 ;
        RECT 119.710 138.250 119.970 138.510 ;
        RECT 27.870 130.110 28.130 130.370 ;
        RECT 28.190 130.110 28.450 130.370 ;
        RECT 28.510 130.110 28.770 130.370 ;
        RECT 28.830 130.110 29.090 130.370 ;
        RECT 73.310 130.110 73.570 130.370 ;
        RECT 73.630 130.110 73.890 130.370 ;
        RECT 73.950 130.110 74.210 130.370 ;
        RECT 74.270 130.110 74.530 130.370 ;
        RECT 118.750 130.110 119.010 130.370 ;
        RECT 119.070 130.110 119.330 130.370 ;
        RECT 119.390 130.110 119.650 130.370 ;
        RECT 119.710 130.110 119.970 130.370 ;
        RECT 27.870 121.970 28.130 122.230 ;
        RECT 28.190 121.970 28.450 122.230 ;
        RECT 28.510 121.970 28.770 122.230 ;
        RECT 28.830 121.970 29.090 122.230 ;
        RECT 73.310 121.970 73.570 122.230 ;
        RECT 73.630 121.970 73.890 122.230 ;
        RECT 73.950 121.970 74.210 122.230 ;
        RECT 74.270 121.970 74.530 122.230 ;
        RECT 118.750 121.970 119.010 122.230 ;
        RECT 119.070 121.970 119.330 122.230 ;
        RECT 119.390 121.970 119.650 122.230 ;
        RECT 119.710 121.970 119.970 122.230 ;
        RECT 27.870 113.830 28.130 114.090 ;
        RECT 28.190 113.830 28.450 114.090 ;
        RECT 28.510 113.830 28.770 114.090 ;
        RECT 28.830 113.830 29.090 114.090 ;
        RECT 73.310 113.830 73.570 114.090 ;
        RECT 73.630 113.830 73.890 114.090 ;
        RECT 73.950 113.830 74.210 114.090 ;
        RECT 74.270 113.830 74.530 114.090 ;
        RECT 118.750 113.830 119.010 114.090 ;
        RECT 119.070 113.830 119.330 114.090 ;
        RECT 119.390 113.830 119.650 114.090 ;
        RECT 119.710 113.830 119.970 114.090 ;
        RECT 27.870 105.690 28.130 105.950 ;
        RECT 28.190 105.690 28.450 105.950 ;
        RECT 28.510 105.690 28.770 105.950 ;
        RECT 28.830 105.690 29.090 105.950 ;
        RECT 73.310 105.690 73.570 105.950 ;
        RECT 73.630 105.690 73.890 105.950 ;
        RECT 73.950 105.690 74.210 105.950 ;
        RECT 74.270 105.690 74.530 105.950 ;
        RECT 118.750 105.690 119.010 105.950 ;
        RECT 119.070 105.690 119.330 105.950 ;
        RECT 119.390 105.690 119.650 105.950 ;
        RECT 119.710 105.690 119.970 105.950 ;
        RECT 27.870 97.550 28.130 97.810 ;
        RECT 28.190 97.550 28.450 97.810 ;
        RECT 28.510 97.550 28.770 97.810 ;
        RECT 28.830 97.550 29.090 97.810 ;
        RECT 73.310 97.550 73.570 97.810 ;
        RECT 73.630 97.550 73.890 97.810 ;
        RECT 73.950 97.550 74.210 97.810 ;
        RECT 74.270 97.550 74.530 97.810 ;
        RECT 118.750 97.550 119.010 97.810 ;
        RECT 119.070 97.550 119.330 97.810 ;
        RECT 119.390 97.550 119.650 97.810 ;
        RECT 119.710 97.550 119.970 97.810 ;
        RECT 27.870 89.410 28.130 89.670 ;
        RECT 28.190 89.410 28.450 89.670 ;
        RECT 28.510 89.410 28.770 89.670 ;
        RECT 28.830 89.410 29.090 89.670 ;
        RECT 73.310 89.410 73.570 89.670 ;
        RECT 73.630 89.410 73.890 89.670 ;
        RECT 73.950 89.410 74.210 89.670 ;
        RECT 74.270 89.410 74.530 89.670 ;
        RECT 118.750 89.410 119.010 89.670 ;
        RECT 119.070 89.410 119.330 89.670 ;
        RECT 119.390 89.410 119.650 89.670 ;
        RECT 119.710 89.410 119.970 89.670 ;
        RECT 27.870 81.270 28.130 81.530 ;
        RECT 28.190 81.270 28.450 81.530 ;
        RECT 28.510 81.270 28.770 81.530 ;
        RECT 28.830 81.270 29.090 81.530 ;
        RECT 73.310 81.270 73.570 81.530 ;
        RECT 73.630 81.270 73.890 81.530 ;
        RECT 73.950 81.270 74.210 81.530 ;
        RECT 74.270 81.270 74.530 81.530 ;
        RECT 118.750 81.270 119.010 81.530 ;
        RECT 119.070 81.270 119.330 81.530 ;
        RECT 119.390 81.270 119.650 81.530 ;
        RECT 119.710 81.270 119.970 81.530 ;
        RECT 27.870 73.130 28.130 73.390 ;
        RECT 28.190 73.130 28.450 73.390 ;
        RECT 28.510 73.130 28.770 73.390 ;
        RECT 28.830 73.130 29.090 73.390 ;
        RECT 73.310 73.130 73.570 73.390 ;
        RECT 73.630 73.130 73.890 73.390 ;
        RECT 73.950 73.130 74.210 73.390 ;
        RECT 74.270 73.130 74.530 73.390 ;
        RECT 118.750 73.130 119.010 73.390 ;
        RECT 119.070 73.130 119.330 73.390 ;
        RECT 119.390 73.130 119.650 73.390 ;
        RECT 119.710 73.130 119.970 73.390 ;
        RECT 27.870 64.990 28.130 65.250 ;
        RECT 28.190 64.990 28.450 65.250 ;
        RECT 28.510 64.990 28.770 65.250 ;
        RECT 28.830 64.990 29.090 65.250 ;
        RECT 73.310 64.990 73.570 65.250 ;
        RECT 73.630 64.990 73.890 65.250 ;
        RECT 73.950 64.990 74.210 65.250 ;
        RECT 74.270 64.990 74.530 65.250 ;
        RECT 118.750 64.990 119.010 65.250 ;
        RECT 119.070 64.990 119.330 65.250 ;
        RECT 119.390 64.990 119.650 65.250 ;
        RECT 119.710 64.990 119.970 65.250 ;
        RECT 27.870 56.850 28.130 57.110 ;
        RECT 28.190 56.850 28.450 57.110 ;
        RECT 28.510 56.850 28.770 57.110 ;
        RECT 28.830 56.850 29.090 57.110 ;
        RECT 73.310 56.850 73.570 57.110 ;
        RECT 73.630 56.850 73.890 57.110 ;
        RECT 73.950 56.850 74.210 57.110 ;
        RECT 74.270 56.850 74.530 57.110 ;
        RECT 118.750 56.850 119.010 57.110 ;
        RECT 119.070 56.850 119.330 57.110 ;
        RECT 119.390 56.850 119.650 57.110 ;
        RECT 119.710 56.850 119.970 57.110 ;
        RECT 27.870 48.710 28.130 48.970 ;
        RECT 28.190 48.710 28.450 48.970 ;
        RECT 28.510 48.710 28.770 48.970 ;
        RECT 28.830 48.710 29.090 48.970 ;
        RECT 73.310 48.710 73.570 48.970 ;
        RECT 73.630 48.710 73.890 48.970 ;
        RECT 73.950 48.710 74.210 48.970 ;
        RECT 74.270 48.710 74.530 48.970 ;
        RECT 118.750 48.710 119.010 48.970 ;
        RECT 119.070 48.710 119.330 48.970 ;
        RECT 119.390 48.710 119.650 48.970 ;
        RECT 119.710 48.710 119.970 48.970 ;
        RECT 27.870 40.570 28.130 40.830 ;
        RECT 28.190 40.570 28.450 40.830 ;
        RECT 28.510 40.570 28.770 40.830 ;
        RECT 28.830 40.570 29.090 40.830 ;
        RECT 73.310 40.570 73.570 40.830 ;
        RECT 73.630 40.570 73.890 40.830 ;
        RECT 73.950 40.570 74.210 40.830 ;
        RECT 74.270 40.570 74.530 40.830 ;
        RECT 118.750 40.570 119.010 40.830 ;
        RECT 119.070 40.570 119.330 40.830 ;
        RECT 119.390 40.570 119.650 40.830 ;
        RECT 119.710 40.570 119.970 40.830 ;
        RECT 27.870 32.430 28.130 32.690 ;
        RECT 28.190 32.430 28.450 32.690 ;
        RECT 28.510 32.430 28.770 32.690 ;
        RECT 28.830 32.430 29.090 32.690 ;
        RECT 73.310 32.430 73.570 32.690 ;
        RECT 73.630 32.430 73.890 32.690 ;
        RECT 73.950 32.430 74.210 32.690 ;
        RECT 74.270 32.430 74.530 32.690 ;
        RECT 118.750 32.430 119.010 32.690 ;
        RECT 119.070 32.430 119.330 32.690 ;
        RECT 119.390 32.430 119.650 32.690 ;
        RECT 119.710 32.430 119.970 32.690 ;
        RECT 27.870 24.290 28.130 24.550 ;
        RECT 28.190 24.290 28.450 24.550 ;
        RECT 28.510 24.290 28.770 24.550 ;
        RECT 28.830 24.290 29.090 24.550 ;
        RECT 73.310 24.290 73.570 24.550 ;
        RECT 73.630 24.290 73.890 24.550 ;
        RECT 73.950 24.290 74.210 24.550 ;
        RECT 74.270 24.290 74.530 24.550 ;
        RECT 118.750 24.290 119.010 24.550 ;
        RECT 119.070 24.290 119.330 24.550 ;
        RECT 119.390 24.290 119.650 24.550 ;
        RECT 119.710 24.290 119.970 24.550 ;
        RECT 27.870 16.150 28.130 16.410 ;
        RECT 28.190 16.150 28.450 16.410 ;
        RECT 28.510 16.150 28.770 16.410 ;
        RECT 28.830 16.150 29.090 16.410 ;
        RECT 73.310 16.150 73.570 16.410 ;
        RECT 73.630 16.150 73.890 16.410 ;
        RECT 73.950 16.150 74.210 16.410 ;
        RECT 74.270 16.150 74.530 16.410 ;
        RECT 118.750 16.150 119.010 16.410 ;
        RECT 119.070 16.150 119.330 16.410 ;
        RECT 119.390 16.150 119.650 16.410 ;
        RECT 119.710 16.150 119.970 16.410 ;
      LAYER met2 ;
        RECT 27.740 146.260 29.220 146.770 ;
        RECT 73.180 146.260 74.660 146.770 ;
        RECT 118.620 146.260 120.100 146.770 ;
        RECT 27.740 138.120 29.220 138.630 ;
        RECT 73.180 138.120 74.660 138.630 ;
        RECT 118.620 138.120 120.100 138.630 ;
        RECT 27.740 129.980 29.220 130.490 ;
        RECT 73.180 129.980 74.660 130.490 ;
        RECT 118.620 129.980 120.100 130.490 ;
        RECT 27.740 121.840 29.220 122.350 ;
        RECT 73.180 121.840 74.660 122.350 ;
        RECT 118.620 121.840 120.100 122.350 ;
        RECT 27.740 113.700 29.220 114.210 ;
        RECT 73.180 113.700 74.660 114.210 ;
        RECT 118.620 113.700 120.100 114.210 ;
        RECT 27.740 105.560 29.220 106.070 ;
        RECT 73.180 105.560 74.660 106.070 ;
        RECT 118.620 105.560 120.100 106.070 ;
        RECT 27.740 97.420 29.220 97.930 ;
        RECT 73.180 97.420 74.660 97.930 ;
        RECT 118.620 97.420 120.100 97.930 ;
        RECT 27.740 89.280 29.220 89.790 ;
        RECT 73.180 89.280 74.660 89.790 ;
        RECT 118.620 89.280 120.100 89.790 ;
        RECT 27.740 81.140 29.220 81.650 ;
        RECT 73.180 81.140 74.660 81.650 ;
        RECT 118.620 81.140 120.100 81.650 ;
        RECT 27.740 73.000 29.220 73.510 ;
        RECT 73.180 73.000 74.660 73.510 ;
        RECT 118.620 73.000 120.100 73.510 ;
        RECT 27.740 64.860 29.220 65.370 ;
        RECT 73.180 64.860 74.660 65.370 ;
        RECT 118.620 64.860 120.100 65.370 ;
        RECT 27.740 56.720 29.220 57.230 ;
        RECT 73.180 56.720 74.660 57.230 ;
        RECT 118.620 56.720 120.100 57.230 ;
        RECT 27.740 48.580 29.220 49.090 ;
        RECT 73.180 48.580 74.660 49.090 ;
        RECT 118.620 48.580 120.100 49.090 ;
        RECT 27.740 40.440 29.220 40.950 ;
        RECT 73.180 40.440 74.660 40.950 ;
        RECT 118.620 40.440 120.100 40.950 ;
        RECT 27.740 32.300 29.220 32.810 ;
        RECT 73.180 32.300 74.660 32.810 ;
        RECT 118.620 32.300 120.100 32.810 ;
        RECT 27.740 24.160 29.220 24.670 ;
        RECT 73.180 24.160 74.660 24.670 ;
        RECT 118.620 24.160 120.100 24.670 ;
        RECT 27.740 16.020 29.220 16.530 ;
        RECT 73.180 16.020 74.660 16.530 ;
        RECT 118.620 16.020 120.100 16.530 ;
      LAYER via2 ;
        RECT 27.740 146.380 28.020 146.660 ;
        RECT 28.140 146.380 28.420 146.660 ;
        RECT 28.540 146.380 28.820 146.660 ;
        RECT 28.940 146.380 29.220 146.660 ;
        RECT 73.180 146.380 73.460 146.660 ;
        RECT 73.580 146.380 73.860 146.660 ;
        RECT 73.980 146.380 74.260 146.660 ;
        RECT 74.380 146.380 74.660 146.660 ;
        RECT 118.620 146.380 118.900 146.660 ;
        RECT 119.020 146.380 119.300 146.660 ;
        RECT 119.420 146.380 119.700 146.660 ;
        RECT 119.820 146.380 120.100 146.660 ;
        RECT 27.740 138.240 28.020 138.520 ;
        RECT 28.140 138.240 28.420 138.520 ;
        RECT 28.540 138.240 28.820 138.520 ;
        RECT 28.940 138.240 29.220 138.520 ;
        RECT 73.180 138.240 73.460 138.520 ;
        RECT 73.580 138.240 73.860 138.520 ;
        RECT 73.980 138.240 74.260 138.520 ;
        RECT 74.380 138.240 74.660 138.520 ;
        RECT 118.620 138.240 118.900 138.520 ;
        RECT 119.020 138.240 119.300 138.520 ;
        RECT 119.420 138.240 119.700 138.520 ;
        RECT 119.820 138.240 120.100 138.520 ;
        RECT 27.740 130.100 28.020 130.380 ;
        RECT 28.140 130.100 28.420 130.380 ;
        RECT 28.540 130.100 28.820 130.380 ;
        RECT 28.940 130.100 29.220 130.380 ;
        RECT 73.180 130.100 73.460 130.380 ;
        RECT 73.580 130.100 73.860 130.380 ;
        RECT 73.980 130.100 74.260 130.380 ;
        RECT 74.380 130.100 74.660 130.380 ;
        RECT 118.620 130.100 118.900 130.380 ;
        RECT 119.020 130.100 119.300 130.380 ;
        RECT 119.420 130.100 119.700 130.380 ;
        RECT 119.820 130.100 120.100 130.380 ;
        RECT 27.740 121.960 28.020 122.240 ;
        RECT 28.140 121.960 28.420 122.240 ;
        RECT 28.540 121.960 28.820 122.240 ;
        RECT 28.940 121.960 29.220 122.240 ;
        RECT 73.180 121.960 73.460 122.240 ;
        RECT 73.580 121.960 73.860 122.240 ;
        RECT 73.980 121.960 74.260 122.240 ;
        RECT 74.380 121.960 74.660 122.240 ;
        RECT 118.620 121.960 118.900 122.240 ;
        RECT 119.020 121.960 119.300 122.240 ;
        RECT 119.420 121.960 119.700 122.240 ;
        RECT 119.820 121.960 120.100 122.240 ;
        RECT 27.740 113.820 28.020 114.100 ;
        RECT 28.140 113.820 28.420 114.100 ;
        RECT 28.540 113.820 28.820 114.100 ;
        RECT 28.940 113.820 29.220 114.100 ;
        RECT 73.180 113.820 73.460 114.100 ;
        RECT 73.580 113.820 73.860 114.100 ;
        RECT 73.980 113.820 74.260 114.100 ;
        RECT 74.380 113.820 74.660 114.100 ;
        RECT 118.620 113.820 118.900 114.100 ;
        RECT 119.020 113.820 119.300 114.100 ;
        RECT 119.420 113.820 119.700 114.100 ;
        RECT 119.820 113.820 120.100 114.100 ;
        RECT 27.740 105.680 28.020 105.960 ;
        RECT 28.140 105.680 28.420 105.960 ;
        RECT 28.540 105.680 28.820 105.960 ;
        RECT 28.940 105.680 29.220 105.960 ;
        RECT 73.180 105.680 73.460 105.960 ;
        RECT 73.580 105.680 73.860 105.960 ;
        RECT 73.980 105.680 74.260 105.960 ;
        RECT 74.380 105.680 74.660 105.960 ;
        RECT 118.620 105.680 118.900 105.960 ;
        RECT 119.020 105.680 119.300 105.960 ;
        RECT 119.420 105.680 119.700 105.960 ;
        RECT 119.820 105.680 120.100 105.960 ;
        RECT 27.740 97.540 28.020 97.820 ;
        RECT 28.140 97.540 28.420 97.820 ;
        RECT 28.540 97.540 28.820 97.820 ;
        RECT 28.940 97.540 29.220 97.820 ;
        RECT 73.180 97.540 73.460 97.820 ;
        RECT 73.580 97.540 73.860 97.820 ;
        RECT 73.980 97.540 74.260 97.820 ;
        RECT 74.380 97.540 74.660 97.820 ;
        RECT 118.620 97.540 118.900 97.820 ;
        RECT 119.020 97.540 119.300 97.820 ;
        RECT 119.420 97.540 119.700 97.820 ;
        RECT 119.820 97.540 120.100 97.820 ;
        RECT 27.740 89.400 28.020 89.680 ;
        RECT 28.140 89.400 28.420 89.680 ;
        RECT 28.540 89.400 28.820 89.680 ;
        RECT 28.940 89.400 29.220 89.680 ;
        RECT 73.180 89.400 73.460 89.680 ;
        RECT 73.580 89.400 73.860 89.680 ;
        RECT 73.980 89.400 74.260 89.680 ;
        RECT 74.380 89.400 74.660 89.680 ;
        RECT 118.620 89.400 118.900 89.680 ;
        RECT 119.020 89.400 119.300 89.680 ;
        RECT 119.420 89.400 119.700 89.680 ;
        RECT 119.820 89.400 120.100 89.680 ;
        RECT 27.740 81.260 28.020 81.540 ;
        RECT 28.140 81.260 28.420 81.540 ;
        RECT 28.540 81.260 28.820 81.540 ;
        RECT 28.940 81.260 29.220 81.540 ;
        RECT 73.180 81.260 73.460 81.540 ;
        RECT 73.580 81.260 73.860 81.540 ;
        RECT 73.980 81.260 74.260 81.540 ;
        RECT 74.380 81.260 74.660 81.540 ;
        RECT 118.620 81.260 118.900 81.540 ;
        RECT 119.020 81.260 119.300 81.540 ;
        RECT 119.420 81.260 119.700 81.540 ;
        RECT 119.820 81.260 120.100 81.540 ;
        RECT 27.740 73.120 28.020 73.400 ;
        RECT 28.140 73.120 28.420 73.400 ;
        RECT 28.540 73.120 28.820 73.400 ;
        RECT 28.940 73.120 29.220 73.400 ;
        RECT 73.180 73.120 73.460 73.400 ;
        RECT 73.580 73.120 73.860 73.400 ;
        RECT 73.980 73.120 74.260 73.400 ;
        RECT 74.380 73.120 74.660 73.400 ;
        RECT 118.620 73.120 118.900 73.400 ;
        RECT 119.020 73.120 119.300 73.400 ;
        RECT 119.420 73.120 119.700 73.400 ;
        RECT 119.820 73.120 120.100 73.400 ;
        RECT 27.740 64.980 28.020 65.260 ;
        RECT 28.140 64.980 28.420 65.260 ;
        RECT 28.540 64.980 28.820 65.260 ;
        RECT 28.940 64.980 29.220 65.260 ;
        RECT 73.180 64.980 73.460 65.260 ;
        RECT 73.580 64.980 73.860 65.260 ;
        RECT 73.980 64.980 74.260 65.260 ;
        RECT 74.380 64.980 74.660 65.260 ;
        RECT 118.620 64.980 118.900 65.260 ;
        RECT 119.020 64.980 119.300 65.260 ;
        RECT 119.420 64.980 119.700 65.260 ;
        RECT 119.820 64.980 120.100 65.260 ;
        RECT 27.740 56.840 28.020 57.120 ;
        RECT 28.140 56.840 28.420 57.120 ;
        RECT 28.540 56.840 28.820 57.120 ;
        RECT 28.940 56.840 29.220 57.120 ;
        RECT 73.180 56.840 73.460 57.120 ;
        RECT 73.580 56.840 73.860 57.120 ;
        RECT 73.980 56.840 74.260 57.120 ;
        RECT 74.380 56.840 74.660 57.120 ;
        RECT 118.620 56.840 118.900 57.120 ;
        RECT 119.020 56.840 119.300 57.120 ;
        RECT 119.420 56.840 119.700 57.120 ;
        RECT 119.820 56.840 120.100 57.120 ;
        RECT 27.740 48.700 28.020 48.980 ;
        RECT 28.140 48.700 28.420 48.980 ;
        RECT 28.540 48.700 28.820 48.980 ;
        RECT 28.940 48.700 29.220 48.980 ;
        RECT 73.180 48.700 73.460 48.980 ;
        RECT 73.580 48.700 73.860 48.980 ;
        RECT 73.980 48.700 74.260 48.980 ;
        RECT 74.380 48.700 74.660 48.980 ;
        RECT 118.620 48.700 118.900 48.980 ;
        RECT 119.020 48.700 119.300 48.980 ;
        RECT 119.420 48.700 119.700 48.980 ;
        RECT 119.820 48.700 120.100 48.980 ;
        RECT 27.740 40.560 28.020 40.840 ;
        RECT 28.140 40.560 28.420 40.840 ;
        RECT 28.540 40.560 28.820 40.840 ;
        RECT 28.940 40.560 29.220 40.840 ;
        RECT 73.180 40.560 73.460 40.840 ;
        RECT 73.580 40.560 73.860 40.840 ;
        RECT 73.980 40.560 74.260 40.840 ;
        RECT 74.380 40.560 74.660 40.840 ;
        RECT 118.620 40.560 118.900 40.840 ;
        RECT 119.020 40.560 119.300 40.840 ;
        RECT 119.420 40.560 119.700 40.840 ;
        RECT 119.820 40.560 120.100 40.840 ;
        RECT 27.740 32.420 28.020 32.700 ;
        RECT 28.140 32.420 28.420 32.700 ;
        RECT 28.540 32.420 28.820 32.700 ;
        RECT 28.940 32.420 29.220 32.700 ;
        RECT 73.180 32.420 73.460 32.700 ;
        RECT 73.580 32.420 73.860 32.700 ;
        RECT 73.980 32.420 74.260 32.700 ;
        RECT 74.380 32.420 74.660 32.700 ;
        RECT 118.620 32.420 118.900 32.700 ;
        RECT 119.020 32.420 119.300 32.700 ;
        RECT 119.420 32.420 119.700 32.700 ;
        RECT 119.820 32.420 120.100 32.700 ;
        RECT 27.740 24.280 28.020 24.560 ;
        RECT 28.140 24.280 28.420 24.560 ;
        RECT 28.540 24.280 28.820 24.560 ;
        RECT 28.940 24.280 29.220 24.560 ;
        RECT 73.180 24.280 73.460 24.560 ;
        RECT 73.580 24.280 73.860 24.560 ;
        RECT 73.980 24.280 74.260 24.560 ;
        RECT 74.380 24.280 74.660 24.560 ;
        RECT 118.620 24.280 118.900 24.560 ;
        RECT 119.020 24.280 119.300 24.560 ;
        RECT 119.420 24.280 119.700 24.560 ;
        RECT 119.820 24.280 120.100 24.560 ;
        RECT 27.740 16.140 28.020 16.420 ;
        RECT 28.140 16.140 28.420 16.420 ;
        RECT 28.540 16.140 28.820 16.420 ;
        RECT 28.940 16.140 29.220 16.420 ;
        RECT 73.180 16.140 73.460 16.420 ;
        RECT 73.580 16.140 73.860 16.420 ;
        RECT 73.980 16.140 74.260 16.420 ;
        RECT 74.380 16.140 74.660 16.420 ;
        RECT 118.620 16.140 118.900 16.420 ;
        RECT 119.020 16.140 119.300 16.420 ;
        RECT 119.420 16.140 119.700 16.420 ;
        RECT 119.820 16.140 120.100 16.420 ;
      LAYER met3 ;
        RECT 27.680 146.350 29.280 146.680 ;
        RECT 73.120 146.350 74.720 146.680 ;
        RECT 118.560 146.350 120.160 146.680 ;
        RECT 27.680 138.210 29.280 138.540 ;
        RECT 73.120 138.210 74.720 138.540 ;
        RECT 118.560 138.210 120.160 138.540 ;
        RECT 27.680 130.070 29.280 130.400 ;
        RECT 73.120 130.070 74.720 130.400 ;
        RECT 118.560 130.070 120.160 130.400 ;
        RECT 27.680 121.930 29.280 122.260 ;
        RECT 73.120 121.930 74.720 122.260 ;
        RECT 118.560 121.930 120.160 122.260 ;
        RECT 27.680 113.790 29.280 114.120 ;
        RECT 73.120 113.790 74.720 114.120 ;
        RECT 118.560 113.790 120.160 114.120 ;
        RECT 27.680 105.650 29.280 105.980 ;
        RECT 73.120 105.650 74.720 105.980 ;
        RECT 118.560 105.650 120.160 105.980 ;
        RECT 27.680 97.510 29.280 97.840 ;
        RECT 73.120 97.510 74.720 97.840 ;
        RECT 118.560 97.510 120.160 97.840 ;
        RECT 27.680 89.370 29.280 89.700 ;
        RECT 73.120 89.370 74.720 89.700 ;
        RECT 118.560 89.370 120.160 89.700 ;
        RECT 27.680 81.230 29.280 81.560 ;
        RECT 73.120 81.230 74.720 81.560 ;
        RECT 118.560 81.230 120.160 81.560 ;
        RECT 27.680 73.090 29.280 73.420 ;
        RECT 73.120 73.090 74.720 73.420 ;
        RECT 118.560 73.090 120.160 73.420 ;
        RECT 27.680 64.950 29.280 65.280 ;
        RECT 73.120 64.950 74.720 65.280 ;
        RECT 118.560 64.950 120.160 65.280 ;
        RECT 27.680 56.810 29.280 57.140 ;
        RECT 73.120 56.810 74.720 57.140 ;
        RECT 118.560 56.810 120.160 57.140 ;
        RECT 27.680 48.670 29.280 49.000 ;
        RECT 73.120 48.670 74.720 49.000 ;
        RECT 118.560 48.670 120.160 49.000 ;
        RECT 27.680 40.530 29.280 40.860 ;
        RECT 73.120 40.530 74.720 40.860 ;
        RECT 118.560 40.530 120.160 40.860 ;
        RECT 27.680 32.390 29.280 32.720 ;
        RECT 73.120 32.390 74.720 32.720 ;
        RECT 118.560 32.390 120.160 32.720 ;
        RECT 27.680 24.250 29.280 24.580 ;
        RECT 73.120 24.250 74.720 24.580 ;
        RECT 118.560 24.250 120.160 24.580 ;
        RECT 27.680 16.110 29.280 16.440 ;
        RECT 73.120 16.110 74.720 16.440 ;
        RECT 118.560 16.110 120.160 16.440 ;
      LAYER via3 ;
        RECT 27.720 146.360 28.040 146.680 ;
        RECT 28.120 146.360 28.440 146.680 ;
        RECT 28.520 146.360 28.840 146.680 ;
        RECT 28.920 146.360 29.240 146.680 ;
        RECT 73.160 146.360 73.480 146.680 ;
        RECT 73.560 146.360 73.880 146.680 ;
        RECT 73.960 146.360 74.280 146.680 ;
        RECT 74.360 146.360 74.680 146.680 ;
        RECT 118.600 146.360 118.920 146.680 ;
        RECT 119.000 146.360 119.320 146.680 ;
        RECT 119.400 146.360 119.720 146.680 ;
        RECT 119.800 146.360 120.120 146.680 ;
        RECT 27.720 138.220 28.040 138.540 ;
        RECT 28.120 138.220 28.440 138.540 ;
        RECT 28.520 138.220 28.840 138.540 ;
        RECT 28.920 138.220 29.240 138.540 ;
        RECT 73.160 138.220 73.480 138.540 ;
        RECT 73.560 138.220 73.880 138.540 ;
        RECT 73.960 138.220 74.280 138.540 ;
        RECT 74.360 138.220 74.680 138.540 ;
        RECT 118.600 138.220 118.920 138.540 ;
        RECT 119.000 138.220 119.320 138.540 ;
        RECT 119.400 138.220 119.720 138.540 ;
        RECT 119.800 138.220 120.120 138.540 ;
        RECT 27.720 130.080 28.040 130.400 ;
        RECT 28.120 130.080 28.440 130.400 ;
        RECT 28.520 130.080 28.840 130.400 ;
        RECT 28.920 130.080 29.240 130.400 ;
        RECT 73.160 130.080 73.480 130.400 ;
        RECT 73.560 130.080 73.880 130.400 ;
        RECT 73.960 130.080 74.280 130.400 ;
        RECT 74.360 130.080 74.680 130.400 ;
        RECT 118.600 130.080 118.920 130.400 ;
        RECT 119.000 130.080 119.320 130.400 ;
        RECT 119.400 130.080 119.720 130.400 ;
        RECT 119.800 130.080 120.120 130.400 ;
        RECT 27.720 121.940 28.040 122.260 ;
        RECT 28.120 121.940 28.440 122.260 ;
        RECT 28.520 121.940 28.840 122.260 ;
        RECT 28.920 121.940 29.240 122.260 ;
        RECT 73.160 121.940 73.480 122.260 ;
        RECT 73.560 121.940 73.880 122.260 ;
        RECT 73.960 121.940 74.280 122.260 ;
        RECT 74.360 121.940 74.680 122.260 ;
        RECT 118.600 121.940 118.920 122.260 ;
        RECT 119.000 121.940 119.320 122.260 ;
        RECT 119.400 121.940 119.720 122.260 ;
        RECT 119.800 121.940 120.120 122.260 ;
        RECT 27.720 113.800 28.040 114.120 ;
        RECT 28.120 113.800 28.440 114.120 ;
        RECT 28.520 113.800 28.840 114.120 ;
        RECT 28.920 113.800 29.240 114.120 ;
        RECT 73.160 113.800 73.480 114.120 ;
        RECT 73.560 113.800 73.880 114.120 ;
        RECT 73.960 113.800 74.280 114.120 ;
        RECT 74.360 113.800 74.680 114.120 ;
        RECT 118.600 113.800 118.920 114.120 ;
        RECT 119.000 113.800 119.320 114.120 ;
        RECT 119.400 113.800 119.720 114.120 ;
        RECT 119.800 113.800 120.120 114.120 ;
        RECT 27.720 105.660 28.040 105.980 ;
        RECT 28.120 105.660 28.440 105.980 ;
        RECT 28.520 105.660 28.840 105.980 ;
        RECT 28.920 105.660 29.240 105.980 ;
        RECT 73.160 105.660 73.480 105.980 ;
        RECT 73.560 105.660 73.880 105.980 ;
        RECT 73.960 105.660 74.280 105.980 ;
        RECT 74.360 105.660 74.680 105.980 ;
        RECT 118.600 105.660 118.920 105.980 ;
        RECT 119.000 105.660 119.320 105.980 ;
        RECT 119.400 105.660 119.720 105.980 ;
        RECT 119.800 105.660 120.120 105.980 ;
        RECT 27.720 97.520 28.040 97.840 ;
        RECT 28.120 97.520 28.440 97.840 ;
        RECT 28.520 97.520 28.840 97.840 ;
        RECT 28.920 97.520 29.240 97.840 ;
        RECT 73.160 97.520 73.480 97.840 ;
        RECT 73.560 97.520 73.880 97.840 ;
        RECT 73.960 97.520 74.280 97.840 ;
        RECT 74.360 97.520 74.680 97.840 ;
        RECT 118.600 97.520 118.920 97.840 ;
        RECT 119.000 97.520 119.320 97.840 ;
        RECT 119.400 97.520 119.720 97.840 ;
        RECT 119.800 97.520 120.120 97.840 ;
        RECT 27.720 89.380 28.040 89.700 ;
        RECT 28.120 89.380 28.440 89.700 ;
        RECT 28.520 89.380 28.840 89.700 ;
        RECT 28.920 89.380 29.240 89.700 ;
        RECT 73.160 89.380 73.480 89.700 ;
        RECT 73.560 89.380 73.880 89.700 ;
        RECT 73.960 89.380 74.280 89.700 ;
        RECT 74.360 89.380 74.680 89.700 ;
        RECT 118.600 89.380 118.920 89.700 ;
        RECT 119.000 89.380 119.320 89.700 ;
        RECT 119.400 89.380 119.720 89.700 ;
        RECT 119.800 89.380 120.120 89.700 ;
        RECT 27.720 81.240 28.040 81.560 ;
        RECT 28.120 81.240 28.440 81.560 ;
        RECT 28.520 81.240 28.840 81.560 ;
        RECT 28.920 81.240 29.240 81.560 ;
        RECT 73.160 81.240 73.480 81.560 ;
        RECT 73.560 81.240 73.880 81.560 ;
        RECT 73.960 81.240 74.280 81.560 ;
        RECT 74.360 81.240 74.680 81.560 ;
        RECT 118.600 81.240 118.920 81.560 ;
        RECT 119.000 81.240 119.320 81.560 ;
        RECT 119.400 81.240 119.720 81.560 ;
        RECT 119.800 81.240 120.120 81.560 ;
        RECT 27.720 73.100 28.040 73.420 ;
        RECT 28.120 73.100 28.440 73.420 ;
        RECT 28.520 73.100 28.840 73.420 ;
        RECT 28.920 73.100 29.240 73.420 ;
        RECT 73.160 73.100 73.480 73.420 ;
        RECT 73.560 73.100 73.880 73.420 ;
        RECT 73.960 73.100 74.280 73.420 ;
        RECT 74.360 73.100 74.680 73.420 ;
        RECT 118.600 73.100 118.920 73.420 ;
        RECT 119.000 73.100 119.320 73.420 ;
        RECT 119.400 73.100 119.720 73.420 ;
        RECT 119.800 73.100 120.120 73.420 ;
        RECT 27.720 64.960 28.040 65.280 ;
        RECT 28.120 64.960 28.440 65.280 ;
        RECT 28.520 64.960 28.840 65.280 ;
        RECT 28.920 64.960 29.240 65.280 ;
        RECT 73.160 64.960 73.480 65.280 ;
        RECT 73.560 64.960 73.880 65.280 ;
        RECT 73.960 64.960 74.280 65.280 ;
        RECT 74.360 64.960 74.680 65.280 ;
        RECT 118.600 64.960 118.920 65.280 ;
        RECT 119.000 64.960 119.320 65.280 ;
        RECT 119.400 64.960 119.720 65.280 ;
        RECT 119.800 64.960 120.120 65.280 ;
        RECT 27.720 56.820 28.040 57.140 ;
        RECT 28.120 56.820 28.440 57.140 ;
        RECT 28.520 56.820 28.840 57.140 ;
        RECT 28.920 56.820 29.240 57.140 ;
        RECT 73.160 56.820 73.480 57.140 ;
        RECT 73.560 56.820 73.880 57.140 ;
        RECT 73.960 56.820 74.280 57.140 ;
        RECT 74.360 56.820 74.680 57.140 ;
        RECT 118.600 56.820 118.920 57.140 ;
        RECT 119.000 56.820 119.320 57.140 ;
        RECT 119.400 56.820 119.720 57.140 ;
        RECT 119.800 56.820 120.120 57.140 ;
        RECT 27.720 48.680 28.040 49.000 ;
        RECT 28.120 48.680 28.440 49.000 ;
        RECT 28.520 48.680 28.840 49.000 ;
        RECT 28.920 48.680 29.240 49.000 ;
        RECT 73.160 48.680 73.480 49.000 ;
        RECT 73.560 48.680 73.880 49.000 ;
        RECT 73.960 48.680 74.280 49.000 ;
        RECT 74.360 48.680 74.680 49.000 ;
        RECT 118.600 48.680 118.920 49.000 ;
        RECT 119.000 48.680 119.320 49.000 ;
        RECT 119.400 48.680 119.720 49.000 ;
        RECT 119.800 48.680 120.120 49.000 ;
        RECT 27.720 40.540 28.040 40.860 ;
        RECT 28.120 40.540 28.440 40.860 ;
        RECT 28.520 40.540 28.840 40.860 ;
        RECT 28.920 40.540 29.240 40.860 ;
        RECT 73.160 40.540 73.480 40.860 ;
        RECT 73.560 40.540 73.880 40.860 ;
        RECT 73.960 40.540 74.280 40.860 ;
        RECT 74.360 40.540 74.680 40.860 ;
        RECT 118.600 40.540 118.920 40.860 ;
        RECT 119.000 40.540 119.320 40.860 ;
        RECT 119.400 40.540 119.720 40.860 ;
        RECT 119.800 40.540 120.120 40.860 ;
        RECT 27.720 32.400 28.040 32.720 ;
        RECT 28.120 32.400 28.440 32.720 ;
        RECT 28.520 32.400 28.840 32.720 ;
        RECT 28.920 32.400 29.240 32.720 ;
        RECT 73.160 32.400 73.480 32.720 ;
        RECT 73.560 32.400 73.880 32.720 ;
        RECT 73.960 32.400 74.280 32.720 ;
        RECT 74.360 32.400 74.680 32.720 ;
        RECT 118.600 32.400 118.920 32.720 ;
        RECT 119.000 32.400 119.320 32.720 ;
        RECT 119.400 32.400 119.720 32.720 ;
        RECT 119.800 32.400 120.120 32.720 ;
        RECT 27.720 24.260 28.040 24.580 ;
        RECT 28.120 24.260 28.440 24.580 ;
        RECT 28.520 24.260 28.840 24.580 ;
        RECT 28.920 24.260 29.240 24.580 ;
        RECT 73.160 24.260 73.480 24.580 ;
        RECT 73.560 24.260 73.880 24.580 ;
        RECT 73.960 24.260 74.280 24.580 ;
        RECT 74.360 24.260 74.680 24.580 ;
        RECT 118.600 24.260 118.920 24.580 ;
        RECT 119.000 24.260 119.320 24.580 ;
        RECT 119.400 24.260 119.720 24.580 ;
        RECT 119.800 24.260 120.120 24.580 ;
        RECT 27.720 16.120 28.040 16.440 ;
        RECT 28.120 16.120 28.440 16.440 ;
        RECT 28.520 16.120 28.840 16.440 ;
        RECT 28.920 16.120 29.240 16.440 ;
        RECT 73.160 16.120 73.480 16.440 ;
        RECT 73.560 16.120 73.880 16.440 ;
        RECT 73.960 16.120 74.280 16.440 ;
        RECT 74.360 16.120 74.680 16.440 ;
        RECT 118.600 16.120 118.920 16.440 ;
        RECT 119.000 16.120 119.320 16.440 ;
        RECT 119.400 16.120 119.720 16.440 ;
        RECT 119.800 16.120 120.120 16.440 ;
      LAYER met4 ;
        RECT 27.680 16.020 29.280 150.850 ;
        RECT 73.120 16.020 74.720 150.850 ;
        RECT 118.560 16.020 120.160 150.850 ;
      LAYER M4M5_PR_C ;
        RECT 27.890 127.360 29.070 128.540 ;
        RECT 27.890 82.590 29.070 83.770 ;
        RECT 27.890 37.820 29.070 39.000 ;
        RECT 73.330 127.360 74.510 128.540 ;
        RECT 73.330 82.590 74.510 83.770 ;
        RECT 73.330 37.820 74.510 39.000 ;
        RECT 118.770 127.360 119.950 128.540 ;
        RECT 118.770 82.590 119.950 83.770 ;
        RECT 118.770 37.820 119.950 39.000 ;
      LAYER met5 ;
        RECT 5.760 127.150 142.080 128.750 ;
        RECT 5.760 82.380 142.080 83.980 ;
        RECT 5.760 37.610 142.080 39.210 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    PORT
      LAYER li1 ;
        RECT 5.920 150.500 6.090 150.680 ;
        RECT 6.400 150.500 6.570 150.680 ;
        RECT 6.880 150.500 7.050 150.680 ;
        RECT 7.360 150.500 7.530 150.680 ;
        RECT 7.840 150.500 8.010 150.680 ;
        RECT 8.320 150.500 8.490 150.680 ;
        RECT 8.800 150.500 8.970 150.680 ;
        RECT 9.280 150.500 9.450 150.680 ;
        RECT 9.760 150.500 9.930 150.680 ;
        RECT 10.240 150.500 10.410 150.680 ;
        RECT 10.720 150.500 10.890 150.680 ;
        RECT 11.200 150.500 11.370 150.680 ;
        RECT 11.680 150.500 11.850 150.680 ;
        RECT 12.160 150.500 12.330 150.680 ;
        RECT 12.640 150.500 12.810 150.680 ;
        RECT 13.120 150.500 13.290 150.680 ;
        RECT 13.600 150.500 13.770 150.680 ;
        RECT 14.080 150.500 14.250 150.680 ;
        RECT 14.560 150.500 14.730 150.680 ;
        RECT 15.040 150.500 15.210 150.680 ;
        RECT 15.520 150.500 15.690 150.680 ;
        RECT 16.000 150.500 16.170 150.680 ;
        RECT 16.480 150.500 16.650 150.680 ;
        RECT 16.960 150.500 17.130 150.680 ;
        RECT 17.440 150.500 17.610 150.680 ;
        RECT 17.920 150.500 18.090 150.680 ;
        RECT 18.400 150.500 18.570 150.680 ;
        RECT 18.880 150.500 19.050 150.680 ;
        RECT 19.360 150.500 19.530 150.680 ;
        RECT 19.840 150.500 20.010 150.680 ;
        RECT 20.320 150.500 20.490 150.680 ;
        RECT 20.800 150.500 20.970 150.680 ;
        RECT 21.280 150.500 21.450 150.680 ;
        RECT 21.760 150.500 21.930 150.680 ;
        RECT 22.240 150.500 22.410 150.680 ;
        RECT 22.720 150.500 22.890 150.680 ;
        RECT 23.200 150.500 23.370 150.680 ;
        RECT 23.680 150.500 23.850 150.680 ;
        RECT 24.160 150.500 24.330 150.680 ;
        RECT 24.640 150.500 24.810 150.680 ;
        RECT 25.120 150.500 25.290 150.680 ;
        RECT 25.600 150.500 25.770 150.680 ;
        RECT 26.080 150.500 26.250 150.680 ;
        RECT 26.560 150.500 26.730 150.680 ;
        RECT 27.040 150.500 27.210 150.680 ;
        RECT 27.520 150.500 27.690 150.680 ;
        RECT 28.000 150.500 28.170 150.680 ;
        RECT 28.480 150.500 28.650 150.680 ;
        RECT 28.960 150.500 29.130 150.680 ;
        RECT 29.440 150.500 29.610 150.680 ;
        RECT 29.920 150.500 30.090 150.680 ;
        RECT 30.400 150.500 30.570 150.680 ;
        RECT 30.880 150.500 31.050 150.680 ;
        RECT 31.360 150.500 31.530 150.680 ;
        RECT 31.840 150.500 32.010 150.680 ;
        RECT 32.320 150.500 32.490 150.680 ;
        RECT 32.800 150.500 32.970 150.680 ;
        RECT 33.280 150.500 33.450 150.680 ;
        RECT 33.760 150.500 33.930 150.680 ;
        RECT 34.240 150.500 34.410 150.680 ;
        RECT 34.720 150.500 34.890 150.680 ;
        RECT 35.200 150.500 35.370 150.680 ;
        RECT 35.680 150.500 35.850 150.680 ;
        RECT 36.160 150.500 36.330 150.680 ;
        RECT 36.640 150.500 36.810 150.680 ;
        RECT 37.120 150.500 37.290 150.680 ;
        RECT 37.600 150.500 37.770 150.680 ;
        RECT 38.080 150.500 38.250 150.680 ;
        RECT 38.560 150.500 38.730 150.680 ;
        RECT 39.040 150.500 39.210 150.680 ;
        RECT 39.520 150.500 39.690 150.680 ;
        RECT 40.000 150.500 40.170 150.680 ;
        RECT 40.480 150.500 40.650 150.680 ;
        RECT 40.960 150.500 41.130 150.680 ;
        RECT 41.440 150.500 41.610 150.680 ;
        RECT 41.920 150.500 42.090 150.680 ;
        RECT 42.400 150.500 42.570 150.680 ;
        RECT 42.880 150.500 43.050 150.680 ;
        RECT 43.360 150.500 43.530 150.680 ;
        RECT 43.840 150.500 44.010 150.680 ;
        RECT 44.320 150.500 44.490 150.680 ;
        RECT 44.800 150.500 44.970 150.680 ;
        RECT 45.280 150.500 45.450 150.680 ;
        RECT 45.760 150.500 45.930 150.680 ;
        RECT 46.240 150.500 46.410 150.680 ;
        RECT 46.720 150.500 46.890 150.680 ;
        RECT 47.200 150.500 47.370 150.680 ;
        RECT 47.680 150.500 47.850 150.680 ;
        RECT 48.160 150.500 48.330 150.680 ;
        RECT 48.640 150.500 48.810 150.680 ;
        RECT 49.120 150.500 49.290 150.680 ;
        RECT 49.600 150.500 49.770 150.680 ;
        RECT 50.080 150.500 50.250 150.680 ;
        RECT 50.560 150.500 50.730 150.680 ;
        RECT 51.040 150.500 51.210 150.680 ;
        RECT 51.520 150.500 51.690 150.680 ;
        RECT 52.000 150.500 52.170 150.680 ;
        RECT 52.480 150.500 52.650 150.680 ;
        RECT 52.960 150.500 53.130 150.680 ;
        RECT 53.440 150.500 53.610 150.680 ;
        RECT 53.920 150.500 54.090 150.680 ;
        RECT 54.400 150.500 54.570 150.680 ;
        RECT 54.880 150.500 55.050 150.680 ;
        RECT 55.360 150.500 55.530 150.680 ;
        RECT 55.840 150.500 56.010 150.680 ;
        RECT 56.320 150.500 56.490 150.680 ;
        RECT 56.800 150.500 56.970 150.680 ;
        RECT 57.280 150.500 57.450 150.680 ;
        RECT 57.760 150.500 57.930 150.680 ;
        RECT 58.240 150.500 58.410 150.680 ;
        RECT 58.720 150.500 58.890 150.680 ;
        RECT 59.200 150.500 59.370 150.680 ;
        RECT 59.680 150.500 59.850 150.680 ;
        RECT 60.160 150.500 60.330 150.680 ;
        RECT 60.640 150.500 60.810 150.680 ;
        RECT 61.120 150.500 61.290 150.680 ;
        RECT 61.600 150.500 61.770 150.680 ;
        RECT 62.080 150.500 62.250 150.680 ;
        RECT 62.560 150.500 62.730 150.680 ;
        RECT 63.040 150.500 63.210 150.680 ;
        RECT 63.520 150.500 63.690 150.680 ;
        RECT 64.000 150.500 64.170 150.680 ;
        RECT 64.480 150.500 64.650 150.680 ;
        RECT 64.960 150.500 65.130 150.680 ;
        RECT 65.440 150.500 65.610 150.680 ;
        RECT 65.920 150.500 66.090 150.680 ;
        RECT 66.400 150.500 66.570 150.680 ;
        RECT 66.880 150.500 67.050 150.680 ;
        RECT 67.360 150.500 67.530 150.680 ;
        RECT 67.840 150.500 68.010 150.680 ;
        RECT 68.320 150.500 68.490 150.680 ;
        RECT 68.800 150.500 68.970 150.680 ;
        RECT 69.280 150.500 69.450 150.680 ;
        RECT 69.760 150.500 69.930 150.680 ;
        RECT 70.240 150.500 70.410 150.680 ;
        RECT 70.720 150.500 70.890 150.680 ;
        RECT 71.200 150.500 71.370 150.680 ;
        RECT 71.680 150.500 71.850 150.680 ;
        RECT 72.160 150.500 72.330 150.680 ;
        RECT 72.640 150.500 72.810 150.680 ;
        RECT 73.120 150.500 73.290 150.680 ;
        RECT 73.600 150.500 73.770 150.680 ;
        RECT 74.080 150.500 74.250 150.680 ;
        RECT 74.560 150.500 74.730 150.680 ;
        RECT 75.040 150.500 75.210 150.680 ;
        RECT 75.520 150.500 75.690 150.680 ;
        RECT 76.000 150.500 76.170 150.680 ;
        RECT 76.480 150.500 76.650 150.680 ;
        RECT 76.960 150.500 77.130 150.680 ;
        RECT 77.440 150.500 77.610 150.680 ;
        RECT 77.920 150.500 78.090 150.680 ;
        RECT 78.400 150.500 78.570 150.680 ;
        RECT 78.880 150.500 79.050 150.680 ;
        RECT 79.360 150.500 79.530 150.680 ;
        RECT 79.840 150.500 80.010 150.680 ;
        RECT 80.320 150.500 80.490 150.680 ;
        RECT 80.800 150.500 80.970 150.680 ;
        RECT 81.280 150.500 81.450 150.680 ;
        RECT 81.760 150.500 81.930 150.680 ;
        RECT 82.240 150.500 82.410 150.680 ;
        RECT 82.720 150.500 82.890 150.680 ;
        RECT 83.200 150.500 83.370 150.680 ;
        RECT 83.680 150.500 83.850 150.680 ;
        RECT 84.160 150.500 84.330 150.680 ;
        RECT 84.640 150.500 84.810 150.680 ;
        RECT 85.120 150.500 85.290 150.680 ;
        RECT 85.600 150.500 85.770 150.680 ;
        RECT 86.080 150.500 86.250 150.680 ;
        RECT 86.560 150.500 86.730 150.680 ;
        RECT 87.040 150.500 87.210 150.680 ;
        RECT 87.520 150.500 87.690 150.680 ;
        RECT 88.000 150.500 88.170 150.680 ;
        RECT 88.480 150.500 88.650 150.680 ;
        RECT 88.960 150.500 89.130 150.680 ;
        RECT 89.440 150.500 89.610 150.680 ;
        RECT 89.920 150.500 90.090 150.680 ;
        RECT 90.400 150.500 90.570 150.680 ;
        RECT 90.880 150.500 91.050 150.680 ;
        RECT 91.360 150.500 91.530 150.680 ;
        RECT 91.840 150.500 92.010 150.680 ;
        RECT 92.320 150.500 92.490 150.680 ;
        RECT 92.800 150.500 92.970 150.680 ;
        RECT 93.280 150.500 93.450 150.680 ;
        RECT 93.760 150.500 93.930 150.680 ;
        RECT 94.240 150.500 94.410 150.680 ;
        RECT 94.720 150.500 94.890 150.680 ;
        RECT 95.200 150.500 95.370 150.680 ;
        RECT 95.680 150.500 95.850 150.680 ;
        RECT 96.160 150.500 96.330 150.680 ;
        RECT 96.640 150.500 96.810 150.680 ;
        RECT 97.120 150.500 97.290 150.680 ;
        RECT 97.600 150.500 97.770 150.680 ;
        RECT 98.080 150.500 98.250 150.680 ;
        RECT 98.560 150.500 98.730 150.680 ;
        RECT 99.040 150.500 99.210 150.680 ;
        RECT 99.520 150.500 99.690 150.680 ;
        RECT 100.000 150.500 100.170 150.680 ;
        RECT 100.480 150.500 100.650 150.680 ;
        RECT 100.960 150.500 101.130 150.680 ;
        RECT 101.440 150.500 101.610 150.680 ;
        RECT 101.920 150.500 102.090 150.680 ;
        RECT 102.400 150.500 102.570 150.680 ;
        RECT 102.880 150.500 103.050 150.680 ;
        RECT 103.360 150.500 103.530 150.680 ;
        RECT 103.840 150.500 104.010 150.680 ;
        RECT 104.320 150.500 104.490 150.680 ;
        RECT 104.800 150.500 104.970 150.680 ;
        RECT 105.280 150.500 105.450 150.680 ;
        RECT 105.760 150.500 105.930 150.680 ;
        RECT 106.240 150.500 106.410 150.680 ;
        RECT 106.720 150.500 106.890 150.680 ;
        RECT 107.200 150.500 107.370 150.680 ;
        RECT 107.680 150.500 107.850 150.680 ;
        RECT 108.160 150.500 108.330 150.680 ;
        RECT 108.640 150.500 108.810 150.680 ;
        RECT 109.120 150.500 109.290 150.680 ;
        RECT 109.600 150.500 109.770 150.680 ;
        RECT 110.080 150.500 110.250 150.680 ;
        RECT 110.560 150.500 110.730 150.680 ;
        RECT 111.040 150.500 111.210 150.680 ;
        RECT 111.520 150.500 111.690 150.680 ;
        RECT 112.000 150.500 112.170 150.680 ;
        RECT 112.480 150.500 112.650 150.680 ;
        RECT 112.960 150.500 113.130 150.680 ;
        RECT 113.440 150.500 113.610 150.680 ;
        RECT 113.920 150.500 114.090 150.680 ;
        RECT 114.400 150.500 114.570 150.680 ;
        RECT 114.880 150.500 115.050 150.680 ;
        RECT 115.360 150.500 115.530 150.680 ;
        RECT 115.840 150.500 116.010 150.680 ;
        RECT 116.320 150.500 116.490 150.680 ;
        RECT 116.800 150.500 116.970 150.680 ;
        RECT 117.280 150.500 117.450 150.680 ;
        RECT 117.760 150.500 117.930 150.680 ;
        RECT 118.240 150.500 118.410 150.680 ;
        RECT 118.720 150.500 118.890 150.680 ;
        RECT 119.200 150.500 119.370 150.680 ;
        RECT 119.680 150.500 119.850 150.680 ;
        RECT 120.160 150.500 120.330 150.680 ;
        RECT 120.640 150.500 120.810 150.680 ;
        RECT 121.120 150.500 121.290 150.680 ;
        RECT 121.600 150.500 121.770 150.680 ;
        RECT 122.080 150.500 122.250 150.680 ;
        RECT 122.560 150.500 122.730 150.680 ;
        RECT 123.040 150.500 123.210 150.680 ;
        RECT 123.520 150.500 123.690 150.680 ;
        RECT 124.000 150.500 124.170 150.680 ;
        RECT 124.480 150.500 124.650 150.680 ;
        RECT 124.960 150.500 125.130 150.680 ;
        RECT 125.440 150.500 125.610 150.680 ;
        RECT 125.920 150.500 126.090 150.680 ;
        RECT 126.400 150.500 126.570 150.680 ;
        RECT 126.880 150.500 127.050 150.680 ;
        RECT 127.360 150.500 127.530 150.680 ;
        RECT 127.840 150.500 128.010 150.680 ;
        RECT 128.320 150.500 128.490 150.680 ;
        RECT 128.800 150.500 128.970 150.680 ;
        RECT 129.280 150.500 129.450 150.680 ;
        RECT 129.760 150.500 129.930 150.680 ;
        RECT 130.240 150.500 130.410 150.680 ;
        RECT 130.720 150.500 130.890 150.680 ;
        RECT 131.200 150.500 131.370 150.680 ;
        RECT 131.680 150.500 131.850 150.680 ;
        RECT 132.160 150.500 132.330 150.680 ;
        RECT 132.640 150.500 132.810 150.680 ;
        RECT 133.120 150.500 133.290 150.680 ;
        RECT 133.600 150.500 133.770 150.680 ;
        RECT 134.080 150.500 134.250 150.680 ;
        RECT 134.560 150.500 134.730 150.680 ;
        RECT 135.040 150.500 135.210 150.680 ;
        RECT 135.520 150.500 135.690 150.680 ;
        RECT 136.000 150.500 136.170 150.680 ;
        RECT 136.480 150.500 136.650 150.680 ;
        RECT 136.960 150.500 137.130 150.680 ;
        RECT 137.440 150.500 137.610 150.680 ;
        RECT 137.920 150.500 138.090 150.680 ;
        RECT 138.400 150.500 138.570 150.680 ;
        RECT 138.880 150.500 139.050 150.680 ;
        RECT 139.360 150.500 139.530 150.680 ;
        RECT 139.840 150.500 140.010 150.680 ;
        RECT 140.320 150.500 140.490 150.680 ;
        RECT 140.800 150.500 140.970 150.680 ;
        RECT 141.280 150.500 141.450 150.680 ;
      LAYER li1 ;
        RECT 141.600 150.500 142.080 150.680 ;
      LAYER li1 ;
        RECT 6.510 150.030 6.680 150.200 ;
        RECT 6.950 150.030 7.120 150.200 ;
        RECT 7.360 150.030 7.530 150.200 ;
        RECT 7.790 150.030 7.960 150.200 ;
        RECT 8.230 150.030 8.400 150.200 ;
        RECT 8.640 150.030 8.810 150.200 ;
        RECT 10.350 150.030 10.520 150.200 ;
        RECT 10.790 150.030 10.960 150.200 ;
        RECT 11.200 150.030 11.370 150.200 ;
        RECT 11.630 150.030 11.800 150.200 ;
        RECT 12.070 150.030 12.240 150.200 ;
        RECT 12.480 150.030 12.650 150.200 ;
        RECT 14.190 150.030 14.360 150.200 ;
        RECT 14.630 150.030 14.800 150.200 ;
        RECT 15.040 150.030 15.210 150.200 ;
        RECT 15.470 150.030 15.640 150.200 ;
        RECT 15.910 150.030 16.080 150.200 ;
        RECT 16.320 150.030 16.490 150.200 ;
        RECT 18.030 150.030 18.200 150.200 ;
        RECT 18.470 150.030 18.640 150.200 ;
        RECT 18.880 150.030 19.050 150.200 ;
        RECT 19.310 150.030 19.480 150.200 ;
        RECT 19.750 150.030 19.920 150.200 ;
        RECT 20.160 150.030 20.330 150.200 ;
        RECT 23.680 150.020 23.850 150.190 ;
        RECT 24.040 150.020 24.210 150.190 ;
        RECT 25.230 150.030 25.400 150.200 ;
        RECT 25.670 150.030 25.840 150.200 ;
        RECT 26.080 150.030 26.250 150.200 ;
        RECT 26.510 150.030 26.680 150.200 ;
        RECT 26.950 150.030 27.120 150.200 ;
        RECT 27.360 150.030 27.530 150.200 ;
        RECT 29.070 150.030 29.240 150.200 ;
        RECT 29.510 150.030 29.680 150.200 ;
        RECT 29.920 150.030 30.090 150.200 ;
        RECT 30.350 150.030 30.520 150.200 ;
        RECT 30.790 150.030 30.960 150.200 ;
        RECT 31.200 150.030 31.370 150.200 ;
        RECT 32.910 150.030 33.080 150.200 ;
        RECT 33.350 150.030 33.520 150.200 ;
        RECT 33.760 150.030 33.930 150.200 ;
        RECT 34.190 150.030 34.360 150.200 ;
        RECT 34.630 150.030 34.800 150.200 ;
        RECT 35.040 150.030 35.210 150.200 ;
        RECT 36.750 150.030 36.920 150.200 ;
        RECT 37.190 150.030 37.360 150.200 ;
        RECT 37.600 150.030 37.770 150.200 ;
        RECT 38.030 150.030 38.200 150.200 ;
        RECT 38.470 150.030 38.640 150.200 ;
        RECT 38.880 150.030 39.050 150.200 ;
        RECT 40.590 150.030 40.760 150.200 ;
        RECT 41.030 150.030 41.200 150.200 ;
        RECT 41.440 150.030 41.610 150.200 ;
        RECT 41.870 150.030 42.040 150.200 ;
        RECT 42.310 150.030 42.480 150.200 ;
        RECT 42.720 150.030 42.890 150.200 ;
        RECT 44.430 150.030 44.600 150.200 ;
        RECT 44.870 150.030 45.040 150.200 ;
        RECT 45.280 150.030 45.450 150.200 ;
        RECT 45.710 150.030 45.880 150.200 ;
        RECT 46.150 150.030 46.320 150.200 ;
        RECT 46.560 150.030 46.730 150.200 ;
        RECT 48.270 150.030 48.440 150.200 ;
        RECT 48.710 150.030 48.880 150.200 ;
        RECT 49.120 150.030 49.290 150.200 ;
        RECT 49.550 150.030 49.720 150.200 ;
        RECT 49.990 150.030 50.160 150.200 ;
        RECT 50.400 150.030 50.570 150.200 ;
        RECT 52.110 150.030 52.280 150.200 ;
        RECT 52.550 150.030 52.720 150.200 ;
        RECT 52.960 150.030 53.130 150.200 ;
        RECT 53.390 150.030 53.560 150.200 ;
        RECT 53.830 150.030 54.000 150.200 ;
        RECT 54.240 150.030 54.410 150.200 ;
        RECT 55.950 150.030 56.120 150.200 ;
        RECT 56.390 150.030 56.560 150.200 ;
        RECT 56.800 150.030 56.970 150.200 ;
        RECT 57.230 150.030 57.400 150.200 ;
        RECT 57.670 150.030 57.840 150.200 ;
        RECT 58.080 150.030 58.250 150.200 ;
        RECT 59.790 150.030 59.960 150.200 ;
        RECT 60.230 150.030 60.400 150.200 ;
        RECT 60.640 150.030 60.810 150.200 ;
        RECT 61.070 150.030 61.240 150.200 ;
        RECT 61.510 150.030 61.680 150.200 ;
        RECT 61.920 150.030 62.090 150.200 ;
        RECT 63.100 150.020 63.270 150.190 ;
        RECT 63.540 150.020 63.710 150.190 ;
        RECT 63.980 150.020 64.150 150.190 ;
        RECT 64.390 150.020 64.560 150.190 ;
        RECT 66.400 150.020 66.570 150.190 ;
        RECT 66.760 150.020 66.930 150.190 ;
        RECT 67.950 150.030 68.120 150.200 ;
        RECT 68.390 150.030 68.560 150.200 ;
        RECT 68.800 150.030 68.970 150.200 ;
        RECT 69.230 150.030 69.400 150.200 ;
        RECT 69.670 150.030 69.840 150.200 ;
        RECT 70.080 150.030 70.250 150.200 ;
        RECT 71.790 150.030 71.960 150.200 ;
        RECT 72.230 150.030 72.400 150.200 ;
        RECT 72.640 150.030 72.810 150.200 ;
        RECT 73.070 150.030 73.240 150.200 ;
        RECT 73.510 150.030 73.680 150.200 ;
        RECT 73.920 150.030 74.090 150.200 ;
        RECT 76.480 150.020 76.650 150.190 ;
        RECT 76.840 150.020 77.010 150.190 ;
        RECT 78.030 150.030 78.200 150.200 ;
        RECT 78.470 150.030 78.640 150.200 ;
        RECT 78.880 150.030 79.050 150.200 ;
        RECT 79.310 150.030 79.480 150.200 ;
        RECT 79.750 150.030 79.920 150.200 ;
        RECT 80.160 150.030 80.330 150.200 ;
        RECT 81.870 150.030 82.040 150.200 ;
        RECT 82.310 150.030 82.480 150.200 ;
        RECT 82.720 150.030 82.890 150.200 ;
        RECT 83.150 150.030 83.320 150.200 ;
        RECT 83.590 150.030 83.760 150.200 ;
        RECT 84.000 150.030 84.170 150.200 ;
        RECT 85.710 150.030 85.880 150.200 ;
        RECT 86.150 150.030 86.320 150.200 ;
        RECT 86.560 150.030 86.730 150.200 ;
        RECT 86.990 150.030 87.160 150.200 ;
        RECT 87.430 150.030 87.600 150.200 ;
        RECT 87.840 150.030 88.010 150.200 ;
        RECT 89.550 150.030 89.720 150.200 ;
        RECT 89.990 150.030 90.160 150.200 ;
        RECT 90.400 150.030 90.570 150.200 ;
        RECT 90.830 150.030 91.000 150.200 ;
        RECT 91.270 150.030 91.440 150.200 ;
        RECT 91.680 150.030 91.850 150.200 ;
        RECT 93.390 150.030 93.560 150.200 ;
        RECT 93.830 150.030 94.000 150.200 ;
        RECT 94.240 150.030 94.410 150.200 ;
        RECT 94.670 150.030 94.840 150.200 ;
        RECT 95.110 150.030 95.280 150.200 ;
        RECT 95.520 150.030 95.690 150.200 ;
        RECT 97.230 150.030 97.400 150.200 ;
        RECT 97.670 150.030 97.840 150.200 ;
        RECT 98.080 150.030 98.250 150.200 ;
        RECT 98.510 150.030 98.680 150.200 ;
        RECT 98.950 150.030 99.120 150.200 ;
        RECT 99.360 150.030 99.530 150.200 ;
        RECT 101.070 150.030 101.240 150.200 ;
        RECT 101.510 150.030 101.680 150.200 ;
        RECT 101.920 150.030 102.090 150.200 ;
        RECT 102.350 150.030 102.520 150.200 ;
        RECT 102.790 150.030 102.960 150.200 ;
        RECT 103.200 150.030 103.370 150.200 ;
        RECT 104.910 150.030 105.080 150.200 ;
        RECT 105.350 150.030 105.520 150.200 ;
        RECT 105.760 150.030 105.930 150.200 ;
        RECT 106.190 150.030 106.360 150.200 ;
        RECT 106.630 150.030 106.800 150.200 ;
        RECT 107.040 150.030 107.210 150.200 ;
        RECT 108.750 150.030 108.920 150.200 ;
        RECT 109.190 150.030 109.360 150.200 ;
        RECT 109.600 150.030 109.770 150.200 ;
        RECT 110.030 150.030 110.200 150.200 ;
        RECT 110.470 150.030 110.640 150.200 ;
        RECT 110.880 150.030 111.050 150.200 ;
        RECT 112.590 150.030 112.760 150.200 ;
        RECT 113.030 150.030 113.200 150.200 ;
        RECT 113.440 150.030 113.610 150.200 ;
        RECT 113.870 150.030 114.040 150.200 ;
        RECT 114.310 150.030 114.480 150.200 ;
        RECT 114.720 150.030 114.890 150.200 ;
        RECT 116.430 150.030 116.600 150.200 ;
        RECT 116.870 150.030 117.040 150.200 ;
        RECT 117.280 150.030 117.450 150.200 ;
        RECT 117.710 150.030 117.880 150.200 ;
        RECT 118.150 150.030 118.320 150.200 ;
        RECT 118.560 150.030 118.730 150.200 ;
        RECT 120.270 150.030 120.440 150.200 ;
        RECT 120.710 150.030 120.880 150.200 ;
        RECT 121.120 150.030 121.290 150.200 ;
        RECT 121.550 150.030 121.720 150.200 ;
        RECT 121.990 150.030 122.160 150.200 ;
        RECT 122.400 150.030 122.570 150.200 ;
        RECT 124.110 150.030 124.280 150.200 ;
        RECT 124.550 150.030 124.720 150.200 ;
        RECT 124.960 150.030 125.130 150.200 ;
        RECT 125.390 150.030 125.560 150.200 ;
        RECT 125.830 150.030 126.000 150.200 ;
        RECT 126.240 150.030 126.410 150.200 ;
        RECT 127.950 150.030 128.120 150.200 ;
        RECT 128.390 150.030 128.560 150.200 ;
        RECT 128.800 150.030 128.970 150.200 ;
        RECT 129.230 150.030 129.400 150.200 ;
        RECT 129.670 150.030 129.840 150.200 ;
        RECT 130.080 150.030 130.250 150.200 ;
        RECT 131.790 150.030 131.960 150.200 ;
        RECT 132.230 150.030 132.400 150.200 ;
        RECT 132.640 150.030 132.810 150.200 ;
        RECT 133.070 150.030 133.240 150.200 ;
        RECT 133.510 150.030 133.680 150.200 ;
        RECT 133.920 150.030 134.090 150.200 ;
        RECT 135.630 150.030 135.800 150.200 ;
        RECT 136.070 150.030 136.240 150.200 ;
        RECT 136.480 150.030 136.650 150.200 ;
        RECT 136.910 150.030 137.080 150.200 ;
        RECT 137.350 150.030 137.520 150.200 ;
        RECT 137.760 150.030 137.930 150.200 ;
        RECT 138.940 150.020 139.110 150.190 ;
        RECT 139.380 150.020 139.550 150.190 ;
        RECT 139.820 150.020 139.990 150.190 ;
        RECT 140.230 150.020 140.400 150.190 ;
        RECT 5.920 142.360 6.090 142.540 ;
        RECT 6.400 142.360 6.570 142.540 ;
        RECT 6.880 142.360 7.050 142.540 ;
        RECT 7.360 142.360 7.530 142.540 ;
        RECT 7.840 142.360 8.010 142.540 ;
        RECT 8.320 142.360 8.490 142.540 ;
        RECT 8.800 142.360 8.970 142.540 ;
        RECT 9.280 142.360 9.450 142.540 ;
        RECT 9.760 142.360 9.930 142.540 ;
        RECT 10.240 142.360 10.410 142.540 ;
        RECT 10.720 142.360 10.890 142.540 ;
        RECT 11.200 142.360 11.370 142.540 ;
        RECT 11.680 142.360 11.850 142.540 ;
        RECT 12.160 142.360 12.330 142.540 ;
        RECT 12.640 142.360 12.810 142.540 ;
        RECT 13.120 142.360 13.290 142.540 ;
        RECT 13.600 142.360 13.770 142.540 ;
        RECT 14.080 142.360 14.250 142.540 ;
        RECT 14.560 142.360 14.730 142.540 ;
        RECT 15.040 142.360 15.210 142.540 ;
        RECT 15.520 142.360 15.690 142.540 ;
        RECT 16.000 142.360 16.170 142.540 ;
        RECT 16.480 142.360 16.650 142.540 ;
        RECT 16.960 142.360 17.130 142.540 ;
        RECT 17.440 142.360 17.610 142.540 ;
      LAYER li1 ;
        RECT 17.760 142.360 18.240 142.540 ;
      LAYER li1 ;
        RECT 18.400 142.360 18.570 142.540 ;
        RECT 18.880 142.360 19.050 142.540 ;
        RECT 19.360 142.360 19.530 142.540 ;
        RECT 19.840 142.360 20.010 142.540 ;
        RECT 20.320 142.360 20.490 142.540 ;
        RECT 20.800 142.360 20.970 142.540 ;
        RECT 21.280 142.360 21.450 142.540 ;
        RECT 21.760 142.360 21.930 142.540 ;
        RECT 22.240 142.360 22.410 142.540 ;
        RECT 22.720 142.360 22.890 142.540 ;
        RECT 23.200 142.360 23.370 142.540 ;
        RECT 23.680 142.360 23.850 142.540 ;
        RECT 24.160 142.360 24.330 142.540 ;
        RECT 24.640 142.360 24.810 142.540 ;
        RECT 25.120 142.360 25.290 142.540 ;
        RECT 25.600 142.360 25.770 142.540 ;
        RECT 26.080 142.360 26.250 142.540 ;
        RECT 26.560 142.360 26.730 142.540 ;
        RECT 27.040 142.360 27.210 142.540 ;
        RECT 27.520 142.360 27.690 142.540 ;
        RECT 28.000 142.360 28.170 142.540 ;
        RECT 28.480 142.360 28.650 142.540 ;
        RECT 28.960 142.360 29.130 142.540 ;
        RECT 29.440 142.360 29.610 142.540 ;
        RECT 29.920 142.360 30.090 142.540 ;
        RECT 30.400 142.360 30.570 142.540 ;
        RECT 30.880 142.360 31.050 142.540 ;
        RECT 31.360 142.360 31.530 142.540 ;
        RECT 31.840 142.360 32.010 142.540 ;
        RECT 32.320 142.360 32.490 142.540 ;
        RECT 32.800 142.360 32.970 142.540 ;
        RECT 33.280 142.360 33.450 142.540 ;
        RECT 33.760 142.360 33.930 142.540 ;
        RECT 34.240 142.360 34.410 142.540 ;
        RECT 34.720 142.360 34.890 142.540 ;
        RECT 35.200 142.360 35.370 142.540 ;
        RECT 35.680 142.360 35.850 142.540 ;
      LAYER li1 ;
        RECT 36.000 142.360 36.480 142.540 ;
      LAYER li1 ;
        RECT 36.640 142.360 36.810 142.540 ;
        RECT 37.120 142.360 37.290 142.540 ;
        RECT 37.600 142.360 37.770 142.540 ;
        RECT 38.080 142.360 38.250 142.540 ;
        RECT 38.560 142.360 38.730 142.540 ;
        RECT 39.040 142.360 39.210 142.540 ;
        RECT 39.520 142.360 39.690 142.540 ;
        RECT 40.000 142.360 40.170 142.540 ;
        RECT 40.480 142.360 40.650 142.540 ;
        RECT 40.960 142.360 41.130 142.540 ;
        RECT 41.440 142.360 41.610 142.540 ;
        RECT 41.920 142.360 42.090 142.540 ;
        RECT 42.400 142.360 42.570 142.540 ;
        RECT 42.880 142.360 43.050 142.540 ;
        RECT 43.360 142.360 43.530 142.540 ;
      LAYER li1 ;
        RECT 43.680 142.360 44.160 142.540 ;
      LAYER li1 ;
        RECT 44.320 142.360 44.490 142.540 ;
        RECT 44.800 142.360 44.970 142.540 ;
        RECT 45.280 142.360 45.450 142.540 ;
        RECT 45.760 142.360 45.930 142.540 ;
        RECT 46.240 142.360 46.410 142.540 ;
        RECT 46.720 142.360 46.890 142.540 ;
        RECT 47.200 142.360 47.370 142.540 ;
        RECT 47.680 142.360 47.850 142.540 ;
        RECT 48.160 142.360 48.330 142.540 ;
        RECT 48.640 142.360 48.810 142.540 ;
        RECT 49.120 142.360 49.290 142.540 ;
        RECT 49.600 142.360 49.770 142.540 ;
        RECT 50.080 142.360 50.250 142.540 ;
        RECT 50.560 142.360 50.730 142.540 ;
        RECT 51.040 142.360 51.210 142.540 ;
        RECT 51.520 142.360 51.690 142.540 ;
        RECT 52.000 142.360 52.170 142.540 ;
        RECT 52.480 142.360 52.650 142.540 ;
        RECT 52.960 142.360 53.130 142.540 ;
        RECT 53.440 142.360 53.610 142.540 ;
        RECT 53.920 142.360 54.090 142.540 ;
        RECT 54.400 142.360 54.570 142.540 ;
        RECT 54.880 142.360 55.050 142.540 ;
        RECT 55.360 142.360 55.530 142.540 ;
        RECT 55.840 142.360 56.010 142.540 ;
        RECT 56.320 142.360 56.490 142.540 ;
        RECT 56.800 142.360 56.970 142.540 ;
        RECT 57.280 142.360 57.450 142.540 ;
        RECT 57.760 142.360 57.930 142.540 ;
        RECT 58.240 142.360 58.410 142.540 ;
        RECT 58.720 142.360 58.890 142.540 ;
        RECT 59.200 142.360 59.370 142.540 ;
        RECT 59.680 142.360 59.850 142.540 ;
        RECT 60.160 142.360 60.330 142.540 ;
        RECT 60.640 142.360 60.810 142.540 ;
        RECT 61.120 142.360 61.290 142.540 ;
        RECT 61.600 142.360 61.770 142.540 ;
        RECT 62.080 142.360 62.250 142.540 ;
        RECT 62.560 142.360 62.730 142.540 ;
        RECT 63.040 142.360 63.210 142.540 ;
        RECT 63.520 142.360 63.690 142.540 ;
        RECT 64.000 142.360 64.170 142.540 ;
        RECT 64.480 142.360 64.650 142.540 ;
        RECT 64.960 142.360 65.130 142.540 ;
        RECT 65.440 142.360 65.610 142.540 ;
        RECT 65.920 142.360 66.090 142.540 ;
        RECT 66.400 142.360 66.570 142.540 ;
        RECT 66.880 142.360 67.050 142.540 ;
        RECT 67.360 142.360 67.530 142.540 ;
        RECT 67.840 142.360 68.010 142.540 ;
        RECT 68.320 142.360 68.490 142.540 ;
        RECT 68.800 142.360 68.970 142.540 ;
        RECT 69.280 142.360 69.450 142.540 ;
        RECT 69.760 142.360 69.930 142.540 ;
        RECT 70.240 142.360 70.410 142.540 ;
        RECT 70.720 142.360 70.890 142.540 ;
        RECT 71.200 142.360 71.370 142.540 ;
        RECT 71.680 142.360 71.850 142.540 ;
        RECT 72.160 142.360 72.330 142.540 ;
        RECT 72.640 142.360 72.810 142.540 ;
        RECT 73.120 142.360 73.290 142.540 ;
        RECT 73.600 142.360 73.770 142.540 ;
        RECT 74.080 142.360 74.250 142.540 ;
        RECT 74.560 142.360 74.730 142.540 ;
        RECT 75.040 142.360 75.210 142.540 ;
        RECT 75.520 142.360 75.690 142.540 ;
        RECT 76.000 142.360 76.170 142.540 ;
        RECT 76.480 142.360 76.650 142.540 ;
        RECT 76.960 142.360 77.130 142.540 ;
        RECT 77.440 142.360 77.610 142.540 ;
        RECT 77.920 142.360 78.090 142.540 ;
        RECT 78.400 142.360 78.570 142.540 ;
        RECT 78.880 142.360 79.050 142.540 ;
        RECT 79.360 142.360 79.530 142.540 ;
        RECT 79.840 142.360 80.010 142.540 ;
        RECT 80.320 142.360 80.490 142.540 ;
        RECT 80.800 142.360 80.970 142.540 ;
        RECT 81.280 142.360 81.450 142.540 ;
        RECT 81.760 142.360 81.930 142.540 ;
        RECT 82.240 142.360 82.410 142.540 ;
        RECT 82.720 142.360 82.890 142.540 ;
        RECT 83.200 142.360 83.370 142.540 ;
        RECT 83.680 142.360 83.850 142.540 ;
        RECT 84.160 142.360 84.330 142.540 ;
        RECT 84.640 142.360 84.810 142.540 ;
        RECT 85.120 142.360 85.290 142.540 ;
      LAYER li1 ;
        RECT 85.440 142.360 85.920 142.540 ;
      LAYER li1 ;
        RECT 86.080 142.360 86.250 142.540 ;
        RECT 86.560 142.360 86.730 142.540 ;
        RECT 87.040 142.360 87.210 142.540 ;
        RECT 87.520 142.360 87.690 142.540 ;
        RECT 88.000 142.360 88.170 142.540 ;
        RECT 88.480 142.360 88.650 142.540 ;
        RECT 88.960 142.360 89.130 142.540 ;
        RECT 89.440 142.360 89.610 142.540 ;
        RECT 89.920 142.360 90.090 142.540 ;
        RECT 90.400 142.360 90.570 142.540 ;
        RECT 90.880 142.360 91.050 142.540 ;
        RECT 91.360 142.360 91.530 142.540 ;
        RECT 91.840 142.360 92.010 142.540 ;
        RECT 92.320 142.360 92.490 142.540 ;
        RECT 92.800 142.360 92.970 142.540 ;
        RECT 93.280 142.360 93.450 142.540 ;
        RECT 93.760 142.360 93.930 142.540 ;
        RECT 94.240 142.360 94.410 142.540 ;
        RECT 94.720 142.360 94.890 142.540 ;
        RECT 95.200 142.360 95.370 142.540 ;
        RECT 95.680 142.360 95.850 142.540 ;
        RECT 96.160 142.360 96.330 142.540 ;
        RECT 96.640 142.360 96.810 142.540 ;
        RECT 97.120 142.360 97.290 142.540 ;
        RECT 97.600 142.360 97.770 142.540 ;
        RECT 98.080 142.360 98.250 142.540 ;
        RECT 98.560 142.360 98.730 142.540 ;
        RECT 99.040 142.360 99.210 142.540 ;
        RECT 99.520 142.360 99.690 142.540 ;
        RECT 100.000 142.360 100.170 142.540 ;
        RECT 100.480 142.360 100.650 142.540 ;
        RECT 100.960 142.360 101.130 142.540 ;
        RECT 101.440 142.360 101.610 142.540 ;
        RECT 101.920 142.360 102.090 142.540 ;
        RECT 102.400 142.360 102.570 142.540 ;
        RECT 102.880 142.360 103.050 142.540 ;
        RECT 103.360 142.360 103.530 142.540 ;
        RECT 103.840 142.360 104.010 142.540 ;
        RECT 104.320 142.360 104.490 142.540 ;
        RECT 104.800 142.360 104.970 142.540 ;
        RECT 105.280 142.360 105.450 142.540 ;
        RECT 105.760 142.360 105.930 142.540 ;
        RECT 106.240 142.360 106.410 142.540 ;
        RECT 106.720 142.360 106.890 142.540 ;
        RECT 107.200 142.360 107.370 142.540 ;
        RECT 107.680 142.360 107.850 142.540 ;
        RECT 108.160 142.360 108.330 142.540 ;
        RECT 108.640 142.360 108.810 142.540 ;
        RECT 109.120 142.360 109.290 142.540 ;
        RECT 109.600 142.360 109.770 142.540 ;
        RECT 110.080 142.360 110.250 142.540 ;
        RECT 110.560 142.360 110.730 142.540 ;
        RECT 111.040 142.360 111.210 142.540 ;
        RECT 111.520 142.360 111.690 142.540 ;
        RECT 112.000 142.360 112.170 142.540 ;
        RECT 112.480 142.360 112.650 142.540 ;
        RECT 112.960 142.360 113.130 142.540 ;
        RECT 113.440 142.360 113.610 142.540 ;
        RECT 113.920 142.360 114.090 142.540 ;
        RECT 114.400 142.360 114.570 142.540 ;
        RECT 114.880 142.360 115.050 142.540 ;
        RECT 115.360 142.360 115.530 142.540 ;
        RECT 115.840 142.360 116.010 142.540 ;
        RECT 116.320 142.360 116.490 142.540 ;
        RECT 116.800 142.360 116.970 142.540 ;
        RECT 117.280 142.360 117.450 142.540 ;
        RECT 117.760 142.360 117.930 142.540 ;
        RECT 118.240 142.360 118.410 142.540 ;
        RECT 118.720 142.360 118.890 142.540 ;
        RECT 119.200 142.360 119.370 142.540 ;
        RECT 119.680 142.360 119.850 142.540 ;
        RECT 120.160 142.360 120.330 142.540 ;
        RECT 120.640 142.360 120.810 142.540 ;
        RECT 121.120 142.360 121.290 142.540 ;
        RECT 121.600 142.360 121.770 142.540 ;
        RECT 122.080 142.360 122.250 142.540 ;
        RECT 122.560 142.360 122.730 142.540 ;
        RECT 123.040 142.360 123.210 142.540 ;
        RECT 123.520 142.360 123.690 142.540 ;
        RECT 124.000 142.360 124.170 142.540 ;
        RECT 124.480 142.360 124.650 142.540 ;
        RECT 124.960 142.360 125.130 142.540 ;
        RECT 125.440 142.360 125.610 142.540 ;
        RECT 125.920 142.360 126.090 142.540 ;
        RECT 126.400 142.360 126.570 142.540 ;
        RECT 126.880 142.360 127.050 142.540 ;
        RECT 127.360 142.360 127.530 142.540 ;
        RECT 127.840 142.360 128.010 142.540 ;
        RECT 128.320 142.360 128.490 142.540 ;
        RECT 128.800 142.360 128.970 142.540 ;
        RECT 129.280 142.360 129.450 142.540 ;
        RECT 129.760 142.360 129.930 142.540 ;
        RECT 130.240 142.360 130.410 142.540 ;
        RECT 130.720 142.360 130.890 142.540 ;
        RECT 131.200 142.360 131.370 142.540 ;
        RECT 131.680 142.360 131.850 142.540 ;
        RECT 132.160 142.360 132.330 142.540 ;
        RECT 132.640 142.360 132.810 142.540 ;
        RECT 133.120 142.360 133.290 142.540 ;
        RECT 133.600 142.360 133.770 142.540 ;
        RECT 134.080 142.360 134.250 142.540 ;
        RECT 134.560 142.360 134.730 142.540 ;
        RECT 135.040 142.360 135.210 142.540 ;
        RECT 135.520 142.360 135.690 142.540 ;
        RECT 136.000 142.360 136.170 142.540 ;
        RECT 136.480 142.360 136.650 142.540 ;
        RECT 136.960 142.360 137.130 142.540 ;
        RECT 137.440 142.360 137.610 142.540 ;
        RECT 137.920 142.360 138.090 142.540 ;
        RECT 138.400 142.360 138.570 142.540 ;
        RECT 138.880 142.360 139.050 142.540 ;
        RECT 139.360 142.360 139.530 142.540 ;
        RECT 139.840 142.360 140.010 142.540 ;
        RECT 140.320 142.360 140.490 142.540 ;
        RECT 140.800 142.360 140.970 142.540 ;
        RECT 141.280 142.360 141.450 142.540 ;
      LAYER li1 ;
        RECT 141.600 142.360 142.080 142.540 ;
      LAYER li1 ;
        RECT 6.510 141.890 6.680 142.060 ;
        RECT 6.950 141.890 7.120 142.060 ;
        RECT 7.360 141.890 7.530 142.060 ;
        RECT 7.790 141.890 7.960 142.060 ;
        RECT 8.230 141.890 8.400 142.060 ;
        RECT 8.640 141.890 8.810 142.060 ;
        RECT 10.350 141.890 10.520 142.060 ;
        RECT 10.790 141.890 10.960 142.060 ;
        RECT 11.200 141.890 11.370 142.060 ;
        RECT 11.630 141.890 11.800 142.060 ;
        RECT 12.070 141.890 12.240 142.060 ;
        RECT 12.480 141.890 12.650 142.060 ;
        RECT 14.190 141.890 14.360 142.060 ;
        RECT 14.630 141.890 14.800 142.060 ;
        RECT 15.040 141.890 15.210 142.060 ;
        RECT 15.470 141.890 15.640 142.060 ;
        RECT 15.910 141.890 16.080 142.060 ;
        RECT 16.320 141.890 16.490 142.060 ;
        RECT 18.030 141.890 18.200 142.060 ;
        RECT 18.470 141.890 18.640 142.060 ;
        RECT 18.880 141.890 19.050 142.060 ;
        RECT 19.310 141.890 19.480 142.060 ;
        RECT 19.750 141.890 19.920 142.060 ;
        RECT 20.160 141.890 20.330 142.060 ;
        RECT 21.870 141.890 22.040 142.060 ;
        RECT 22.310 141.890 22.480 142.060 ;
        RECT 22.720 141.890 22.890 142.060 ;
        RECT 23.150 141.890 23.320 142.060 ;
        RECT 23.590 141.890 23.760 142.060 ;
        RECT 24.000 141.890 24.170 142.060 ;
        RECT 25.710 141.890 25.880 142.060 ;
        RECT 26.150 141.890 26.320 142.060 ;
        RECT 26.560 141.890 26.730 142.060 ;
        RECT 26.990 141.890 27.160 142.060 ;
        RECT 27.430 141.890 27.600 142.060 ;
        RECT 27.840 141.890 28.010 142.060 ;
        RECT 30.830 141.880 31.000 142.050 ;
        RECT 31.190 141.880 31.360 142.050 ;
        RECT 31.550 141.880 31.720 142.050 ;
        RECT 32.470 141.880 32.640 142.050 ;
        RECT 32.830 141.880 33.000 142.050 ;
        RECT 37.430 141.880 37.600 142.050 ;
        RECT 37.790 141.880 37.960 142.050 ;
        RECT 38.150 141.880 38.320 142.050 ;
        RECT 41.400 141.880 41.570 142.050 ;
        RECT 41.760 141.880 41.930 142.050 ;
        RECT 42.120 141.880 42.290 142.050 ;
        RECT 44.010 141.880 44.180 142.050 ;
        RECT 44.370 141.880 44.540 142.050 ;
        RECT 44.730 141.880 44.900 142.050 ;
        RECT 45.820 141.880 45.990 142.050 ;
        RECT 46.260 141.880 46.430 142.050 ;
        RECT 46.700 141.880 46.870 142.050 ;
        RECT 47.110 141.880 47.280 142.050 ;
        RECT 48.110 141.880 48.280 142.050 ;
        RECT 48.470 141.880 48.640 142.050 ;
        RECT 48.830 141.880 49.000 142.050 ;
        RECT 49.750 141.880 49.920 142.050 ;
        RECT 50.110 141.880 50.280 142.050 ;
        RECT 54.710 141.880 54.880 142.050 ;
        RECT 55.070 141.880 55.240 142.050 ;
        RECT 55.430 141.880 55.600 142.050 ;
        RECT 58.680 141.880 58.850 142.050 ;
        RECT 59.040 141.880 59.210 142.050 ;
        RECT 59.400 141.880 59.570 142.050 ;
        RECT 61.290 141.880 61.460 142.050 ;
        RECT 61.650 141.880 61.820 142.050 ;
        RECT 62.010 141.880 62.180 142.050 ;
        RECT 63.100 141.880 63.270 142.050 ;
        RECT 63.540 141.880 63.710 142.050 ;
        RECT 63.980 141.880 64.150 142.050 ;
        RECT 64.390 141.880 64.560 142.050 ;
        RECT 65.350 141.880 65.520 142.050 ;
        RECT 65.710 141.880 65.880 142.050 ;
        RECT 66.070 141.880 66.240 142.050 ;
        RECT 66.430 141.880 66.600 142.050 ;
        RECT 67.950 141.890 68.120 142.060 ;
        RECT 68.390 141.890 68.560 142.060 ;
        RECT 68.800 141.890 68.970 142.060 ;
        RECT 69.230 141.890 69.400 142.060 ;
        RECT 69.670 141.890 69.840 142.060 ;
        RECT 70.080 141.890 70.250 142.060 ;
        RECT 71.160 141.880 71.330 142.050 ;
        RECT 71.520 141.880 71.690 142.050 ;
        RECT 72.700 141.880 72.870 142.050 ;
        RECT 73.140 141.880 73.310 142.050 ;
        RECT 73.580 141.880 73.750 142.050 ;
        RECT 73.990 141.880 74.160 142.050 ;
        RECT 74.950 141.880 75.120 142.050 ;
        RECT 75.310 141.880 75.480 142.050 ;
        RECT 75.670 141.880 75.840 142.050 ;
        RECT 76.030 141.880 76.200 142.050 ;
        RECT 77.020 141.880 77.190 142.050 ;
        RECT 77.460 141.880 77.630 142.050 ;
        RECT 77.900 141.880 78.070 142.050 ;
        RECT 78.310 141.880 78.480 142.050 ;
        RECT 79.310 141.880 79.480 142.050 ;
        RECT 79.670 141.880 79.840 142.050 ;
        RECT 80.030 141.880 80.200 142.050 ;
        RECT 80.950 141.880 81.120 142.050 ;
        RECT 81.310 141.880 81.480 142.050 ;
        RECT 85.910 141.880 86.080 142.050 ;
        RECT 86.270 141.880 86.440 142.050 ;
        RECT 86.630 141.880 86.800 142.050 ;
        RECT 89.880 141.880 90.050 142.050 ;
        RECT 90.240 141.880 90.410 142.050 ;
        RECT 90.600 141.880 90.770 142.050 ;
        RECT 92.490 141.880 92.660 142.050 ;
        RECT 92.850 141.880 93.020 142.050 ;
        RECT 93.210 141.880 93.380 142.050 ;
        RECT 94.830 141.890 95.000 142.060 ;
        RECT 95.270 141.890 95.440 142.060 ;
        RECT 95.680 141.890 95.850 142.060 ;
        RECT 96.110 141.890 96.280 142.060 ;
        RECT 96.550 141.890 96.720 142.060 ;
        RECT 96.960 141.890 97.130 142.060 ;
        RECT 98.510 141.880 98.680 142.050 ;
        RECT 98.870 141.880 99.040 142.050 ;
        RECT 99.230 141.880 99.400 142.050 ;
        RECT 100.150 141.880 100.320 142.050 ;
        RECT 100.510 141.880 100.680 142.050 ;
        RECT 105.110 141.880 105.280 142.050 ;
        RECT 105.470 141.880 105.640 142.050 ;
        RECT 105.830 141.880 106.000 142.050 ;
        RECT 109.080 141.880 109.250 142.050 ;
        RECT 109.440 141.880 109.610 142.050 ;
        RECT 109.800 141.880 109.970 142.050 ;
        RECT 111.690 141.880 111.860 142.050 ;
        RECT 112.050 141.880 112.220 142.050 ;
        RECT 112.410 141.880 112.580 142.050 ;
        RECT 114.030 141.890 114.200 142.060 ;
        RECT 114.470 141.890 114.640 142.060 ;
        RECT 114.880 141.890 115.050 142.060 ;
        RECT 115.310 141.890 115.480 142.060 ;
        RECT 115.750 141.890 115.920 142.060 ;
        RECT 116.160 141.890 116.330 142.060 ;
        RECT 117.870 141.890 118.040 142.060 ;
        RECT 118.310 141.890 118.480 142.060 ;
        RECT 118.720 141.890 118.890 142.060 ;
        RECT 119.150 141.890 119.320 142.060 ;
        RECT 119.590 141.890 119.760 142.060 ;
        RECT 120.000 141.890 120.170 142.060 ;
        RECT 121.710 141.890 121.880 142.060 ;
        RECT 122.150 141.890 122.320 142.060 ;
        RECT 122.560 141.890 122.730 142.060 ;
        RECT 122.990 141.890 123.160 142.060 ;
        RECT 123.430 141.890 123.600 142.060 ;
        RECT 123.840 141.890 124.010 142.060 ;
        RECT 125.550 141.890 125.720 142.060 ;
        RECT 125.990 141.890 126.160 142.060 ;
        RECT 126.400 141.890 126.570 142.060 ;
        RECT 126.830 141.890 127.000 142.060 ;
        RECT 127.270 141.890 127.440 142.060 ;
        RECT 127.680 141.890 127.850 142.060 ;
        RECT 129.390 141.890 129.560 142.060 ;
        RECT 129.830 141.890 130.000 142.060 ;
        RECT 130.240 141.890 130.410 142.060 ;
        RECT 130.670 141.890 130.840 142.060 ;
        RECT 131.110 141.890 131.280 142.060 ;
        RECT 131.520 141.890 131.690 142.060 ;
        RECT 133.230 141.890 133.400 142.060 ;
        RECT 133.670 141.890 133.840 142.060 ;
        RECT 134.080 141.890 134.250 142.060 ;
        RECT 134.510 141.890 134.680 142.060 ;
        RECT 134.950 141.890 135.120 142.060 ;
        RECT 135.360 141.890 135.530 142.060 ;
        RECT 137.070 141.890 137.240 142.060 ;
        RECT 137.510 141.890 137.680 142.060 ;
        RECT 137.920 141.890 138.090 142.060 ;
        RECT 138.350 141.890 138.520 142.060 ;
        RECT 138.790 141.890 138.960 142.060 ;
        RECT 139.200 141.890 139.370 142.060 ;
        RECT 140.380 141.880 140.550 142.050 ;
        RECT 140.820 141.880 140.990 142.050 ;
        RECT 141.260 141.880 141.430 142.050 ;
        RECT 141.670 141.880 141.840 142.050 ;
        RECT 5.920 134.220 6.090 134.400 ;
        RECT 6.400 134.220 6.570 134.400 ;
        RECT 6.880 134.220 7.050 134.400 ;
        RECT 7.360 134.220 7.530 134.400 ;
        RECT 7.840 134.220 8.010 134.400 ;
        RECT 8.320 134.220 8.490 134.400 ;
        RECT 8.800 134.220 8.970 134.400 ;
        RECT 9.280 134.220 9.450 134.400 ;
        RECT 9.760 134.220 9.930 134.400 ;
        RECT 10.240 134.220 10.410 134.400 ;
        RECT 10.720 134.220 10.890 134.400 ;
        RECT 11.200 134.220 11.370 134.400 ;
        RECT 11.680 134.220 11.850 134.400 ;
        RECT 12.160 134.220 12.330 134.400 ;
        RECT 12.640 134.220 12.810 134.400 ;
        RECT 13.120 134.220 13.290 134.400 ;
        RECT 13.600 134.220 13.770 134.400 ;
        RECT 14.080 134.220 14.250 134.400 ;
        RECT 14.560 134.220 14.730 134.400 ;
        RECT 15.040 134.220 15.210 134.400 ;
        RECT 15.520 134.220 15.690 134.400 ;
        RECT 16.000 134.220 16.170 134.400 ;
        RECT 16.480 134.220 16.650 134.400 ;
        RECT 16.960 134.220 17.130 134.400 ;
        RECT 17.440 134.220 17.610 134.400 ;
        RECT 17.920 134.220 18.090 134.400 ;
        RECT 18.400 134.220 18.570 134.400 ;
        RECT 18.880 134.220 19.050 134.400 ;
        RECT 19.360 134.220 19.530 134.400 ;
        RECT 19.840 134.220 20.010 134.400 ;
        RECT 20.320 134.220 20.490 134.400 ;
        RECT 20.800 134.220 20.970 134.400 ;
        RECT 21.280 134.220 21.450 134.400 ;
        RECT 21.760 134.220 21.930 134.400 ;
        RECT 22.240 134.220 22.410 134.400 ;
        RECT 22.720 134.220 22.890 134.400 ;
        RECT 23.200 134.220 23.370 134.400 ;
        RECT 23.680 134.220 23.850 134.400 ;
        RECT 24.160 134.220 24.330 134.400 ;
        RECT 24.640 134.220 24.810 134.400 ;
        RECT 25.120 134.220 25.290 134.400 ;
        RECT 25.600 134.220 25.770 134.400 ;
        RECT 26.080 134.220 26.250 134.400 ;
        RECT 26.560 134.220 26.730 134.400 ;
        RECT 27.040 134.220 27.210 134.400 ;
        RECT 27.520 134.220 27.690 134.400 ;
        RECT 28.000 134.220 28.170 134.400 ;
        RECT 28.480 134.220 28.650 134.400 ;
        RECT 28.960 134.220 29.130 134.400 ;
        RECT 29.440 134.220 29.610 134.400 ;
        RECT 29.920 134.220 30.090 134.400 ;
      LAYER li1 ;
        RECT 30.240 134.220 30.720 134.400 ;
      LAYER li1 ;
        RECT 30.880 134.220 31.050 134.400 ;
        RECT 31.360 134.220 31.530 134.400 ;
        RECT 31.840 134.220 32.010 134.400 ;
        RECT 32.320 134.220 32.490 134.400 ;
        RECT 32.800 134.220 32.970 134.400 ;
        RECT 33.280 134.220 33.450 134.400 ;
        RECT 33.760 134.220 33.930 134.400 ;
        RECT 34.240 134.220 34.410 134.400 ;
        RECT 34.720 134.220 34.890 134.400 ;
        RECT 35.200 134.220 35.370 134.400 ;
        RECT 35.680 134.220 35.850 134.400 ;
        RECT 36.160 134.220 36.330 134.400 ;
        RECT 36.640 134.220 36.810 134.400 ;
        RECT 37.120 134.220 37.290 134.400 ;
        RECT 37.600 134.220 37.770 134.400 ;
        RECT 38.080 134.220 38.250 134.400 ;
        RECT 38.560 134.220 38.730 134.400 ;
        RECT 39.040 134.220 39.210 134.400 ;
        RECT 39.520 134.220 39.690 134.400 ;
        RECT 40.000 134.220 40.170 134.400 ;
        RECT 40.480 134.220 40.650 134.400 ;
        RECT 40.960 134.220 41.130 134.400 ;
        RECT 41.440 134.220 41.610 134.400 ;
        RECT 41.920 134.220 42.090 134.400 ;
        RECT 42.400 134.220 42.570 134.400 ;
        RECT 42.880 134.220 43.050 134.400 ;
        RECT 43.360 134.220 43.530 134.400 ;
        RECT 43.840 134.220 44.010 134.400 ;
        RECT 44.320 134.220 44.490 134.400 ;
        RECT 44.800 134.220 44.970 134.400 ;
        RECT 45.280 134.220 45.450 134.400 ;
        RECT 45.760 134.220 45.930 134.400 ;
        RECT 46.240 134.220 46.410 134.400 ;
        RECT 46.720 134.220 46.890 134.400 ;
        RECT 47.200 134.220 47.370 134.400 ;
        RECT 47.680 134.220 47.850 134.400 ;
        RECT 48.160 134.220 48.330 134.400 ;
        RECT 48.640 134.220 48.810 134.400 ;
        RECT 49.120 134.220 49.290 134.400 ;
        RECT 49.600 134.220 49.770 134.400 ;
        RECT 50.080 134.220 50.250 134.400 ;
        RECT 50.560 134.220 50.730 134.400 ;
        RECT 51.040 134.220 51.210 134.400 ;
        RECT 51.520 134.220 51.690 134.400 ;
        RECT 52.000 134.220 52.170 134.400 ;
        RECT 52.480 134.220 52.650 134.400 ;
        RECT 52.960 134.220 53.130 134.400 ;
        RECT 53.440 134.220 53.610 134.400 ;
        RECT 53.920 134.220 54.090 134.400 ;
        RECT 54.400 134.220 54.570 134.400 ;
        RECT 54.880 134.220 55.050 134.400 ;
        RECT 55.360 134.220 55.530 134.400 ;
        RECT 55.840 134.220 56.010 134.400 ;
        RECT 56.320 134.220 56.490 134.400 ;
        RECT 56.800 134.220 56.970 134.400 ;
        RECT 57.280 134.220 57.450 134.400 ;
        RECT 57.760 134.220 57.930 134.400 ;
        RECT 58.240 134.220 58.410 134.400 ;
        RECT 58.720 134.220 58.890 134.400 ;
        RECT 59.200 134.220 59.370 134.400 ;
        RECT 59.680 134.220 59.850 134.400 ;
        RECT 60.160 134.220 60.330 134.400 ;
        RECT 60.640 134.220 60.810 134.400 ;
        RECT 61.120 134.220 61.290 134.400 ;
        RECT 61.600 134.220 61.770 134.400 ;
        RECT 62.080 134.220 62.250 134.400 ;
      LAYER li1 ;
        RECT 62.400 134.220 62.880 134.400 ;
      LAYER li1 ;
        RECT 63.040 134.220 63.210 134.400 ;
        RECT 63.520 134.220 63.690 134.400 ;
        RECT 64.000 134.220 64.170 134.400 ;
        RECT 64.480 134.220 64.650 134.400 ;
        RECT 64.960 134.220 65.130 134.400 ;
        RECT 65.440 134.220 65.610 134.400 ;
        RECT 65.920 134.220 66.090 134.400 ;
        RECT 66.400 134.220 66.570 134.400 ;
        RECT 66.880 134.220 67.050 134.400 ;
        RECT 67.360 134.220 67.530 134.400 ;
        RECT 67.840 134.220 68.010 134.400 ;
        RECT 68.320 134.220 68.490 134.400 ;
        RECT 68.800 134.220 68.970 134.400 ;
        RECT 69.280 134.220 69.450 134.400 ;
        RECT 69.760 134.220 69.930 134.400 ;
        RECT 70.240 134.220 70.410 134.400 ;
        RECT 70.720 134.220 70.890 134.400 ;
        RECT 71.200 134.220 71.370 134.400 ;
        RECT 71.680 134.220 71.850 134.400 ;
        RECT 72.160 134.220 72.330 134.400 ;
        RECT 72.640 134.220 72.810 134.400 ;
        RECT 73.120 134.220 73.290 134.400 ;
        RECT 73.600 134.220 73.770 134.400 ;
        RECT 74.080 134.220 74.250 134.400 ;
        RECT 74.560 134.220 74.730 134.400 ;
      LAYER li1 ;
        RECT 74.880 134.220 75.360 134.400 ;
      LAYER li1 ;
        RECT 75.520 134.220 75.690 134.400 ;
        RECT 76.000 134.220 76.170 134.400 ;
        RECT 76.480 134.220 76.650 134.400 ;
        RECT 76.960 134.220 77.130 134.400 ;
        RECT 77.440 134.220 77.610 134.400 ;
        RECT 77.920 134.220 78.090 134.400 ;
        RECT 78.400 134.220 78.570 134.400 ;
        RECT 78.880 134.220 79.050 134.400 ;
        RECT 79.360 134.220 79.530 134.400 ;
        RECT 79.840 134.220 80.010 134.400 ;
        RECT 80.320 134.220 80.490 134.400 ;
        RECT 80.800 134.220 80.970 134.400 ;
        RECT 81.280 134.220 81.450 134.400 ;
        RECT 81.760 134.220 81.930 134.400 ;
        RECT 82.240 134.220 82.410 134.400 ;
        RECT 82.720 134.220 82.890 134.400 ;
        RECT 83.200 134.220 83.370 134.400 ;
        RECT 83.680 134.220 83.850 134.400 ;
        RECT 84.160 134.220 84.330 134.400 ;
        RECT 84.640 134.220 84.810 134.400 ;
        RECT 85.120 134.220 85.290 134.400 ;
        RECT 85.600 134.220 85.770 134.400 ;
        RECT 86.080 134.220 86.250 134.400 ;
        RECT 86.560 134.220 86.730 134.400 ;
        RECT 87.040 134.220 87.210 134.400 ;
        RECT 87.520 134.220 87.690 134.400 ;
        RECT 88.000 134.220 88.170 134.400 ;
        RECT 88.480 134.220 88.650 134.400 ;
        RECT 88.960 134.220 89.130 134.400 ;
        RECT 89.440 134.220 89.610 134.400 ;
        RECT 89.920 134.220 90.090 134.400 ;
        RECT 90.400 134.220 90.570 134.400 ;
        RECT 90.880 134.220 91.050 134.400 ;
        RECT 91.360 134.220 91.530 134.400 ;
        RECT 91.840 134.220 92.010 134.400 ;
        RECT 92.320 134.220 92.490 134.400 ;
        RECT 92.800 134.220 92.970 134.400 ;
        RECT 93.280 134.220 93.450 134.400 ;
        RECT 93.760 134.220 93.930 134.400 ;
        RECT 94.240 134.220 94.410 134.400 ;
        RECT 94.720 134.220 94.890 134.400 ;
        RECT 95.200 134.220 95.370 134.400 ;
        RECT 95.680 134.220 95.850 134.400 ;
        RECT 96.160 134.220 96.330 134.400 ;
        RECT 96.640 134.220 96.810 134.400 ;
        RECT 97.120 134.220 97.290 134.400 ;
        RECT 97.600 134.220 97.770 134.400 ;
      LAYER li1 ;
        RECT 97.920 134.220 98.400 134.400 ;
      LAYER li1 ;
        RECT 98.560 134.220 98.730 134.400 ;
        RECT 99.040 134.220 99.210 134.400 ;
        RECT 99.520 134.220 99.690 134.400 ;
        RECT 100.000 134.220 100.170 134.400 ;
        RECT 100.480 134.220 100.650 134.400 ;
        RECT 100.960 134.220 101.130 134.400 ;
        RECT 101.440 134.220 101.610 134.400 ;
        RECT 101.920 134.220 102.090 134.400 ;
        RECT 102.400 134.220 102.570 134.400 ;
        RECT 102.880 134.220 103.050 134.400 ;
        RECT 103.360 134.220 103.530 134.400 ;
        RECT 103.840 134.220 104.010 134.400 ;
        RECT 104.320 134.220 104.490 134.400 ;
        RECT 104.800 134.220 104.970 134.400 ;
        RECT 105.280 134.220 105.450 134.400 ;
        RECT 105.760 134.220 105.930 134.400 ;
        RECT 106.240 134.220 106.410 134.400 ;
        RECT 106.720 134.220 106.890 134.400 ;
        RECT 107.200 134.220 107.370 134.400 ;
        RECT 107.680 134.220 107.850 134.400 ;
        RECT 108.160 134.220 108.330 134.400 ;
        RECT 108.640 134.220 108.810 134.400 ;
        RECT 109.120 134.220 109.290 134.400 ;
      LAYER li1 ;
        RECT 109.440 134.220 109.920 134.400 ;
      LAYER li1 ;
        RECT 110.080 134.220 110.250 134.400 ;
        RECT 110.560 134.220 110.730 134.400 ;
        RECT 111.040 134.220 111.210 134.400 ;
        RECT 111.520 134.220 111.690 134.400 ;
        RECT 112.000 134.220 112.170 134.400 ;
        RECT 112.480 134.220 112.650 134.400 ;
        RECT 112.960 134.220 113.130 134.400 ;
        RECT 113.440 134.220 113.610 134.400 ;
        RECT 113.920 134.220 114.090 134.400 ;
        RECT 114.400 134.220 114.570 134.400 ;
        RECT 114.880 134.220 115.050 134.400 ;
        RECT 115.360 134.220 115.530 134.400 ;
        RECT 115.840 134.220 116.010 134.400 ;
        RECT 116.320 134.220 116.490 134.400 ;
        RECT 116.800 134.220 116.970 134.400 ;
        RECT 117.280 134.220 117.450 134.400 ;
        RECT 117.760 134.220 117.930 134.400 ;
        RECT 118.240 134.220 118.410 134.400 ;
        RECT 118.720 134.220 118.890 134.400 ;
        RECT 119.200 134.220 119.370 134.400 ;
        RECT 119.680 134.220 119.850 134.400 ;
        RECT 120.160 134.220 120.330 134.400 ;
        RECT 120.640 134.220 120.810 134.400 ;
        RECT 121.120 134.220 121.290 134.400 ;
        RECT 121.600 134.220 121.770 134.400 ;
        RECT 122.080 134.220 122.250 134.400 ;
        RECT 122.560 134.220 122.730 134.400 ;
        RECT 123.040 134.220 123.210 134.400 ;
        RECT 123.520 134.220 123.690 134.400 ;
        RECT 124.000 134.220 124.170 134.400 ;
        RECT 124.480 134.220 124.650 134.400 ;
        RECT 124.960 134.220 125.130 134.400 ;
        RECT 125.440 134.220 125.610 134.400 ;
        RECT 125.920 134.220 126.090 134.400 ;
        RECT 126.400 134.220 126.570 134.400 ;
        RECT 126.880 134.220 127.050 134.400 ;
        RECT 127.360 134.220 127.530 134.400 ;
        RECT 127.840 134.220 128.010 134.400 ;
        RECT 128.320 134.220 128.490 134.400 ;
        RECT 128.800 134.220 128.970 134.400 ;
        RECT 129.280 134.220 129.450 134.400 ;
        RECT 129.760 134.220 129.930 134.400 ;
        RECT 130.240 134.220 130.410 134.400 ;
        RECT 130.720 134.220 130.890 134.400 ;
        RECT 131.200 134.220 131.370 134.400 ;
        RECT 131.680 134.220 131.850 134.400 ;
        RECT 132.160 134.220 132.330 134.400 ;
        RECT 132.640 134.220 132.810 134.400 ;
        RECT 133.120 134.220 133.290 134.400 ;
        RECT 133.600 134.220 133.770 134.400 ;
        RECT 134.080 134.220 134.250 134.400 ;
        RECT 134.560 134.220 134.730 134.400 ;
        RECT 135.040 134.220 135.210 134.400 ;
        RECT 135.520 134.220 135.690 134.400 ;
        RECT 136.000 134.220 136.170 134.400 ;
        RECT 136.480 134.220 136.650 134.400 ;
        RECT 136.960 134.220 137.130 134.400 ;
        RECT 137.440 134.220 137.610 134.400 ;
        RECT 137.920 134.220 138.090 134.400 ;
        RECT 138.400 134.220 138.570 134.400 ;
        RECT 138.880 134.220 139.050 134.400 ;
        RECT 139.360 134.220 139.530 134.400 ;
        RECT 139.840 134.220 140.010 134.400 ;
        RECT 140.320 134.220 140.490 134.400 ;
        RECT 140.800 134.220 140.970 134.400 ;
        RECT 141.280 134.220 141.450 134.400 ;
      LAYER li1 ;
        RECT 141.600 134.220 142.080 134.400 ;
      LAYER li1 ;
        RECT 6.510 133.750 6.680 133.920 ;
        RECT 6.950 133.750 7.120 133.920 ;
        RECT 7.360 133.750 7.530 133.920 ;
        RECT 7.790 133.750 7.960 133.920 ;
        RECT 8.230 133.750 8.400 133.920 ;
        RECT 8.640 133.750 8.810 133.920 ;
        RECT 12.160 133.740 12.330 133.910 ;
        RECT 12.520 133.740 12.690 133.910 ;
        RECT 13.710 133.750 13.880 133.920 ;
        RECT 14.150 133.750 14.320 133.920 ;
        RECT 14.560 133.750 14.730 133.920 ;
        RECT 14.990 133.750 15.160 133.920 ;
        RECT 15.430 133.750 15.600 133.920 ;
        RECT 15.840 133.750 16.010 133.920 ;
        RECT 17.550 133.750 17.720 133.920 ;
        RECT 17.990 133.750 18.160 133.920 ;
        RECT 18.400 133.750 18.570 133.920 ;
        RECT 18.830 133.750 19.000 133.920 ;
        RECT 19.270 133.750 19.440 133.920 ;
        RECT 19.680 133.750 19.850 133.920 ;
        RECT 21.390 133.750 21.560 133.920 ;
        RECT 21.830 133.750 22.000 133.920 ;
        RECT 22.240 133.750 22.410 133.920 ;
        RECT 22.670 133.750 22.840 133.920 ;
        RECT 23.110 133.750 23.280 133.920 ;
        RECT 23.520 133.750 23.690 133.920 ;
        RECT 25.230 133.750 25.400 133.920 ;
        RECT 25.670 133.750 25.840 133.920 ;
        RECT 26.080 133.750 26.250 133.920 ;
        RECT 26.510 133.750 26.680 133.920 ;
        RECT 26.950 133.750 27.120 133.920 ;
        RECT 27.360 133.750 27.530 133.920 ;
        RECT 28.540 133.740 28.710 133.910 ;
        RECT 28.980 133.740 29.150 133.910 ;
        RECT 29.420 133.740 29.590 133.910 ;
        RECT 29.830 133.740 30.000 133.910 ;
        RECT 33.880 133.740 34.050 133.910 ;
        RECT 34.240 133.740 34.410 133.910 ;
        RECT 34.600 133.740 34.770 133.910 ;
        RECT 36.270 133.750 36.440 133.920 ;
        RECT 36.710 133.750 36.880 133.920 ;
        RECT 37.120 133.750 37.290 133.920 ;
        RECT 37.550 133.750 37.720 133.920 ;
        RECT 37.990 133.750 38.160 133.920 ;
        RECT 38.400 133.750 38.570 133.920 ;
        RECT 40.110 133.750 40.280 133.920 ;
        RECT 40.550 133.750 40.720 133.920 ;
        RECT 40.960 133.750 41.130 133.920 ;
        RECT 41.390 133.750 41.560 133.920 ;
        RECT 41.830 133.750 42.000 133.920 ;
        RECT 42.240 133.750 42.410 133.920 ;
        RECT 43.950 133.750 44.120 133.920 ;
        RECT 44.390 133.750 44.560 133.920 ;
        RECT 44.800 133.750 44.970 133.920 ;
        RECT 45.230 133.750 45.400 133.920 ;
        RECT 45.670 133.750 45.840 133.920 ;
        RECT 46.080 133.750 46.250 133.920 ;
        RECT 47.790 133.750 47.960 133.920 ;
        RECT 48.230 133.750 48.400 133.920 ;
        RECT 48.640 133.750 48.810 133.920 ;
        RECT 49.070 133.750 49.240 133.920 ;
        RECT 49.510 133.750 49.680 133.920 ;
        RECT 49.920 133.750 50.090 133.920 ;
        RECT 51.630 133.750 51.800 133.920 ;
        RECT 52.070 133.750 52.240 133.920 ;
        RECT 52.480 133.750 52.650 133.920 ;
        RECT 52.910 133.750 53.080 133.920 ;
        RECT 53.350 133.750 53.520 133.920 ;
        RECT 53.760 133.750 53.930 133.920 ;
        RECT 55.470 133.750 55.640 133.920 ;
        RECT 55.910 133.750 56.080 133.920 ;
        RECT 56.320 133.750 56.490 133.920 ;
        RECT 56.750 133.750 56.920 133.920 ;
        RECT 57.190 133.750 57.360 133.920 ;
        RECT 57.600 133.750 57.770 133.920 ;
        RECT 59.310 133.750 59.480 133.920 ;
        RECT 59.750 133.750 59.920 133.920 ;
        RECT 60.160 133.750 60.330 133.920 ;
        RECT 60.590 133.750 60.760 133.920 ;
        RECT 61.030 133.750 61.200 133.920 ;
        RECT 61.440 133.750 61.610 133.920 ;
        RECT 63.150 133.750 63.320 133.920 ;
        RECT 63.590 133.750 63.760 133.920 ;
        RECT 64.000 133.750 64.170 133.920 ;
        RECT 64.430 133.750 64.600 133.920 ;
        RECT 64.870 133.750 65.040 133.920 ;
        RECT 65.280 133.750 65.450 133.920 ;
        RECT 66.990 133.750 67.160 133.920 ;
        RECT 67.430 133.750 67.600 133.920 ;
        RECT 67.840 133.750 68.010 133.920 ;
        RECT 68.270 133.750 68.440 133.920 ;
        RECT 68.710 133.750 68.880 133.920 ;
        RECT 69.120 133.750 69.290 133.920 ;
        RECT 70.300 133.740 70.470 133.910 ;
        RECT 70.740 133.740 70.910 133.910 ;
        RECT 71.180 133.740 71.350 133.910 ;
        RECT 71.590 133.740 71.760 133.910 ;
        RECT 75.130 133.740 75.300 133.910 ;
        RECT 75.490 133.740 75.660 133.910 ;
        RECT 75.850 133.740 76.020 133.910 ;
        RECT 77.020 133.740 77.190 133.910 ;
        RECT 77.460 133.740 77.630 133.910 ;
        RECT 77.900 133.740 78.070 133.910 ;
        RECT 78.310 133.740 78.480 133.910 ;
        RECT 78.840 133.740 79.010 133.910 ;
        RECT 79.200 133.740 79.370 133.910 ;
        RECT 80.110 133.740 80.280 133.910 ;
        RECT 80.470 133.740 80.640 133.910 ;
        RECT 80.830 133.740 81.000 133.910 ;
        RECT 82.300 133.740 82.470 133.910 ;
        RECT 82.740 133.740 82.910 133.910 ;
        RECT 83.180 133.740 83.350 133.910 ;
        RECT 83.590 133.740 83.760 133.910 ;
        RECT 85.520 133.740 85.690 133.910 ;
        RECT 85.880 133.740 86.050 133.910 ;
        RECT 86.240 133.740 86.410 133.910 ;
        RECT 88.880 133.740 89.050 133.910 ;
        RECT 89.240 133.740 89.410 133.910 ;
        RECT 89.600 133.740 89.770 133.910 ;
        RECT 89.960 133.740 90.130 133.910 ;
        RECT 90.990 133.750 91.160 133.920 ;
        RECT 91.430 133.750 91.600 133.920 ;
        RECT 91.840 133.750 92.010 133.920 ;
        RECT 92.270 133.750 92.440 133.920 ;
        RECT 92.710 133.750 92.880 133.920 ;
        RECT 93.120 133.750 93.290 133.920 ;
        RECT 94.830 133.750 95.000 133.920 ;
        RECT 95.270 133.750 95.440 133.920 ;
        RECT 95.680 133.750 95.850 133.920 ;
        RECT 96.110 133.750 96.280 133.920 ;
        RECT 96.550 133.750 96.720 133.920 ;
        RECT 96.960 133.750 97.130 133.920 ;
        RECT 98.480 133.740 98.650 133.910 ;
        RECT 98.840 133.740 99.010 133.910 ;
        RECT 99.200 133.740 99.370 133.910 ;
        RECT 101.840 133.740 102.010 133.910 ;
        RECT 102.200 133.740 102.370 133.910 ;
        RECT 102.560 133.740 102.730 133.910 ;
        RECT 102.920 133.740 103.090 133.910 ;
        RECT 103.420 133.740 103.590 133.910 ;
        RECT 103.860 133.740 104.030 133.910 ;
        RECT 104.300 133.740 104.470 133.910 ;
        RECT 104.710 133.740 104.880 133.910 ;
        RECT 105.760 133.740 105.930 133.910 ;
        RECT 106.120 133.740 106.290 133.910 ;
        RECT 106.480 133.740 106.650 133.910 ;
        RECT 108.700 133.740 108.870 133.910 ;
        RECT 109.140 133.740 109.310 133.910 ;
        RECT 109.580 133.740 109.750 133.910 ;
        RECT 109.990 133.740 110.160 133.910 ;
        RECT 111.470 133.740 111.640 133.910 ;
        RECT 111.830 133.740 112.000 133.910 ;
        RECT 112.190 133.740 112.360 133.910 ;
        RECT 113.110 133.740 113.280 133.910 ;
        RECT 113.470 133.740 113.640 133.910 ;
        RECT 118.070 133.740 118.240 133.910 ;
        RECT 118.430 133.740 118.600 133.910 ;
        RECT 118.790 133.740 118.960 133.910 ;
        RECT 122.040 133.740 122.210 133.910 ;
        RECT 122.400 133.740 122.570 133.910 ;
        RECT 122.760 133.740 122.930 133.910 ;
        RECT 124.650 133.740 124.820 133.910 ;
        RECT 125.010 133.740 125.180 133.910 ;
        RECT 125.370 133.740 125.540 133.910 ;
        RECT 126.990 133.750 127.160 133.920 ;
        RECT 127.430 133.750 127.600 133.920 ;
        RECT 127.840 133.750 128.010 133.920 ;
        RECT 128.270 133.750 128.440 133.920 ;
        RECT 128.710 133.750 128.880 133.920 ;
        RECT 129.120 133.750 129.290 133.920 ;
        RECT 130.830 133.750 131.000 133.920 ;
        RECT 131.270 133.750 131.440 133.920 ;
        RECT 131.680 133.750 131.850 133.920 ;
        RECT 132.110 133.750 132.280 133.920 ;
        RECT 132.550 133.750 132.720 133.920 ;
        RECT 132.960 133.750 133.130 133.920 ;
        RECT 134.670 133.750 134.840 133.920 ;
        RECT 135.110 133.750 135.280 133.920 ;
        RECT 135.520 133.750 135.690 133.920 ;
        RECT 135.950 133.750 136.120 133.920 ;
        RECT 136.390 133.750 136.560 133.920 ;
        RECT 136.800 133.750 136.970 133.920 ;
        RECT 138.510 133.750 138.680 133.920 ;
        RECT 138.950 133.750 139.120 133.920 ;
        RECT 139.360 133.750 139.530 133.920 ;
        RECT 139.790 133.750 139.960 133.920 ;
        RECT 140.230 133.750 140.400 133.920 ;
        RECT 140.640 133.750 140.810 133.920 ;
        RECT 5.920 126.080 6.090 126.260 ;
        RECT 6.400 126.080 6.570 126.260 ;
        RECT 6.880 126.080 7.050 126.260 ;
        RECT 7.360 126.080 7.530 126.260 ;
        RECT 7.840 126.080 8.010 126.260 ;
        RECT 8.320 126.080 8.490 126.260 ;
        RECT 8.800 126.080 8.970 126.260 ;
        RECT 9.280 126.080 9.450 126.260 ;
        RECT 9.760 126.080 9.930 126.260 ;
        RECT 10.240 126.080 10.410 126.260 ;
        RECT 10.720 126.080 10.890 126.260 ;
        RECT 11.200 126.080 11.370 126.260 ;
        RECT 11.680 126.080 11.850 126.260 ;
        RECT 12.160 126.080 12.330 126.260 ;
        RECT 12.640 126.080 12.810 126.260 ;
        RECT 13.120 126.080 13.290 126.260 ;
        RECT 13.600 126.080 13.770 126.260 ;
        RECT 14.080 126.080 14.250 126.260 ;
        RECT 14.560 126.080 14.730 126.260 ;
        RECT 15.040 126.080 15.210 126.260 ;
        RECT 15.520 126.080 15.690 126.260 ;
        RECT 16.000 126.080 16.170 126.260 ;
        RECT 16.480 126.080 16.650 126.260 ;
        RECT 16.960 126.080 17.130 126.260 ;
        RECT 17.440 126.080 17.610 126.260 ;
        RECT 17.920 126.080 18.090 126.260 ;
        RECT 18.400 126.080 18.570 126.260 ;
        RECT 18.880 126.080 19.050 126.260 ;
        RECT 19.360 126.080 19.530 126.260 ;
        RECT 19.840 126.080 20.010 126.260 ;
        RECT 20.320 126.080 20.490 126.260 ;
        RECT 20.800 126.080 20.970 126.260 ;
        RECT 21.280 126.080 21.450 126.260 ;
        RECT 21.760 126.080 21.930 126.260 ;
        RECT 22.240 126.080 22.410 126.260 ;
        RECT 22.720 126.080 22.890 126.260 ;
        RECT 23.200 126.080 23.370 126.260 ;
        RECT 23.680 126.080 23.850 126.260 ;
        RECT 24.160 126.080 24.330 126.260 ;
        RECT 24.640 126.080 24.810 126.260 ;
        RECT 25.120 126.080 25.290 126.260 ;
        RECT 25.600 126.080 25.770 126.260 ;
        RECT 26.080 126.080 26.250 126.260 ;
        RECT 26.560 126.080 26.730 126.260 ;
        RECT 27.040 126.080 27.210 126.260 ;
        RECT 27.520 126.080 27.690 126.260 ;
        RECT 28.000 126.080 28.170 126.260 ;
        RECT 28.480 126.080 28.650 126.260 ;
        RECT 28.960 126.080 29.130 126.260 ;
        RECT 29.440 126.080 29.610 126.260 ;
        RECT 29.920 126.080 30.090 126.260 ;
        RECT 30.400 126.080 30.570 126.260 ;
        RECT 30.880 126.080 31.050 126.260 ;
        RECT 31.360 126.080 31.530 126.260 ;
        RECT 31.840 126.080 32.010 126.260 ;
        RECT 32.320 126.080 32.490 126.260 ;
        RECT 32.800 126.080 32.970 126.260 ;
        RECT 33.280 126.080 33.450 126.260 ;
        RECT 33.760 126.080 33.930 126.260 ;
      LAYER li1 ;
        RECT 34.080 126.080 34.560 126.260 ;
      LAYER li1 ;
        RECT 34.720 126.080 34.890 126.260 ;
        RECT 35.200 126.080 35.370 126.260 ;
        RECT 35.680 126.080 35.850 126.260 ;
        RECT 36.160 126.080 36.330 126.260 ;
        RECT 36.640 126.080 36.810 126.260 ;
        RECT 37.120 126.080 37.290 126.260 ;
        RECT 37.600 126.080 37.770 126.260 ;
        RECT 38.080 126.080 38.250 126.260 ;
        RECT 38.560 126.080 38.730 126.260 ;
        RECT 39.040 126.080 39.210 126.260 ;
        RECT 39.520 126.080 39.690 126.260 ;
        RECT 40.000 126.080 40.170 126.260 ;
        RECT 40.480 126.080 40.650 126.260 ;
        RECT 40.960 126.080 41.130 126.260 ;
        RECT 41.440 126.080 41.610 126.260 ;
        RECT 41.920 126.080 42.090 126.260 ;
        RECT 42.400 126.080 42.570 126.260 ;
        RECT 42.880 126.080 43.050 126.260 ;
        RECT 43.360 126.080 43.530 126.260 ;
      LAYER li1 ;
        RECT 43.680 126.080 44.160 126.260 ;
      LAYER li1 ;
        RECT 44.320 126.080 44.490 126.260 ;
        RECT 44.800 126.080 44.970 126.260 ;
        RECT 45.280 126.080 45.450 126.260 ;
        RECT 45.760 126.080 45.930 126.260 ;
        RECT 46.240 126.080 46.410 126.260 ;
        RECT 46.720 126.080 46.890 126.260 ;
        RECT 47.200 126.080 47.370 126.260 ;
        RECT 47.680 126.080 47.850 126.260 ;
        RECT 48.160 126.080 48.330 126.260 ;
        RECT 48.640 126.080 48.810 126.260 ;
        RECT 49.120 126.080 49.290 126.260 ;
        RECT 49.600 126.080 49.770 126.260 ;
        RECT 50.080 126.080 50.250 126.260 ;
        RECT 50.560 126.080 50.730 126.260 ;
        RECT 51.040 126.080 51.210 126.260 ;
        RECT 51.520 126.080 51.690 126.260 ;
        RECT 52.000 126.080 52.170 126.260 ;
        RECT 52.480 126.080 52.650 126.260 ;
        RECT 52.960 126.080 53.130 126.260 ;
        RECT 53.440 126.080 53.610 126.260 ;
        RECT 53.920 126.080 54.090 126.260 ;
        RECT 54.400 126.080 54.570 126.260 ;
        RECT 54.880 126.080 55.050 126.260 ;
        RECT 55.360 126.080 55.530 126.260 ;
        RECT 55.840 126.080 56.010 126.260 ;
        RECT 56.320 126.080 56.490 126.260 ;
        RECT 56.800 126.080 56.970 126.260 ;
        RECT 57.280 126.080 57.450 126.260 ;
        RECT 57.760 126.080 57.930 126.260 ;
        RECT 58.240 126.080 58.410 126.260 ;
        RECT 58.720 126.080 58.890 126.260 ;
        RECT 59.200 126.080 59.370 126.260 ;
        RECT 59.680 126.080 59.850 126.260 ;
        RECT 60.160 126.080 60.330 126.260 ;
        RECT 60.640 126.080 60.810 126.260 ;
        RECT 61.120 126.080 61.290 126.260 ;
        RECT 61.600 126.080 61.770 126.260 ;
        RECT 62.080 126.080 62.250 126.260 ;
        RECT 62.560 126.080 62.730 126.260 ;
        RECT 63.040 126.080 63.210 126.260 ;
        RECT 63.520 126.080 63.690 126.260 ;
        RECT 64.000 126.080 64.170 126.260 ;
        RECT 64.480 126.080 64.650 126.260 ;
        RECT 64.960 126.080 65.130 126.260 ;
        RECT 65.440 126.080 65.610 126.260 ;
        RECT 65.920 126.080 66.090 126.260 ;
        RECT 66.400 126.080 66.570 126.260 ;
        RECT 66.880 126.080 67.050 126.260 ;
        RECT 67.360 126.080 67.530 126.260 ;
        RECT 67.840 126.080 68.010 126.260 ;
        RECT 68.320 126.080 68.490 126.260 ;
        RECT 68.800 126.080 68.970 126.260 ;
        RECT 69.280 126.080 69.450 126.260 ;
        RECT 69.760 126.080 69.930 126.260 ;
        RECT 70.240 126.080 70.410 126.260 ;
        RECT 70.720 126.080 70.890 126.260 ;
        RECT 71.200 126.080 71.370 126.260 ;
        RECT 71.680 126.080 71.850 126.260 ;
        RECT 72.160 126.080 72.330 126.260 ;
        RECT 72.640 126.080 72.810 126.260 ;
        RECT 73.120 126.080 73.290 126.260 ;
        RECT 73.600 126.080 73.770 126.260 ;
      LAYER li1 ;
        RECT 73.920 126.080 74.400 126.260 ;
      LAYER li1 ;
        RECT 74.560 126.080 74.730 126.260 ;
        RECT 75.040 126.080 75.210 126.260 ;
        RECT 75.520 126.080 75.690 126.260 ;
        RECT 76.000 126.080 76.170 126.260 ;
        RECT 76.480 126.080 76.650 126.260 ;
        RECT 76.960 126.080 77.130 126.260 ;
        RECT 77.440 126.080 77.610 126.260 ;
        RECT 77.920 126.080 78.090 126.260 ;
        RECT 78.400 126.080 78.570 126.260 ;
        RECT 78.880 126.080 79.050 126.260 ;
        RECT 79.360 126.080 79.530 126.260 ;
        RECT 79.840 126.080 80.010 126.260 ;
        RECT 80.320 126.080 80.490 126.260 ;
        RECT 80.800 126.080 80.970 126.260 ;
        RECT 81.280 126.080 81.450 126.260 ;
        RECT 81.760 126.080 81.930 126.260 ;
        RECT 82.240 126.080 82.410 126.260 ;
        RECT 82.720 126.080 82.890 126.260 ;
        RECT 83.200 126.080 83.370 126.260 ;
        RECT 83.680 126.080 83.850 126.260 ;
        RECT 84.160 126.080 84.330 126.260 ;
        RECT 84.640 126.080 84.810 126.260 ;
        RECT 85.120 126.080 85.290 126.260 ;
        RECT 85.600 126.080 85.770 126.260 ;
        RECT 86.080 126.080 86.250 126.260 ;
        RECT 86.560 126.080 86.730 126.260 ;
        RECT 87.040 126.080 87.210 126.260 ;
        RECT 87.520 126.080 87.690 126.260 ;
        RECT 88.000 126.080 88.170 126.260 ;
        RECT 88.480 126.080 88.650 126.260 ;
        RECT 88.960 126.080 89.130 126.260 ;
        RECT 89.440 126.080 89.610 126.260 ;
        RECT 89.920 126.080 90.090 126.260 ;
        RECT 90.400 126.080 90.570 126.260 ;
        RECT 90.880 126.080 91.050 126.260 ;
        RECT 91.360 126.080 91.530 126.260 ;
        RECT 91.840 126.080 92.010 126.260 ;
        RECT 92.320 126.080 92.490 126.260 ;
        RECT 92.800 126.080 92.970 126.260 ;
        RECT 93.280 126.080 93.450 126.260 ;
        RECT 93.760 126.080 93.930 126.260 ;
        RECT 94.240 126.080 94.410 126.260 ;
        RECT 94.720 126.080 94.890 126.260 ;
        RECT 95.200 126.080 95.370 126.260 ;
        RECT 95.680 126.080 95.850 126.260 ;
        RECT 96.160 126.080 96.330 126.260 ;
        RECT 96.640 126.080 96.810 126.260 ;
        RECT 97.120 126.080 97.290 126.260 ;
        RECT 97.600 126.080 97.770 126.260 ;
        RECT 98.080 126.080 98.250 126.260 ;
        RECT 98.560 126.080 98.730 126.260 ;
        RECT 99.040 126.080 99.210 126.260 ;
        RECT 99.520 126.080 99.690 126.260 ;
        RECT 100.000 126.080 100.170 126.260 ;
        RECT 100.480 126.080 100.650 126.260 ;
        RECT 100.960 126.080 101.130 126.260 ;
        RECT 101.440 126.080 101.610 126.260 ;
        RECT 101.920 126.080 102.090 126.260 ;
        RECT 102.400 126.080 102.570 126.260 ;
        RECT 102.880 126.080 103.050 126.260 ;
        RECT 103.360 126.080 103.530 126.260 ;
        RECT 103.840 126.080 104.010 126.260 ;
        RECT 104.320 126.080 104.490 126.260 ;
        RECT 104.800 126.080 104.970 126.260 ;
        RECT 105.280 126.080 105.450 126.260 ;
        RECT 105.760 126.080 105.930 126.260 ;
        RECT 106.240 126.080 106.410 126.260 ;
        RECT 106.720 126.080 106.890 126.260 ;
        RECT 107.200 126.080 107.370 126.260 ;
        RECT 107.680 126.080 107.850 126.260 ;
        RECT 108.160 126.080 108.330 126.260 ;
        RECT 108.640 126.080 108.810 126.260 ;
        RECT 109.120 126.080 109.290 126.260 ;
        RECT 109.600 126.080 109.770 126.260 ;
        RECT 110.080 126.080 110.250 126.260 ;
      LAYER li1 ;
        RECT 110.400 126.080 110.880 126.260 ;
      LAYER li1 ;
        RECT 111.040 126.080 111.210 126.260 ;
        RECT 111.520 126.080 111.690 126.260 ;
        RECT 112.000 126.080 112.170 126.260 ;
        RECT 112.480 126.080 112.650 126.260 ;
        RECT 112.960 126.080 113.130 126.260 ;
        RECT 113.440 126.080 113.610 126.260 ;
        RECT 113.920 126.080 114.090 126.260 ;
        RECT 114.400 126.080 114.570 126.260 ;
        RECT 114.880 126.080 115.050 126.260 ;
        RECT 115.360 126.080 115.530 126.260 ;
        RECT 115.840 126.080 116.010 126.260 ;
        RECT 116.320 126.080 116.490 126.260 ;
        RECT 116.800 126.080 116.970 126.260 ;
        RECT 117.280 126.080 117.450 126.260 ;
        RECT 117.760 126.080 117.930 126.260 ;
      LAYER li1 ;
        RECT 118.080 126.080 118.560 126.260 ;
      LAYER li1 ;
        RECT 118.720 126.080 118.890 126.260 ;
        RECT 119.200 126.080 119.370 126.260 ;
        RECT 119.680 126.080 119.850 126.260 ;
        RECT 120.160 126.080 120.330 126.260 ;
        RECT 120.640 126.080 120.810 126.260 ;
        RECT 121.120 126.080 121.290 126.260 ;
        RECT 121.600 126.080 121.770 126.260 ;
        RECT 122.080 126.080 122.250 126.260 ;
        RECT 122.560 126.080 122.730 126.260 ;
        RECT 123.040 126.080 123.210 126.260 ;
        RECT 123.520 126.080 123.690 126.260 ;
        RECT 124.000 126.080 124.170 126.260 ;
        RECT 124.480 126.080 124.650 126.260 ;
        RECT 124.960 126.080 125.130 126.260 ;
        RECT 125.440 126.080 125.610 126.260 ;
        RECT 125.920 126.080 126.090 126.260 ;
        RECT 126.400 126.080 126.570 126.260 ;
        RECT 126.880 126.080 127.050 126.260 ;
        RECT 127.360 126.080 127.530 126.260 ;
        RECT 127.840 126.080 128.010 126.260 ;
        RECT 128.320 126.080 128.490 126.260 ;
        RECT 128.800 126.080 128.970 126.260 ;
        RECT 129.280 126.080 129.450 126.260 ;
        RECT 129.760 126.080 129.930 126.260 ;
        RECT 130.240 126.080 130.410 126.260 ;
        RECT 130.720 126.080 130.890 126.260 ;
        RECT 131.200 126.080 131.370 126.260 ;
        RECT 131.680 126.080 131.850 126.260 ;
        RECT 132.160 126.080 132.330 126.260 ;
        RECT 132.640 126.080 132.810 126.260 ;
        RECT 133.120 126.080 133.290 126.260 ;
        RECT 133.600 126.080 133.770 126.260 ;
        RECT 134.080 126.080 134.250 126.260 ;
        RECT 134.560 126.080 134.730 126.260 ;
        RECT 135.040 126.080 135.210 126.260 ;
        RECT 135.520 126.080 135.690 126.260 ;
        RECT 136.000 126.080 136.170 126.260 ;
        RECT 136.480 126.080 136.650 126.260 ;
        RECT 136.960 126.080 137.130 126.260 ;
        RECT 137.440 126.080 137.610 126.260 ;
        RECT 137.920 126.080 138.090 126.260 ;
        RECT 138.400 126.080 138.570 126.260 ;
        RECT 138.880 126.080 139.050 126.260 ;
        RECT 139.360 126.080 139.530 126.260 ;
        RECT 139.840 126.080 140.010 126.260 ;
        RECT 140.320 126.080 140.490 126.260 ;
        RECT 140.800 126.080 140.970 126.260 ;
        RECT 141.280 126.080 141.450 126.260 ;
        RECT 141.760 126.080 141.930 126.260 ;
        RECT 5.980 125.600 6.150 125.770 ;
        RECT 6.420 125.600 6.590 125.770 ;
        RECT 6.860 125.600 7.030 125.770 ;
        RECT 7.270 125.600 7.440 125.770 ;
        RECT 8.750 125.600 8.920 125.770 ;
        RECT 9.110 125.600 9.280 125.770 ;
        RECT 9.470 125.600 9.640 125.770 ;
        RECT 10.390 125.600 10.560 125.770 ;
        RECT 10.750 125.600 10.920 125.770 ;
        RECT 15.350 125.600 15.520 125.770 ;
        RECT 15.710 125.600 15.880 125.770 ;
        RECT 16.070 125.600 16.240 125.770 ;
        RECT 19.320 125.600 19.490 125.770 ;
        RECT 19.680 125.600 19.850 125.770 ;
        RECT 20.040 125.600 20.210 125.770 ;
        RECT 21.930 125.600 22.100 125.770 ;
        RECT 22.290 125.600 22.460 125.770 ;
        RECT 22.650 125.600 22.820 125.770 ;
        RECT 23.740 125.600 23.910 125.770 ;
        RECT 24.180 125.600 24.350 125.770 ;
        RECT 24.620 125.600 24.790 125.770 ;
        RECT 25.030 125.600 25.200 125.770 ;
        RECT 26.990 125.600 27.160 125.770 ;
        RECT 27.350 125.600 27.520 125.770 ;
        RECT 27.710 125.600 27.880 125.770 ;
        RECT 28.630 125.600 28.800 125.770 ;
        RECT 28.990 125.600 29.160 125.770 ;
        RECT 33.590 125.600 33.760 125.770 ;
        RECT 33.950 125.600 34.120 125.770 ;
        RECT 34.310 125.600 34.480 125.770 ;
        RECT 37.560 125.600 37.730 125.770 ;
        RECT 37.920 125.600 38.090 125.770 ;
        RECT 38.280 125.600 38.450 125.770 ;
        RECT 40.170 125.600 40.340 125.770 ;
        RECT 40.530 125.600 40.700 125.770 ;
        RECT 40.890 125.600 41.060 125.770 ;
        RECT 41.980 125.600 42.150 125.770 ;
        RECT 42.420 125.600 42.590 125.770 ;
        RECT 42.860 125.600 43.030 125.770 ;
        RECT 43.270 125.600 43.440 125.770 ;
        RECT 44.760 125.600 44.930 125.770 ;
        RECT 45.120 125.600 45.290 125.770 ;
        RECT 45.480 125.600 45.650 125.770 ;
        RECT 45.840 125.600 46.010 125.770 ;
        RECT 46.200 125.600 46.370 125.770 ;
        RECT 48.010 125.600 48.180 125.770 ;
        RECT 48.370 125.600 48.540 125.770 ;
        RECT 48.730 125.600 48.900 125.770 ;
        RECT 49.090 125.600 49.260 125.770 ;
        RECT 50.190 125.610 50.360 125.780 ;
        RECT 50.630 125.610 50.800 125.780 ;
        RECT 51.040 125.610 51.210 125.780 ;
        RECT 51.470 125.610 51.640 125.780 ;
        RECT 51.910 125.610 52.080 125.780 ;
        RECT 52.320 125.610 52.490 125.780 ;
        RECT 54.030 125.610 54.200 125.780 ;
        RECT 54.470 125.610 54.640 125.780 ;
        RECT 54.880 125.610 55.050 125.780 ;
        RECT 55.310 125.610 55.480 125.780 ;
        RECT 55.750 125.610 55.920 125.780 ;
        RECT 56.160 125.610 56.330 125.780 ;
        RECT 58.630 125.600 58.800 125.770 ;
        RECT 58.990 125.600 59.160 125.770 ;
        RECT 59.350 125.600 59.520 125.770 ;
        RECT 59.710 125.600 59.880 125.770 ;
        RECT 61.230 125.610 61.400 125.780 ;
        RECT 61.670 125.610 61.840 125.780 ;
        RECT 62.080 125.610 62.250 125.780 ;
        RECT 62.510 125.610 62.680 125.780 ;
        RECT 62.950 125.610 63.120 125.780 ;
        RECT 63.360 125.610 63.530 125.780 ;
        RECT 65.070 125.610 65.240 125.780 ;
        RECT 65.510 125.610 65.680 125.780 ;
        RECT 65.920 125.610 66.090 125.780 ;
        RECT 66.350 125.610 66.520 125.780 ;
        RECT 66.790 125.610 66.960 125.780 ;
        RECT 67.200 125.610 67.370 125.780 ;
        RECT 68.910 125.610 69.080 125.780 ;
        RECT 69.350 125.610 69.520 125.780 ;
        RECT 69.760 125.610 69.930 125.780 ;
        RECT 70.190 125.610 70.360 125.780 ;
        RECT 70.630 125.610 70.800 125.780 ;
        RECT 71.040 125.610 71.210 125.780 ;
        RECT 72.220 125.600 72.390 125.770 ;
        RECT 72.660 125.600 72.830 125.770 ;
        RECT 73.100 125.600 73.270 125.770 ;
        RECT 73.510 125.600 73.680 125.770 ;
        RECT 75.000 125.600 75.170 125.770 ;
        RECT 75.360 125.600 75.530 125.770 ;
        RECT 76.270 125.600 76.440 125.770 ;
        RECT 76.630 125.600 76.800 125.770 ;
        RECT 76.990 125.600 77.160 125.770 ;
        RECT 78.990 125.610 79.160 125.780 ;
        RECT 79.430 125.610 79.600 125.780 ;
        RECT 79.840 125.610 80.010 125.780 ;
        RECT 80.270 125.610 80.440 125.780 ;
        RECT 80.710 125.610 80.880 125.780 ;
        RECT 81.120 125.610 81.290 125.780 ;
        RECT 82.830 125.610 83.000 125.780 ;
        RECT 83.270 125.610 83.440 125.780 ;
        RECT 83.680 125.610 83.850 125.780 ;
        RECT 84.110 125.610 84.280 125.780 ;
        RECT 84.550 125.610 84.720 125.780 ;
        RECT 84.960 125.610 85.130 125.780 ;
        RECT 86.670 125.610 86.840 125.780 ;
        RECT 87.110 125.610 87.280 125.780 ;
        RECT 87.520 125.610 87.690 125.780 ;
        RECT 87.950 125.610 88.120 125.780 ;
        RECT 88.390 125.610 88.560 125.780 ;
        RECT 88.800 125.610 88.970 125.780 ;
        RECT 90.840 125.600 91.010 125.770 ;
        RECT 91.200 125.600 91.370 125.770 ;
        RECT 92.380 125.600 92.550 125.770 ;
        RECT 92.820 125.600 92.990 125.770 ;
        RECT 93.260 125.600 93.430 125.770 ;
        RECT 93.670 125.600 93.840 125.770 ;
        RECT 94.640 125.600 94.810 125.770 ;
        RECT 95.000 125.600 95.170 125.770 ;
        RECT 95.360 125.600 95.530 125.770 ;
        RECT 98.000 125.600 98.170 125.770 ;
        RECT 98.360 125.600 98.530 125.770 ;
        RECT 98.720 125.600 98.890 125.770 ;
        RECT 99.080 125.600 99.250 125.770 ;
        RECT 99.580 125.600 99.750 125.770 ;
        RECT 100.020 125.600 100.190 125.770 ;
        RECT 100.460 125.600 100.630 125.770 ;
        RECT 100.870 125.600 101.040 125.770 ;
        RECT 103.480 125.600 103.650 125.770 ;
        RECT 103.840 125.600 104.010 125.770 ;
        RECT 104.200 125.600 104.370 125.770 ;
        RECT 105.340 125.600 105.510 125.770 ;
        RECT 105.780 125.600 105.950 125.770 ;
        RECT 106.220 125.600 106.390 125.770 ;
        RECT 106.630 125.600 106.800 125.770 ;
        RECT 107.160 125.600 107.330 125.770 ;
        RECT 107.520 125.600 107.690 125.770 ;
        RECT 108.700 125.600 108.870 125.770 ;
        RECT 109.140 125.600 109.310 125.770 ;
        RECT 109.580 125.600 109.750 125.770 ;
        RECT 109.990 125.600 110.160 125.770 ;
        RECT 111.950 125.600 112.120 125.770 ;
        RECT 112.310 125.600 112.480 125.770 ;
        RECT 112.670 125.600 112.840 125.770 ;
        RECT 113.590 125.600 113.760 125.770 ;
        RECT 113.950 125.600 114.120 125.770 ;
        RECT 118.550 125.600 118.720 125.770 ;
        RECT 118.910 125.600 119.080 125.770 ;
        RECT 119.270 125.600 119.440 125.770 ;
        RECT 122.520 125.600 122.690 125.770 ;
        RECT 122.880 125.600 123.050 125.770 ;
        RECT 123.240 125.600 123.410 125.770 ;
        RECT 125.130 125.600 125.300 125.770 ;
        RECT 125.490 125.600 125.660 125.770 ;
        RECT 125.850 125.600 126.020 125.770 ;
        RECT 127.470 125.610 127.640 125.780 ;
        RECT 127.910 125.610 128.080 125.780 ;
        RECT 128.320 125.610 128.490 125.780 ;
        RECT 128.750 125.610 128.920 125.780 ;
        RECT 129.190 125.610 129.360 125.780 ;
        RECT 129.600 125.610 129.770 125.780 ;
        RECT 131.310 125.610 131.480 125.780 ;
        RECT 131.750 125.610 131.920 125.780 ;
        RECT 132.160 125.610 132.330 125.780 ;
        RECT 132.590 125.610 132.760 125.780 ;
        RECT 133.030 125.610 133.200 125.780 ;
        RECT 133.440 125.610 133.610 125.780 ;
        RECT 135.150 125.610 135.320 125.780 ;
        RECT 135.590 125.610 135.760 125.780 ;
        RECT 136.000 125.610 136.170 125.780 ;
        RECT 136.430 125.610 136.600 125.780 ;
        RECT 136.870 125.610 137.040 125.780 ;
        RECT 137.280 125.610 137.450 125.780 ;
        RECT 138.990 125.610 139.160 125.780 ;
        RECT 139.430 125.610 139.600 125.780 ;
        RECT 139.840 125.610 140.010 125.780 ;
        RECT 140.270 125.610 140.440 125.780 ;
        RECT 140.710 125.610 140.880 125.780 ;
        RECT 141.120 125.610 141.290 125.780 ;
        RECT 5.920 117.940 6.090 118.120 ;
        RECT 6.400 117.940 6.570 118.120 ;
        RECT 6.880 117.940 7.050 118.120 ;
        RECT 7.360 117.940 7.530 118.120 ;
        RECT 7.840 117.940 8.010 118.120 ;
        RECT 8.320 117.940 8.490 118.120 ;
        RECT 8.800 117.940 8.970 118.120 ;
        RECT 9.280 117.940 9.450 118.120 ;
        RECT 9.760 117.940 9.930 118.120 ;
        RECT 10.240 117.940 10.410 118.120 ;
      LAYER li1 ;
        RECT 10.560 117.940 11.040 118.120 ;
      LAYER li1 ;
        RECT 11.200 117.940 11.370 118.120 ;
        RECT 11.680 117.940 11.850 118.120 ;
        RECT 12.160 117.940 12.330 118.120 ;
        RECT 12.640 117.940 12.810 118.120 ;
        RECT 13.120 117.940 13.290 118.120 ;
        RECT 13.600 117.940 13.770 118.120 ;
        RECT 14.080 117.940 14.250 118.120 ;
        RECT 14.560 117.940 14.730 118.120 ;
        RECT 15.040 117.940 15.210 118.120 ;
        RECT 15.520 117.940 15.690 118.120 ;
        RECT 16.000 117.940 16.170 118.120 ;
        RECT 16.480 117.940 16.650 118.120 ;
        RECT 16.960 117.940 17.130 118.120 ;
        RECT 17.440 117.940 17.610 118.120 ;
        RECT 17.920 117.940 18.090 118.120 ;
        RECT 18.400 117.940 18.570 118.120 ;
        RECT 18.880 117.940 19.050 118.120 ;
        RECT 19.360 117.940 19.530 118.120 ;
        RECT 19.840 117.940 20.010 118.120 ;
        RECT 20.320 117.940 20.490 118.120 ;
        RECT 20.800 117.940 20.970 118.120 ;
        RECT 21.280 117.940 21.450 118.120 ;
        RECT 21.760 117.940 21.930 118.120 ;
        RECT 22.240 117.940 22.410 118.120 ;
        RECT 22.720 117.940 22.890 118.120 ;
        RECT 23.200 117.940 23.370 118.120 ;
        RECT 23.680 117.940 23.850 118.120 ;
        RECT 24.160 117.940 24.330 118.120 ;
        RECT 24.640 117.940 24.810 118.120 ;
        RECT 25.120 117.940 25.290 118.120 ;
        RECT 25.600 117.940 25.770 118.120 ;
        RECT 26.080 117.940 26.250 118.120 ;
        RECT 26.560 117.940 26.730 118.120 ;
        RECT 27.040 117.940 27.210 118.120 ;
        RECT 27.520 117.940 27.690 118.120 ;
        RECT 28.000 117.940 28.170 118.120 ;
      LAYER li1 ;
        RECT 28.320 117.940 28.800 118.120 ;
      LAYER li1 ;
        RECT 28.960 117.940 29.130 118.120 ;
        RECT 29.440 117.940 29.610 118.120 ;
        RECT 29.920 117.940 30.090 118.120 ;
        RECT 30.400 117.940 30.570 118.120 ;
        RECT 30.880 117.940 31.050 118.120 ;
        RECT 31.360 117.940 31.530 118.120 ;
        RECT 31.840 117.940 32.010 118.120 ;
        RECT 32.320 117.940 32.490 118.120 ;
        RECT 32.800 117.940 32.970 118.120 ;
        RECT 33.280 117.940 33.450 118.120 ;
        RECT 33.760 117.940 33.930 118.120 ;
        RECT 34.240 117.940 34.410 118.120 ;
        RECT 34.720 117.940 34.890 118.120 ;
        RECT 35.200 117.940 35.370 118.120 ;
        RECT 35.680 117.940 35.850 118.120 ;
        RECT 36.160 117.940 36.330 118.120 ;
        RECT 36.640 117.940 36.810 118.120 ;
        RECT 37.120 117.940 37.290 118.120 ;
        RECT 37.600 117.940 37.770 118.120 ;
        RECT 38.080 117.940 38.250 118.120 ;
        RECT 38.560 117.940 38.730 118.120 ;
        RECT 39.040 117.940 39.210 118.120 ;
        RECT 39.520 117.940 39.690 118.120 ;
        RECT 40.000 117.940 40.170 118.120 ;
        RECT 40.480 117.940 40.650 118.120 ;
        RECT 40.960 117.940 41.130 118.120 ;
        RECT 41.440 117.940 41.610 118.120 ;
        RECT 41.920 117.940 42.090 118.120 ;
        RECT 42.400 117.940 42.570 118.120 ;
        RECT 42.880 117.940 43.050 118.120 ;
      LAYER li1 ;
        RECT 43.200 117.940 43.680 118.120 ;
      LAYER li1 ;
        RECT 43.840 117.940 44.010 118.120 ;
        RECT 44.320 117.940 44.490 118.120 ;
        RECT 44.800 117.940 44.970 118.120 ;
        RECT 45.280 117.940 45.450 118.120 ;
        RECT 45.760 117.940 45.930 118.120 ;
        RECT 46.240 117.940 46.410 118.120 ;
        RECT 46.720 117.940 46.890 118.120 ;
        RECT 47.200 117.940 47.370 118.120 ;
        RECT 47.680 117.940 47.850 118.120 ;
        RECT 48.160 117.940 48.330 118.120 ;
        RECT 48.640 117.940 48.810 118.120 ;
        RECT 49.120 117.940 49.290 118.120 ;
        RECT 49.600 117.940 49.770 118.120 ;
      LAYER li1 ;
        RECT 49.920 117.940 50.400 118.120 ;
      LAYER li1 ;
        RECT 50.560 117.940 50.730 118.120 ;
        RECT 51.040 117.940 51.210 118.120 ;
        RECT 51.520 117.940 51.690 118.120 ;
        RECT 52.000 117.940 52.170 118.120 ;
        RECT 52.480 117.940 52.650 118.120 ;
        RECT 52.960 117.940 53.130 118.120 ;
        RECT 53.440 117.940 53.610 118.120 ;
        RECT 53.920 117.940 54.090 118.120 ;
        RECT 54.400 117.940 54.570 118.120 ;
        RECT 54.880 117.940 55.050 118.120 ;
        RECT 55.360 117.940 55.530 118.120 ;
        RECT 55.840 117.940 56.010 118.120 ;
        RECT 56.320 117.940 56.490 118.120 ;
        RECT 56.800 117.940 56.970 118.120 ;
        RECT 57.280 117.940 57.450 118.120 ;
        RECT 57.760 117.940 57.930 118.120 ;
        RECT 58.240 117.940 58.410 118.120 ;
        RECT 58.720 117.940 58.890 118.120 ;
        RECT 59.200 117.940 59.370 118.120 ;
        RECT 59.680 117.940 59.850 118.120 ;
        RECT 60.160 117.940 60.330 118.120 ;
        RECT 60.640 117.940 60.810 118.120 ;
        RECT 61.120 117.940 61.290 118.120 ;
        RECT 61.600 117.940 61.770 118.120 ;
        RECT 62.080 117.940 62.250 118.120 ;
        RECT 62.560 117.940 62.730 118.120 ;
        RECT 63.040 117.940 63.210 118.120 ;
        RECT 63.520 117.940 63.690 118.120 ;
        RECT 64.000 117.940 64.170 118.120 ;
        RECT 64.480 117.940 64.650 118.120 ;
        RECT 64.960 117.940 65.130 118.120 ;
        RECT 65.440 117.940 65.610 118.120 ;
        RECT 65.920 117.940 66.090 118.120 ;
        RECT 66.400 117.940 66.570 118.120 ;
        RECT 66.880 117.940 67.050 118.120 ;
      LAYER li1 ;
        RECT 67.200 117.940 67.680 118.120 ;
      LAYER li1 ;
        RECT 67.840 117.940 68.010 118.120 ;
        RECT 68.320 117.940 68.490 118.120 ;
        RECT 68.800 117.940 68.970 118.120 ;
        RECT 69.280 117.940 69.450 118.120 ;
        RECT 69.760 117.940 69.930 118.120 ;
        RECT 70.240 117.940 70.410 118.120 ;
        RECT 70.720 117.940 70.890 118.120 ;
        RECT 71.200 117.940 71.370 118.120 ;
        RECT 71.680 117.940 71.850 118.120 ;
        RECT 72.160 117.940 72.330 118.120 ;
        RECT 72.640 117.940 72.810 118.120 ;
        RECT 73.120 117.940 73.290 118.120 ;
        RECT 73.600 117.940 73.770 118.120 ;
        RECT 74.080 117.940 74.250 118.120 ;
        RECT 74.560 117.940 74.730 118.120 ;
        RECT 75.040 117.940 75.210 118.120 ;
        RECT 75.520 117.940 75.690 118.120 ;
        RECT 76.000 117.940 76.170 118.120 ;
        RECT 76.480 117.940 76.650 118.120 ;
        RECT 76.960 117.940 77.130 118.120 ;
        RECT 77.440 117.940 77.610 118.120 ;
        RECT 77.920 117.940 78.090 118.120 ;
        RECT 78.400 117.940 78.570 118.120 ;
        RECT 78.880 117.940 79.050 118.120 ;
        RECT 79.360 117.940 79.530 118.120 ;
        RECT 79.840 117.940 80.010 118.120 ;
        RECT 80.320 117.940 80.490 118.120 ;
        RECT 80.800 117.940 80.970 118.120 ;
        RECT 81.280 117.940 81.450 118.120 ;
        RECT 81.760 117.940 81.930 118.120 ;
        RECT 82.240 117.940 82.410 118.120 ;
        RECT 82.720 117.940 82.890 118.120 ;
        RECT 83.200 117.940 83.370 118.120 ;
        RECT 83.680 117.940 83.850 118.120 ;
        RECT 84.160 117.940 84.330 118.120 ;
        RECT 84.640 117.940 84.810 118.120 ;
        RECT 85.120 117.940 85.290 118.120 ;
        RECT 85.600 117.940 85.770 118.120 ;
        RECT 86.080 117.940 86.250 118.120 ;
        RECT 86.560 117.940 86.730 118.120 ;
        RECT 87.040 117.940 87.210 118.120 ;
        RECT 87.520 117.940 87.690 118.120 ;
        RECT 88.000 117.940 88.170 118.120 ;
        RECT 88.480 117.940 88.650 118.120 ;
        RECT 88.960 117.940 89.130 118.120 ;
        RECT 89.440 117.940 89.610 118.120 ;
        RECT 89.920 117.940 90.090 118.120 ;
        RECT 90.400 117.940 90.570 118.120 ;
        RECT 90.880 117.940 91.050 118.120 ;
        RECT 91.360 117.940 91.530 118.120 ;
        RECT 91.840 117.940 92.010 118.120 ;
        RECT 92.320 117.940 92.490 118.120 ;
        RECT 92.800 117.940 92.970 118.120 ;
        RECT 93.280 117.940 93.450 118.120 ;
        RECT 93.760 117.940 93.930 118.120 ;
        RECT 94.240 117.940 94.410 118.120 ;
        RECT 94.720 117.940 94.890 118.120 ;
        RECT 95.200 117.940 95.370 118.120 ;
        RECT 95.680 117.940 95.850 118.120 ;
        RECT 96.160 117.940 96.330 118.120 ;
        RECT 96.640 117.940 96.810 118.120 ;
        RECT 97.120 117.940 97.290 118.120 ;
        RECT 97.600 117.940 97.770 118.120 ;
        RECT 98.080 117.940 98.250 118.120 ;
        RECT 98.560 117.940 98.730 118.120 ;
        RECT 99.040 117.940 99.210 118.120 ;
        RECT 99.520 117.940 99.690 118.120 ;
        RECT 100.000 117.940 100.170 118.120 ;
      LAYER li1 ;
        RECT 100.320 117.940 100.800 118.120 ;
      LAYER li1 ;
        RECT 100.960 117.940 101.130 118.120 ;
        RECT 101.440 117.940 101.610 118.120 ;
        RECT 101.920 117.940 102.090 118.120 ;
        RECT 102.400 117.940 102.570 118.120 ;
        RECT 102.880 117.940 103.050 118.120 ;
        RECT 103.360 117.940 103.530 118.120 ;
        RECT 103.840 117.940 104.010 118.120 ;
        RECT 104.320 117.940 104.490 118.120 ;
        RECT 104.800 117.940 104.970 118.120 ;
        RECT 105.280 117.940 105.450 118.120 ;
        RECT 105.760 117.940 105.930 118.120 ;
        RECT 106.240 117.940 106.410 118.120 ;
        RECT 106.720 117.940 106.890 118.120 ;
        RECT 107.200 117.940 107.370 118.120 ;
        RECT 107.680 117.940 107.850 118.120 ;
        RECT 108.160 117.940 108.330 118.120 ;
        RECT 108.640 117.940 108.810 118.120 ;
        RECT 109.120 117.940 109.290 118.120 ;
        RECT 109.600 117.940 109.770 118.120 ;
        RECT 110.080 117.940 110.250 118.120 ;
        RECT 110.560 117.940 110.730 118.120 ;
        RECT 111.040 117.940 111.210 118.120 ;
        RECT 111.520 117.940 111.690 118.120 ;
        RECT 112.000 117.940 112.170 118.120 ;
        RECT 112.480 117.940 112.650 118.120 ;
        RECT 112.960 117.940 113.130 118.120 ;
        RECT 113.440 117.940 113.610 118.120 ;
        RECT 113.920 117.940 114.090 118.120 ;
        RECT 114.400 117.940 114.570 118.120 ;
        RECT 114.880 117.940 115.050 118.120 ;
        RECT 115.360 117.940 115.530 118.120 ;
        RECT 115.840 117.940 116.010 118.120 ;
        RECT 116.320 117.940 116.490 118.120 ;
        RECT 116.800 117.940 116.970 118.120 ;
        RECT 117.280 117.940 117.450 118.120 ;
        RECT 117.760 117.940 117.930 118.120 ;
        RECT 118.240 117.940 118.410 118.120 ;
        RECT 118.720 117.940 118.890 118.120 ;
        RECT 119.200 117.940 119.370 118.120 ;
        RECT 119.680 117.940 119.850 118.120 ;
        RECT 120.160 117.940 120.330 118.120 ;
        RECT 120.640 117.940 120.810 118.120 ;
        RECT 121.120 117.940 121.290 118.120 ;
        RECT 121.600 117.940 121.770 118.120 ;
        RECT 122.080 117.940 122.250 118.120 ;
        RECT 122.560 117.940 122.730 118.120 ;
        RECT 123.040 117.940 123.210 118.120 ;
        RECT 123.520 117.940 123.690 118.120 ;
        RECT 124.000 117.940 124.170 118.120 ;
        RECT 124.480 117.940 124.650 118.120 ;
        RECT 124.960 117.940 125.130 118.120 ;
        RECT 125.440 117.940 125.610 118.120 ;
        RECT 125.920 117.940 126.090 118.120 ;
        RECT 126.400 117.940 126.570 118.120 ;
        RECT 126.880 117.940 127.050 118.120 ;
        RECT 127.360 117.940 127.530 118.120 ;
        RECT 127.840 117.940 128.010 118.120 ;
        RECT 128.320 117.940 128.490 118.120 ;
        RECT 128.800 117.940 128.970 118.120 ;
        RECT 129.280 117.940 129.450 118.120 ;
        RECT 129.760 117.940 129.930 118.120 ;
        RECT 130.240 117.940 130.410 118.120 ;
        RECT 130.720 117.940 130.890 118.120 ;
        RECT 131.200 117.940 131.370 118.120 ;
        RECT 131.680 117.940 131.850 118.120 ;
        RECT 132.160 117.940 132.330 118.120 ;
        RECT 132.640 117.940 132.810 118.120 ;
        RECT 133.120 117.940 133.290 118.120 ;
        RECT 133.600 117.940 133.770 118.120 ;
        RECT 134.080 117.940 134.250 118.120 ;
        RECT 134.560 117.940 134.730 118.120 ;
        RECT 135.040 117.940 135.210 118.120 ;
        RECT 135.520 117.940 135.690 118.120 ;
        RECT 136.000 117.940 136.170 118.120 ;
        RECT 136.480 117.940 136.650 118.120 ;
        RECT 136.960 117.940 137.130 118.120 ;
        RECT 137.440 117.940 137.610 118.120 ;
        RECT 137.920 117.940 138.090 118.120 ;
        RECT 138.400 117.940 138.570 118.120 ;
        RECT 138.880 117.940 139.050 118.120 ;
        RECT 139.360 117.940 139.530 118.120 ;
        RECT 139.840 117.940 140.010 118.120 ;
        RECT 140.320 117.940 140.490 118.120 ;
        RECT 140.800 117.940 140.970 118.120 ;
        RECT 141.280 117.940 141.450 118.120 ;
      LAYER li1 ;
        RECT 141.600 117.940 142.080 118.120 ;
      LAYER li1 ;
        RECT 6.510 117.470 6.680 117.640 ;
        RECT 6.950 117.470 7.120 117.640 ;
        RECT 7.360 117.470 7.530 117.640 ;
        RECT 7.790 117.470 7.960 117.640 ;
        RECT 8.230 117.470 8.400 117.640 ;
        RECT 8.640 117.470 8.810 117.640 ;
        RECT 10.350 117.470 10.520 117.640 ;
        RECT 10.790 117.470 10.960 117.640 ;
        RECT 11.200 117.470 11.370 117.640 ;
        RECT 11.630 117.470 11.800 117.640 ;
        RECT 12.070 117.470 12.240 117.640 ;
        RECT 12.480 117.470 12.650 117.640 ;
        RECT 14.470 117.460 14.640 117.630 ;
        RECT 14.830 117.460 15.000 117.630 ;
        RECT 15.190 117.460 15.360 117.630 ;
        RECT 15.550 117.460 15.720 117.630 ;
        RECT 17.070 117.470 17.240 117.640 ;
        RECT 17.510 117.470 17.680 117.640 ;
        RECT 17.920 117.470 18.090 117.640 ;
        RECT 18.350 117.470 18.520 117.640 ;
        RECT 18.790 117.470 18.960 117.640 ;
        RECT 19.200 117.470 19.370 117.640 ;
        RECT 20.910 117.470 21.080 117.640 ;
        RECT 21.350 117.470 21.520 117.640 ;
        RECT 21.760 117.470 21.930 117.640 ;
        RECT 22.190 117.470 22.360 117.640 ;
        RECT 22.630 117.470 22.800 117.640 ;
        RECT 23.040 117.470 23.210 117.640 ;
        RECT 25.080 117.460 25.250 117.630 ;
        RECT 25.440 117.460 25.610 117.630 ;
        RECT 27.150 117.470 27.320 117.640 ;
        RECT 27.590 117.470 27.760 117.640 ;
        RECT 28.000 117.470 28.170 117.640 ;
        RECT 28.430 117.470 28.600 117.640 ;
        RECT 28.870 117.470 29.040 117.640 ;
        RECT 29.280 117.470 29.450 117.640 ;
        RECT 30.990 117.470 31.160 117.640 ;
        RECT 31.430 117.470 31.600 117.640 ;
        RECT 31.840 117.470 32.010 117.640 ;
        RECT 32.270 117.470 32.440 117.640 ;
        RECT 32.710 117.470 32.880 117.640 ;
        RECT 33.120 117.470 33.290 117.640 ;
        RECT 34.830 117.470 35.000 117.640 ;
        RECT 35.270 117.470 35.440 117.640 ;
        RECT 35.680 117.470 35.850 117.640 ;
        RECT 36.110 117.470 36.280 117.640 ;
        RECT 36.550 117.470 36.720 117.640 ;
        RECT 36.960 117.470 37.130 117.640 ;
        RECT 38.670 117.470 38.840 117.640 ;
        RECT 39.110 117.470 39.280 117.640 ;
        RECT 39.520 117.470 39.690 117.640 ;
        RECT 39.950 117.470 40.120 117.640 ;
        RECT 40.390 117.470 40.560 117.640 ;
        RECT 40.800 117.470 40.970 117.640 ;
        RECT 44.920 117.460 45.090 117.630 ;
        RECT 45.280 117.460 45.450 117.630 ;
        RECT 45.640 117.460 45.810 117.630 ;
        RECT 46.780 117.460 46.950 117.630 ;
        RECT 47.220 117.460 47.390 117.630 ;
        RECT 47.660 117.460 47.830 117.630 ;
        RECT 48.070 117.460 48.240 117.630 ;
        RECT 48.600 117.460 48.770 117.630 ;
        RECT 48.960 117.460 49.130 117.630 ;
        RECT 49.320 117.460 49.490 117.630 ;
        RECT 50.160 117.460 50.330 117.630 ;
        RECT 50.520 117.460 50.690 117.630 ;
        RECT 50.880 117.460 51.050 117.630 ;
        RECT 51.720 117.460 51.890 117.630 ;
        RECT 52.080 117.460 52.250 117.630 ;
        RECT 52.440 117.460 52.610 117.630 ;
        RECT 53.500 117.460 53.670 117.630 ;
        RECT 53.940 117.460 54.110 117.630 ;
        RECT 54.380 117.460 54.550 117.630 ;
        RECT 54.790 117.460 54.960 117.630 ;
        RECT 56.710 117.460 56.880 117.630 ;
        RECT 57.070 117.460 57.240 117.630 ;
        RECT 57.430 117.460 57.600 117.630 ;
        RECT 57.790 117.460 57.960 117.630 ;
        RECT 58.780 117.460 58.950 117.630 ;
        RECT 59.220 117.460 59.390 117.630 ;
        RECT 59.660 117.460 59.830 117.630 ;
        RECT 60.070 117.460 60.240 117.630 ;
        RECT 61.030 117.460 61.200 117.630 ;
        RECT 61.390 117.460 61.560 117.630 ;
        RECT 61.750 117.460 61.920 117.630 ;
        RECT 62.110 117.460 62.280 117.630 ;
        RECT 63.630 117.470 63.800 117.640 ;
        RECT 64.070 117.470 64.240 117.640 ;
        RECT 64.480 117.470 64.650 117.640 ;
        RECT 64.910 117.470 65.080 117.640 ;
        RECT 65.350 117.470 65.520 117.640 ;
        RECT 65.760 117.470 65.930 117.640 ;
        RECT 67.270 117.460 67.440 117.630 ;
        RECT 67.630 117.460 67.800 117.630 ;
        RECT 67.990 117.460 68.160 117.630 ;
        RECT 68.350 117.460 68.520 117.630 ;
        RECT 69.340 117.460 69.510 117.630 ;
        RECT 69.780 117.460 69.950 117.630 ;
        RECT 70.220 117.460 70.390 117.630 ;
        RECT 70.630 117.460 70.800 117.630 ;
        RECT 71.630 117.460 71.800 117.630 ;
        RECT 71.990 117.460 72.160 117.630 ;
        RECT 72.350 117.460 72.520 117.630 ;
        RECT 73.270 117.460 73.440 117.630 ;
        RECT 73.630 117.460 73.800 117.630 ;
        RECT 78.230 117.460 78.400 117.630 ;
        RECT 78.590 117.460 78.760 117.630 ;
        RECT 78.950 117.460 79.120 117.630 ;
        RECT 82.200 117.460 82.370 117.630 ;
        RECT 82.560 117.460 82.730 117.630 ;
        RECT 82.920 117.460 83.090 117.630 ;
        RECT 84.810 117.460 84.980 117.630 ;
        RECT 85.170 117.460 85.340 117.630 ;
        RECT 85.530 117.460 85.700 117.630 ;
        RECT 86.620 117.460 86.790 117.630 ;
        RECT 87.060 117.460 87.230 117.630 ;
        RECT 87.500 117.460 87.670 117.630 ;
        RECT 87.910 117.460 88.080 117.630 ;
        RECT 89.350 117.460 89.520 117.630 ;
        RECT 89.710 117.460 89.880 117.630 ;
        RECT 90.070 117.460 90.240 117.630 ;
        RECT 90.430 117.460 90.600 117.630 ;
        RECT 91.420 117.460 91.590 117.630 ;
        RECT 91.860 117.460 92.030 117.630 ;
        RECT 92.300 117.460 92.470 117.630 ;
        RECT 92.710 117.460 92.880 117.630 ;
        RECT 93.680 117.460 93.850 117.630 ;
        RECT 94.040 117.460 94.210 117.630 ;
        RECT 94.400 117.460 94.570 117.630 ;
        RECT 97.040 117.460 97.210 117.630 ;
        RECT 97.400 117.460 97.570 117.630 ;
        RECT 97.760 117.460 97.930 117.630 ;
        RECT 98.120 117.460 98.290 117.630 ;
        RECT 98.620 117.460 98.790 117.630 ;
        RECT 99.060 117.460 99.230 117.630 ;
        RECT 99.500 117.460 99.670 117.630 ;
        RECT 99.910 117.460 100.080 117.630 ;
        RECT 100.870 117.460 101.040 117.630 ;
        RECT 101.230 117.460 101.400 117.630 ;
        RECT 101.590 117.460 101.760 117.630 ;
        RECT 101.950 117.460 102.120 117.630 ;
        RECT 102.940 117.460 103.110 117.630 ;
        RECT 103.380 117.460 103.550 117.630 ;
        RECT 103.820 117.460 103.990 117.630 ;
        RECT 104.230 117.460 104.400 117.630 ;
        RECT 104.760 117.460 104.930 117.630 ;
        RECT 105.120 117.460 105.290 117.630 ;
        RECT 105.480 117.460 105.650 117.630 ;
        RECT 106.320 117.460 106.490 117.630 ;
        RECT 106.680 117.460 106.850 117.630 ;
        RECT 107.040 117.460 107.210 117.630 ;
        RECT 107.880 117.460 108.050 117.630 ;
        RECT 108.240 117.460 108.410 117.630 ;
        RECT 108.600 117.460 108.770 117.630 ;
        RECT 109.660 117.460 109.830 117.630 ;
        RECT 110.100 117.460 110.270 117.630 ;
        RECT 110.540 117.460 110.710 117.630 ;
        RECT 110.950 117.460 111.120 117.630 ;
        RECT 111.910 117.460 112.080 117.630 ;
        RECT 112.270 117.460 112.440 117.630 ;
        RECT 112.630 117.460 112.800 117.630 ;
        RECT 112.990 117.460 113.160 117.630 ;
        RECT 113.980 117.460 114.150 117.630 ;
        RECT 114.420 117.460 114.590 117.630 ;
        RECT 114.860 117.460 115.030 117.630 ;
        RECT 115.270 117.460 115.440 117.630 ;
        RECT 117.670 117.460 117.840 117.630 ;
        RECT 118.030 117.460 118.200 117.630 ;
        RECT 118.390 117.460 118.560 117.630 ;
        RECT 118.750 117.460 118.920 117.630 ;
        RECT 119.740 117.460 119.910 117.630 ;
        RECT 120.180 117.460 120.350 117.630 ;
        RECT 120.620 117.460 120.790 117.630 ;
        RECT 121.030 117.460 121.200 117.630 ;
        RECT 121.560 117.460 121.730 117.630 ;
        RECT 121.920 117.460 122.090 117.630 ;
        RECT 123.630 117.470 123.800 117.640 ;
        RECT 124.070 117.470 124.240 117.640 ;
        RECT 124.480 117.470 124.650 117.640 ;
        RECT 124.910 117.470 125.080 117.640 ;
        RECT 125.350 117.470 125.520 117.640 ;
        RECT 125.760 117.470 125.930 117.640 ;
        RECT 127.470 117.470 127.640 117.640 ;
        RECT 127.910 117.470 128.080 117.640 ;
        RECT 128.320 117.470 128.490 117.640 ;
        RECT 128.750 117.470 128.920 117.640 ;
        RECT 129.190 117.470 129.360 117.640 ;
        RECT 129.600 117.470 129.770 117.640 ;
        RECT 131.310 117.470 131.480 117.640 ;
        RECT 131.750 117.470 131.920 117.640 ;
        RECT 132.160 117.470 132.330 117.640 ;
        RECT 132.590 117.470 132.760 117.640 ;
        RECT 133.030 117.470 133.200 117.640 ;
        RECT 133.440 117.470 133.610 117.640 ;
        RECT 135.150 117.470 135.320 117.640 ;
        RECT 135.590 117.470 135.760 117.640 ;
        RECT 136.000 117.470 136.170 117.640 ;
        RECT 136.430 117.470 136.600 117.640 ;
        RECT 136.870 117.470 137.040 117.640 ;
        RECT 137.280 117.470 137.450 117.640 ;
        RECT 138.990 117.470 139.160 117.640 ;
        RECT 139.430 117.470 139.600 117.640 ;
        RECT 139.840 117.470 140.010 117.640 ;
        RECT 140.270 117.470 140.440 117.640 ;
        RECT 140.710 117.470 140.880 117.640 ;
        RECT 141.120 117.470 141.290 117.640 ;
        RECT 5.920 109.800 6.090 109.980 ;
        RECT 6.400 109.800 6.570 109.980 ;
        RECT 6.880 109.800 7.050 109.980 ;
        RECT 7.360 109.800 7.530 109.980 ;
        RECT 7.840 109.800 8.010 109.980 ;
        RECT 8.320 109.800 8.490 109.980 ;
        RECT 8.800 109.800 8.970 109.980 ;
        RECT 9.280 109.800 9.450 109.980 ;
        RECT 9.760 109.800 9.930 109.980 ;
        RECT 10.240 109.800 10.410 109.980 ;
        RECT 10.720 109.800 10.890 109.980 ;
        RECT 11.200 109.800 11.370 109.980 ;
        RECT 11.680 109.800 11.850 109.980 ;
        RECT 12.160 109.800 12.330 109.980 ;
        RECT 12.640 109.800 12.810 109.980 ;
        RECT 13.120 109.800 13.290 109.980 ;
        RECT 13.600 109.800 13.770 109.980 ;
        RECT 14.080 109.800 14.250 109.980 ;
        RECT 14.560 109.800 14.730 109.980 ;
        RECT 15.040 109.800 15.210 109.980 ;
        RECT 15.520 109.800 15.690 109.980 ;
        RECT 16.000 109.800 16.170 109.980 ;
        RECT 16.480 109.800 16.650 109.980 ;
        RECT 16.960 109.800 17.130 109.980 ;
        RECT 17.440 109.800 17.610 109.980 ;
        RECT 17.920 109.800 18.090 109.980 ;
        RECT 18.400 109.800 18.570 109.980 ;
        RECT 18.880 109.800 19.050 109.980 ;
        RECT 19.360 109.800 19.530 109.980 ;
        RECT 19.840 109.800 20.010 109.980 ;
        RECT 20.320 109.800 20.490 109.980 ;
        RECT 20.800 109.800 20.970 109.980 ;
        RECT 21.280 109.800 21.450 109.980 ;
        RECT 21.760 109.800 21.930 109.980 ;
        RECT 22.240 109.800 22.410 109.980 ;
        RECT 22.720 109.800 22.890 109.980 ;
        RECT 23.200 109.800 23.370 109.980 ;
        RECT 23.680 109.800 23.850 109.980 ;
      LAYER li1 ;
        RECT 24.000 109.800 24.480 109.980 ;
      LAYER li1 ;
        RECT 24.640 109.800 24.810 109.980 ;
        RECT 25.120 109.800 25.290 109.980 ;
        RECT 25.600 109.800 25.770 109.980 ;
        RECT 26.080 109.800 26.250 109.980 ;
        RECT 26.560 109.800 26.730 109.980 ;
        RECT 27.040 109.800 27.210 109.980 ;
        RECT 27.520 109.800 27.690 109.980 ;
        RECT 28.000 109.800 28.170 109.980 ;
        RECT 28.480 109.800 28.650 109.980 ;
        RECT 28.960 109.800 29.130 109.980 ;
        RECT 29.440 109.800 29.610 109.980 ;
        RECT 29.920 109.800 30.090 109.980 ;
        RECT 30.400 109.800 30.570 109.980 ;
        RECT 30.880 109.800 31.050 109.980 ;
        RECT 31.360 109.800 31.530 109.980 ;
        RECT 31.840 109.800 32.010 109.980 ;
        RECT 32.320 109.800 32.490 109.980 ;
        RECT 32.800 109.800 32.970 109.980 ;
        RECT 33.280 109.800 33.450 109.980 ;
        RECT 33.760 109.800 33.930 109.980 ;
        RECT 34.240 109.800 34.410 109.980 ;
        RECT 34.720 109.800 34.890 109.980 ;
        RECT 35.200 109.800 35.370 109.980 ;
        RECT 35.680 109.800 35.850 109.980 ;
        RECT 36.160 109.800 36.330 109.980 ;
        RECT 36.640 109.800 36.810 109.980 ;
      LAYER li1 ;
        RECT 36.960 109.800 37.440 109.980 ;
      LAYER li1 ;
        RECT 37.600 109.800 37.770 109.980 ;
        RECT 38.080 109.800 38.250 109.980 ;
        RECT 38.560 109.800 38.730 109.980 ;
        RECT 39.040 109.800 39.210 109.980 ;
        RECT 39.520 109.800 39.690 109.980 ;
        RECT 40.000 109.800 40.170 109.980 ;
        RECT 40.480 109.800 40.650 109.980 ;
        RECT 40.960 109.800 41.130 109.980 ;
        RECT 41.440 109.800 41.610 109.980 ;
        RECT 41.920 109.800 42.090 109.980 ;
        RECT 42.400 109.800 42.570 109.980 ;
        RECT 42.880 109.800 43.050 109.980 ;
        RECT 43.360 109.800 43.530 109.980 ;
        RECT 43.840 109.800 44.010 109.980 ;
        RECT 44.320 109.800 44.490 109.980 ;
        RECT 44.800 109.800 44.970 109.980 ;
        RECT 45.280 109.800 45.450 109.980 ;
        RECT 45.760 109.800 45.930 109.980 ;
        RECT 46.240 109.800 46.410 109.980 ;
        RECT 46.720 109.800 46.890 109.980 ;
        RECT 47.200 109.800 47.370 109.980 ;
        RECT 47.680 109.800 47.850 109.980 ;
        RECT 48.160 109.800 48.330 109.980 ;
        RECT 48.640 109.800 48.810 109.980 ;
        RECT 49.120 109.800 49.290 109.980 ;
        RECT 49.600 109.800 49.770 109.980 ;
        RECT 50.080 109.800 50.250 109.980 ;
        RECT 50.560 109.800 50.730 109.980 ;
        RECT 51.040 109.800 51.210 109.980 ;
        RECT 51.520 109.800 51.690 109.980 ;
        RECT 52.000 109.800 52.170 109.980 ;
        RECT 52.480 109.800 52.650 109.980 ;
        RECT 52.960 109.800 53.130 109.980 ;
        RECT 53.440 109.800 53.610 109.980 ;
        RECT 53.920 109.800 54.090 109.980 ;
        RECT 54.400 109.800 54.570 109.980 ;
        RECT 54.880 109.800 55.050 109.980 ;
        RECT 55.360 109.800 55.530 109.980 ;
        RECT 55.840 109.800 56.010 109.980 ;
        RECT 56.320 109.800 56.490 109.980 ;
        RECT 56.800 109.800 56.970 109.980 ;
        RECT 57.280 109.800 57.450 109.980 ;
        RECT 57.760 109.800 57.930 109.980 ;
        RECT 58.240 109.800 58.410 109.980 ;
        RECT 58.720 109.800 58.890 109.980 ;
        RECT 59.200 109.800 59.370 109.980 ;
        RECT 59.680 109.800 59.850 109.980 ;
        RECT 60.160 109.800 60.330 109.980 ;
        RECT 60.640 109.800 60.810 109.980 ;
        RECT 61.120 109.800 61.290 109.980 ;
        RECT 61.600 109.800 61.770 109.980 ;
        RECT 62.080 109.800 62.250 109.980 ;
        RECT 62.560 109.800 62.730 109.980 ;
        RECT 63.040 109.800 63.210 109.980 ;
        RECT 63.520 109.800 63.690 109.980 ;
        RECT 64.000 109.800 64.170 109.980 ;
        RECT 64.480 109.800 64.650 109.980 ;
        RECT 64.960 109.800 65.130 109.980 ;
        RECT 65.440 109.800 65.610 109.980 ;
        RECT 65.920 109.800 66.090 109.980 ;
        RECT 66.400 109.800 66.570 109.980 ;
        RECT 66.880 109.800 67.050 109.980 ;
        RECT 67.360 109.800 67.530 109.980 ;
        RECT 67.840 109.800 68.010 109.980 ;
        RECT 68.320 109.800 68.490 109.980 ;
        RECT 68.800 109.800 68.970 109.980 ;
        RECT 69.280 109.800 69.450 109.980 ;
        RECT 69.760 109.800 69.930 109.980 ;
        RECT 70.240 109.800 70.410 109.980 ;
        RECT 70.720 109.800 70.890 109.980 ;
        RECT 71.200 109.800 71.370 109.980 ;
      LAYER li1 ;
        RECT 71.520 109.800 72.000 109.980 ;
      LAYER li1 ;
        RECT 72.160 109.800 72.330 109.980 ;
        RECT 72.640 109.800 72.810 109.980 ;
        RECT 73.120 109.800 73.290 109.980 ;
        RECT 73.600 109.800 73.770 109.980 ;
        RECT 74.080 109.800 74.250 109.980 ;
        RECT 74.560 109.800 74.730 109.980 ;
        RECT 75.040 109.800 75.210 109.980 ;
        RECT 75.520 109.800 75.690 109.980 ;
        RECT 76.000 109.800 76.170 109.980 ;
        RECT 76.480 109.800 76.650 109.980 ;
        RECT 76.960 109.800 77.130 109.980 ;
        RECT 77.440 109.800 77.610 109.980 ;
        RECT 77.920 109.800 78.090 109.980 ;
        RECT 78.400 109.800 78.570 109.980 ;
        RECT 78.880 109.800 79.050 109.980 ;
        RECT 79.360 109.800 79.530 109.980 ;
        RECT 79.840 109.800 80.010 109.980 ;
        RECT 80.320 109.800 80.490 109.980 ;
        RECT 80.800 109.800 80.970 109.980 ;
        RECT 81.280 109.800 81.450 109.980 ;
        RECT 81.760 109.800 81.930 109.980 ;
        RECT 82.240 109.800 82.410 109.980 ;
        RECT 82.720 109.800 82.890 109.980 ;
        RECT 83.200 109.800 83.370 109.980 ;
        RECT 83.680 109.800 83.850 109.980 ;
        RECT 84.160 109.800 84.330 109.980 ;
        RECT 84.640 109.800 84.810 109.980 ;
        RECT 85.120 109.800 85.290 109.980 ;
        RECT 85.600 109.800 85.770 109.980 ;
        RECT 86.080 109.800 86.250 109.980 ;
        RECT 86.560 109.800 86.730 109.980 ;
        RECT 87.040 109.800 87.210 109.980 ;
        RECT 87.520 109.800 87.690 109.980 ;
        RECT 88.000 109.800 88.170 109.980 ;
        RECT 88.480 109.800 88.650 109.980 ;
        RECT 88.960 109.800 89.130 109.980 ;
        RECT 89.440 109.800 89.610 109.980 ;
        RECT 89.920 109.800 90.090 109.980 ;
        RECT 90.400 109.800 90.570 109.980 ;
        RECT 90.880 109.800 91.050 109.980 ;
        RECT 91.360 109.800 91.530 109.980 ;
        RECT 91.840 109.800 92.010 109.980 ;
        RECT 92.320 109.800 92.490 109.980 ;
        RECT 92.800 109.800 92.970 109.980 ;
        RECT 93.280 109.800 93.450 109.980 ;
        RECT 93.760 109.800 93.930 109.980 ;
        RECT 94.240 109.800 94.410 109.980 ;
        RECT 94.720 109.800 94.890 109.980 ;
        RECT 95.200 109.800 95.370 109.980 ;
        RECT 95.680 109.800 95.850 109.980 ;
        RECT 96.160 109.800 96.330 109.980 ;
        RECT 96.640 109.800 96.810 109.980 ;
        RECT 97.120 109.800 97.290 109.980 ;
        RECT 97.600 109.800 97.770 109.980 ;
        RECT 98.080 109.800 98.250 109.980 ;
        RECT 98.560 109.800 98.730 109.980 ;
        RECT 99.040 109.800 99.210 109.980 ;
        RECT 99.520 109.800 99.690 109.980 ;
        RECT 100.000 109.800 100.170 109.980 ;
        RECT 100.480 109.800 100.650 109.980 ;
        RECT 100.960 109.800 101.130 109.980 ;
        RECT 101.440 109.800 101.610 109.980 ;
        RECT 101.920 109.800 102.090 109.980 ;
        RECT 102.400 109.800 102.570 109.980 ;
        RECT 102.880 109.800 103.050 109.980 ;
        RECT 103.360 109.800 103.530 109.980 ;
        RECT 103.840 109.800 104.010 109.980 ;
        RECT 104.320 109.800 104.490 109.980 ;
        RECT 104.800 109.800 104.970 109.980 ;
        RECT 105.280 109.800 105.450 109.980 ;
        RECT 105.760 109.800 105.930 109.980 ;
        RECT 106.240 109.800 106.410 109.980 ;
        RECT 106.720 109.800 106.890 109.980 ;
        RECT 107.200 109.800 107.370 109.980 ;
        RECT 107.680 109.800 107.850 109.980 ;
        RECT 108.160 109.800 108.330 109.980 ;
        RECT 108.640 109.800 108.810 109.980 ;
        RECT 109.120 109.800 109.290 109.980 ;
        RECT 109.600 109.800 109.770 109.980 ;
        RECT 110.080 109.800 110.250 109.980 ;
        RECT 110.560 109.800 110.730 109.980 ;
        RECT 111.040 109.800 111.210 109.980 ;
        RECT 111.520 109.800 111.690 109.980 ;
        RECT 112.000 109.800 112.170 109.980 ;
        RECT 112.480 109.800 112.650 109.980 ;
        RECT 112.960 109.800 113.130 109.980 ;
        RECT 113.440 109.800 113.610 109.980 ;
        RECT 113.920 109.800 114.090 109.980 ;
        RECT 114.400 109.800 114.570 109.980 ;
        RECT 114.880 109.800 115.050 109.980 ;
        RECT 115.360 109.800 115.530 109.980 ;
        RECT 115.840 109.800 116.010 109.980 ;
        RECT 116.320 109.800 116.490 109.980 ;
        RECT 116.800 109.800 116.970 109.980 ;
        RECT 117.280 109.800 117.450 109.980 ;
        RECT 117.760 109.800 117.930 109.980 ;
        RECT 118.240 109.800 118.410 109.980 ;
        RECT 118.720 109.800 118.890 109.980 ;
        RECT 119.200 109.800 119.370 109.980 ;
        RECT 119.680 109.800 119.850 109.980 ;
        RECT 120.160 109.800 120.330 109.980 ;
        RECT 120.640 109.800 120.810 109.980 ;
        RECT 121.120 109.800 121.290 109.980 ;
        RECT 121.600 109.800 121.770 109.980 ;
        RECT 122.080 109.800 122.250 109.980 ;
        RECT 122.560 109.800 122.730 109.980 ;
        RECT 123.040 109.800 123.210 109.980 ;
        RECT 123.520 109.800 123.690 109.980 ;
        RECT 124.000 109.800 124.170 109.980 ;
        RECT 124.480 109.800 124.650 109.980 ;
        RECT 124.960 109.800 125.130 109.980 ;
        RECT 125.440 109.800 125.610 109.980 ;
        RECT 125.920 109.800 126.090 109.980 ;
        RECT 126.400 109.800 126.570 109.980 ;
        RECT 126.880 109.800 127.050 109.980 ;
        RECT 127.360 109.800 127.530 109.980 ;
        RECT 127.840 109.800 128.010 109.980 ;
        RECT 128.320 109.800 128.490 109.980 ;
        RECT 128.800 109.800 128.970 109.980 ;
        RECT 129.280 109.800 129.450 109.980 ;
        RECT 129.760 109.800 129.930 109.980 ;
        RECT 130.240 109.800 130.410 109.980 ;
        RECT 130.720 109.800 130.890 109.980 ;
        RECT 131.200 109.800 131.370 109.980 ;
        RECT 131.680 109.800 131.850 109.980 ;
        RECT 132.160 109.800 132.330 109.980 ;
        RECT 132.640 109.800 132.810 109.980 ;
        RECT 133.120 109.800 133.290 109.980 ;
        RECT 133.600 109.800 133.770 109.980 ;
        RECT 134.080 109.800 134.250 109.980 ;
        RECT 134.560 109.800 134.730 109.980 ;
        RECT 135.040 109.800 135.210 109.980 ;
        RECT 135.520 109.800 135.690 109.980 ;
        RECT 136.000 109.800 136.170 109.980 ;
        RECT 136.480 109.800 136.650 109.980 ;
        RECT 136.960 109.800 137.130 109.980 ;
        RECT 137.440 109.800 137.610 109.980 ;
        RECT 137.920 109.800 138.090 109.980 ;
        RECT 138.400 109.800 138.570 109.980 ;
        RECT 138.880 109.800 139.050 109.980 ;
        RECT 139.360 109.800 139.530 109.980 ;
        RECT 139.840 109.800 140.010 109.980 ;
        RECT 140.320 109.800 140.490 109.980 ;
        RECT 140.800 109.800 140.970 109.980 ;
        RECT 141.280 109.800 141.450 109.980 ;
        RECT 141.760 109.800 141.930 109.980 ;
        RECT 6.510 109.330 6.680 109.500 ;
        RECT 6.950 109.330 7.120 109.500 ;
        RECT 7.360 109.330 7.530 109.500 ;
        RECT 7.790 109.330 7.960 109.500 ;
        RECT 8.230 109.330 8.400 109.500 ;
        RECT 8.640 109.330 8.810 109.500 ;
        RECT 10.350 109.330 10.520 109.500 ;
        RECT 10.790 109.330 10.960 109.500 ;
        RECT 11.200 109.330 11.370 109.500 ;
        RECT 11.630 109.330 11.800 109.500 ;
        RECT 12.070 109.330 12.240 109.500 ;
        RECT 12.480 109.330 12.650 109.500 ;
        RECT 14.190 109.330 14.360 109.500 ;
        RECT 14.630 109.330 14.800 109.500 ;
        RECT 15.040 109.330 15.210 109.500 ;
        RECT 15.470 109.330 15.640 109.500 ;
        RECT 15.910 109.330 16.080 109.500 ;
        RECT 16.320 109.330 16.490 109.500 ;
        RECT 18.030 109.330 18.200 109.500 ;
        RECT 18.470 109.330 18.640 109.500 ;
        RECT 18.880 109.330 19.050 109.500 ;
        RECT 19.310 109.330 19.480 109.500 ;
        RECT 19.750 109.330 19.920 109.500 ;
        RECT 20.160 109.330 20.330 109.500 ;
        RECT 21.340 109.320 21.510 109.490 ;
        RECT 21.780 109.320 21.950 109.490 ;
        RECT 22.220 109.320 22.390 109.490 ;
        RECT 22.630 109.320 22.800 109.490 ;
        RECT 25.240 109.320 25.410 109.490 ;
        RECT 25.600 109.320 25.770 109.490 ;
        RECT 25.960 109.320 26.130 109.490 ;
        RECT 27.100 109.320 27.270 109.490 ;
        RECT 27.540 109.320 27.710 109.490 ;
        RECT 27.980 109.320 28.150 109.490 ;
        RECT 28.390 109.320 28.560 109.490 ;
        RECT 29.390 109.320 29.560 109.490 ;
        RECT 29.750 109.320 29.920 109.490 ;
        RECT 30.110 109.320 30.280 109.490 ;
        RECT 31.030 109.320 31.200 109.490 ;
        RECT 31.390 109.320 31.560 109.490 ;
        RECT 35.990 109.320 36.160 109.490 ;
        RECT 36.350 109.320 36.520 109.490 ;
        RECT 36.710 109.320 36.880 109.490 ;
        RECT 39.960 109.320 40.130 109.490 ;
        RECT 40.320 109.320 40.490 109.490 ;
        RECT 40.680 109.320 40.850 109.490 ;
        RECT 42.570 109.320 42.740 109.490 ;
        RECT 42.930 109.320 43.100 109.490 ;
        RECT 43.290 109.320 43.460 109.490 ;
        RECT 44.380 109.320 44.550 109.490 ;
        RECT 44.820 109.320 44.990 109.490 ;
        RECT 45.260 109.320 45.430 109.490 ;
        RECT 45.670 109.320 45.840 109.490 ;
        RECT 46.200 109.320 46.370 109.490 ;
        RECT 46.560 109.320 46.730 109.490 ;
        RECT 47.740 109.320 47.910 109.490 ;
        RECT 48.180 109.320 48.350 109.490 ;
        RECT 48.620 109.320 48.790 109.490 ;
        RECT 49.030 109.320 49.200 109.490 ;
        RECT 50.030 109.320 50.200 109.490 ;
        RECT 50.390 109.320 50.560 109.490 ;
        RECT 50.750 109.320 50.920 109.490 ;
        RECT 51.670 109.320 51.840 109.490 ;
        RECT 52.030 109.320 52.200 109.490 ;
        RECT 56.630 109.320 56.800 109.490 ;
        RECT 56.990 109.320 57.160 109.490 ;
        RECT 57.350 109.320 57.520 109.490 ;
        RECT 60.600 109.320 60.770 109.490 ;
        RECT 60.960 109.320 61.130 109.490 ;
        RECT 61.320 109.320 61.490 109.490 ;
        RECT 63.210 109.320 63.380 109.490 ;
        RECT 63.570 109.320 63.740 109.490 ;
        RECT 63.930 109.320 64.100 109.490 ;
        RECT 65.020 109.320 65.190 109.490 ;
        RECT 65.460 109.320 65.630 109.490 ;
        RECT 65.900 109.320 66.070 109.490 ;
        RECT 66.310 109.320 66.480 109.490 ;
        RECT 66.840 109.320 67.010 109.490 ;
        RECT 67.200 109.320 67.370 109.490 ;
        RECT 67.560 109.320 67.730 109.490 ;
        RECT 68.400 109.320 68.570 109.490 ;
        RECT 68.760 109.320 68.930 109.490 ;
        RECT 69.120 109.320 69.290 109.490 ;
        RECT 69.960 109.320 70.130 109.490 ;
        RECT 70.320 109.320 70.490 109.490 ;
        RECT 70.680 109.320 70.850 109.490 ;
        RECT 71.740 109.320 71.910 109.490 ;
        RECT 72.180 109.320 72.350 109.490 ;
        RECT 72.620 109.320 72.790 109.490 ;
        RECT 73.030 109.320 73.200 109.490 ;
        RECT 74.030 109.320 74.200 109.490 ;
        RECT 74.390 109.320 74.560 109.490 ;
        RECT 74.750 109.320 74.920 109.490 ;
        RECT 75.670 109.320 75.840 109.490 ;
        RECT 76.030 109.320 76.200 109.490 ;
        RECT 76.540 109.320 76.710 109.490 ;
        RECT 76.980 109.320 77.150 109.490 ;
        RECT 77.420 109.320 77.590 109.490 ;
        RECT 77.830 109.320 78.000 109.490 ;
        RECT 80.440 109.320 80.610 109.490 ;
        RECT 80.800 109.320 80.970 109.490 ;
        RECT 81.160 109.320 81.330 109.490 ;
        RECT 82.300 109.320 82.470 109.490 ;
        RECT 82.740 109.320 82.910 109.490 ;
        RECT 83.180 109.320 83.350 109.490 ;
        RECT 83.590 109.320 83.760 109.490 ;
        RECT 84.560 109.320 84.730 109.490 ;
        RECT 84.920 109.320 85.090 109.490 ;
        RECT 85.280 109.320 85.450 109.490 ;
        RECT 87.920 109.320 88.090 109.490 ;
        RECT 88.280 109.320 88.450 109.490 ;
        RECT 88.640 109.320 88.810 109.490 ;
        RECT 89.000 109.320 89.170 109.490 ;
        RECT 89.500 109.320 89.670 109.490 ;
        RECT 89.940 109.320 90.110 109.490 ;
        RECT 90.380 109.320 90.550 109.490 ;
        RECT 90.790 109.320 90.960 109.490 ;
        RECT 92.280 109.320 92.450 109.490 ;
        RECT 92.640 109.320 92.810 109.490 ;
        RECT 93.000 109.320 93.170 109.490 ;
        RECT 93.840 109.320 94.010 109.490 ;
        RECT 94.200 109.320 94.370 109.490 ;
        RECT 94.560 109.320 94.730 109.490 ;
        RECT 95.400 109.320 95.570 109.490 ;
        RECT 95.760 109.320 95.930 109.490 ;
        RECT 96.120 109.320 96.290 109.490 ;
        RECT 97.180 109.320 97.350 109.490 ;
        RECT 97.620 109.320 97.790 109.490 ;
        RECT 98.060 109.320 98.230 109.490 ;
        RECT 98.470 109.320 98.640 109.490 ;
        RECT 99.000 109.320 99.170 109.490 ;
        RECT 99.360 109.320 99.530 109.490 ;
        RECT 99.720 109.320 99.890 109.490 ;
        RECT 100.560 109.320 100.730 109.490 ;
        RECT 100.920 109.320 101.090 109.490 ;
        RECT 101.280 109.320 101.450 109.490 ;
        RECT 102.120 109.320 102.290 109.490 ;
        RECT 102.480 109.320 102.650 109.490 ;
        RECT 102.840 109.320 103.010 109.490 ;
        RECT 103.900 109.320 104.070 109.490 ;
        RECT 104.340 109.320 104.510 109.490 ;
        RECT 104.780 109.320 104.950 109.490 ;
        RECT 105.190 109.320 105.360 109.490 ;
        RECT 105.720 109.320 105.890 109.490 ;
        RECT 106.080 109.320 106.250 109.490 ;
        RECT 106.440 109.320 106.610 109.490 ;
        RECT 107.280 109.320 107.450 109.490 ;
        RECT 107.640 109.320 107.810 109.490 ;
        RECT 108.000 109.320 108.170 109.490 ;
        RECT 108.840 109.320 109.010 109.490 ;
        RECT 109.200 109.320 109.370 109.490 ;
        RECT 109.560 109.320 109.730 109.490 ;
        RECT 110.620 109.320 110.790 109.490 ;
        RECT 111.060 109.320 111.230 109.490 ;
        RECT 111.500 109.320 111.670 109.490 ;
        RECT 111.910 109.320 112.080 109.490 ;
        RECT 112.870 109.320 113.040 109.490 ;
        RECT 113.230 109.320 113.400 109.490 ;
        RECT 113.590 109.320 113.760 109.490 ;
        RECT 113.950 109.320 114.120 109.490 ;
        RECT 114.940 109.320 115.110 109.490 ;
        RECT 115.380 109.320 115.550 109.490 ;
        RECT 115.820 109.320 115.990 109.490 ;
        RECT 116.230 109.320 116.400 109.490 ;
        RECT 117.670 109.320 117.840 109.490 ;
        RECT 118.030 109.320 118.200 109.490 ;
        RECT 118.390 109.320 118.560 109.490 ;
        RECT 118.750 109.320 118.920 109.490 ;
        RECT 119.740 109.320 119.910 109.490 ;
        RECT 120.180 109.320 120.350 109.490 ;
        RECT 120.620 109.320 120.790 109.490 ;
        RECT 121.030 109.320 121.200 109.490 ;
        RECT 121.560 109.320 121.730 109.490 ;
        RECT 121.920 109.320 122.090 109.490 ;
        RECT 122.280 109.320 122.450 109.490 ;
        RECT 123.120 109.320 123.290 109.490 ;
        RECT 123.480 109.320 123.650 109.490 ;
        RECT 123.840 109.320 124.010 109.490 ;
        RECT 124.680 109.320 124.850 109.490 ;
        RECT 125.040 109.320 125.210 109.490 ;
        RECT 125.400 109.320 125.570 109.490 ;
        RECT 126.990 109.330 127.160 109.500 ;
        RECT 127.430 109.330 127.600 109.500 ;
        RECT 127.840 109.330 128.010 109.500 ;
        RECT 128.270 109.330 128.440 109.500 ;
        RECT 128.710 109.330 128.880 109.500 ;
        RECT 129.120 109.330 129.290 109.500 ;
        RECT 130.830 109.330 131.000 109.500 ;
        RECT 131.270 109.330 131.440 109.500 ;
        RECT 131.680 109.330 131.850 109.500 ;
        RECT 132.110 109.330 132.280 109.500 ;
        RECT 132.550 109.330 132.720 109.500 ;
        RECT 132.960 109.330 133.130 109.500 ;
        RECT 134.670 109.330 134.840 109.500 ;
        RECT 135.110 109.330 135.280 109.500 ;
        RECT 135.520 109.330 135.690 109.500 ;
        RECT 135.950 109.330 136.120 109.500 ;
        RECT 136.390 109.330 136.560 109.500 ;
        RECT 136.800 109.330 136.970 109.500 ;
        RECT 138.510 109.330 138.680 109.500 ;
        RECT 138.950 109.330 139.120 109.500 ;
        RECT 139.360 109.330 139.530 109.500 ;
        RECT 139.790 109.330 139.960 109.500 ;
        RECT 140.230 109.330 140.400 109.500 ;
        RECT 140.640 109.330 140.810 109.500 ;
        RECT 5.920 101.660 6.090 101.840 ;
        RECT 6.400 101.660 6.570 101.840 ;
        RECT 6.880 101.660 7.050 101.840 ;
        RECT 7.360 101.660 7.530 101.840 ;
        RECT 7.840 101.660 8.010 101.840 ;
        RECT 8.320 101.660 8.490 101.840 ;
        RECT 8.800 101.660 8.970 101.840 ;
        RECT 9.280 101.660 9.450 101.840 ;
        RECT 9.760 101.660 9.930 101.840 ;
        RECT 10.240 101.660 10.410 101.840 ;
        RECT 10.720 101.660 10.890 101.840 ;
        RECT 11.200 101.660 11.370 101.840 ;
        RECT 11.680 101.660 11.850 101.840 ;
        RECT 12.160 101.660 12.330 101.840 ;
        RECT 12.640 101.660 12.810 101.840 ;
        RECT 13.120 101.660 13.290 101.840 ;
        RECT 13.600 101.660 13.770 101.840 ;
        RECT 14.080 101.660 14.250 101.840 ;
        RECT 14.560 101.660 14.730 101.840 ;
        RECT 15.040 101.660 15.210 101.840 ;
        RECT 15.520 101.660 15.690 101.840 ;
        RECT 16.000 101.660 16.170 101.840 ;
        RECT 16.480 101.660 16.650 101.840 ;
        RECT 16.960 101.660 17.130 101.840 ;
        RECT 17.440 101.660 17.610 101.840 ;
        RECT 17.920 101.660 18.090 101.840 ;
        RECT 18.400 101.660 18.570 101.840 ;
        RECT 18.880 101.660 19.050 101.840 ;
        RECT 19.360 101.660 19.530 101.840 ;
        RECT 19.840 101.660 20.010 101.840 ;
        RECT 20.320 101.660 20.490 101.840 ;
        RECT 20.800 101.660 20.970 101.840 ;
        RECT 21.280 101.660 21.450 101.840 ;
        RECT 21.760 101.660 21.930 101.840 ;
        RECT 22.240 101.660 22.410 101.840 ;
        RECT 22.720 101.660 22.890 101.840 ;
        RECT 23.200 101.660 23.370 101.840 ;
        RECT 23.680 101.660 23.850 101.840 ;
        RECT 24.160 101.660 24.330 101.840 ;
        RECT 24.640 101.660 24.810 101.840 ;
        RECT 25.120 101.660 25.290 101.840 ;
        RECT 25.600 101.660 25.770 101.840 ;
        RECT 26.080 101.660 26.250 101.840 ;
        RECT 26.560 101.660 26.730 101.840 ;
        RECT 27.040 101.660 27.210 101.840 ;
        RECT 27.520 101.660 27.690 101.840 ;
        RECT 28.000 101.660 28.170 101.840 ;
        RECT 28.480 101.660 28.650 101.840 ;
        RECT 28.960 101.660 29.130 101.840 ;
        RECT 29.440 101.660 29.610 101.840 ;
        RECT 29.920 101.660 30.090 101.840 ;
        RECT 30.400 101.660 30.570 101.840 ;
        RECT 30.880 101.660 31.050 101.840 ;
        RECT 31.360 101.660 31.530 101.840 ;
        RECT 31.840 101.660 32.010 101.840 ;
        RECT 32.320 101.660 32.490 101.840 ;
        RECT 32.800 101.660 32.970 101.840 ;
        RECT 33.280 101.660 33.450 101.840 ;
        RECT 33.760 101.660 33.930 101.840 ;
        RECT 34.240 101.660 34.410 101.840 ;
        RECT 34.720 101.660 34.890 101.840 ;
        RECT 35.200 101.660 35.370 101.840 ;
        RECT 35.680 101.660 35.850 101.840 ;
        RECT 36.160 101.660 36.330 101.840 ;
        RECT 36.640 101.660 36.810 101.840 ;
        RECT 37.120 101.660 37.290 101.840 ;
        RECT 37.600 101.660 37.770 101.840 ;
        RECT 38.080 101.660 38.250 101.840 ;
        RECT 38.560 101.660 38.730 101.840 ;
        RECT 39.040 101.660 39.210 101.840 ;
        RECT 39.520 101.660 39.690 101.840 ;
        RECT 40.000 101.660 40.170 101.840 ;
      LAYER li1 ;
        RECT 40.320 101.660 40.800 101.840 ;
      LAYER li1 ;
        RECT 40.960 101.660 41.130 101.840 ;
        RECT 41.440 101.660 41.610 101.840 ;
        RECT 41.920 101.660 42.090 101.840 ;
        RECT 42.400 101.660 42.570 101.840 ;
        RECT 42.880 101.660 43.050 101.840 ;
        RECT 43.360 101.660 43.530 101.840 ;
        RECT 43.840 101.660 44.010 101.840 ;
        RECT 44.320 101.660 44.490 101.840 ;
        RECT 44.800 101.660 44.970 101.840 ;
        RECT 45.280 101.660 45.450 101.840 ;
        RECT 45.760 101.660 45.930 101.840 ;
        RECT 46.240 101.660 46.410 101.840 ;
        RECT 46.720 101.660 46.890 101.840 ;
        RECT 47.200 101.660 47.370 101.840 ;
        RECT 47.680 101.660 47.850 101.840 ;
        RECT 48.160 101.660 48.330 101.840 ;
        RECT 48.640 101.660 48.810 101.840 ;
        RECT 49.120 101.660 49.290 101.840 ;
        RECT 49.600 101.660 49.770 101.840 ;
        RECT 50.080 101.660 50.250 101.840 ;
        RECT 50.560 101.660 50.730 101.840 ;
        RECT 51.040 101.660 51.210 101.840 ;
        RECT 51.520 101.660 51.690 101.840 ;
        RECT 52.000 101.660 52.170 101.840 ;
        RECT 52.480 101.660 52.650 101.840 ;
        RECT 52.960 101.660 53.130 101.840 ;
        RECT 53.440 101.660 53.610 101.840 ;
        RECT 53.920 101.660 54.090 101.840 ;
        RECT 54.400 101.660 54.570 101.840 ;
        RECT 54.880 101.660 55.050 101.840 ;
        RECT 55.360 101.660 55.530 101.840 ;
        RECT 55.840 101.660 56.010 101.840 ;
        RECT 56.320 101.660 56.490 101.840 ;
        RECT 56.800 101.660 56.970 101.840 ;
        RECT 57.280 101.660 57.450 101.840 ;
        RECT 57.760 101.660 57.930 101.840 ;
        RECT 58.240 101.660 58.410 101.840 ;
        RECT 58.720 101.660 58.890 101.840 ;
        RECT 59.200 101.660 59.370 101.840 ;
        RECT 59.680 101.660 59.850 101.840 ;
        RECT 60.160 101.660 60.330 101.840 ;
        RECT 60.640 101.660 60.810 101.840 ;
      LAYER li1 ;
        RECT 60.960 101.660 61.440 101.840 ;
      LAYER li1 ;
        RECT 61.600 101.660 61.770 101.840 ;
        RECT 62.080 101.660 62.250 101.840 ;
        RECT 62.560 101.660 62.730 101.840 ;
        RECT 63.040 101.660 63.210 101.840 ;
        RECT 63.520 101.660 63.690 101.840 ;
        RECT 64.000 101.660 64.170 101.840 ;
        RECT 64.480 101.660 64.650 101.840 ;
        RECT 64.960 101.660 65.130 101.840 ;
        RECT 65.440 101.660 65.610 101.840 ;
        RECT 65.920 101.660 66.090 101.840 ;
        RECT 66.400 101.660 66.570 101.840 ;
        RECT 66.880 101.660 67.050 101.840 ;
        RECT 67.360 101.660 67.530 101.840 ;
        RECT 67.840 101.660 68.010 101.840 ;
        RECT 68.320 101.660 68.490 101.840 ;
        RECT 68.800 101.660 68.970 101.840 ;
        RECT 69.280 101.660 69.450 101.840 ;
        RECT 69.760 101.660 69.930 101.840 ;
        RECT 70.240 101.660 70.410 101.840 ;
        RECT 70.720 101.660 70.890 101.840 ;
        RECT 71.200 101.660 71.370 101.840 ;
        RECT 71.680 101.660 71.850 101.840 ;
        RECT 72.160 101.660 72.330 101.840 ;
        RECT 72.640 101.660 72.810 101.840 ;
        RECT 73.120 101.660 73.290 101.840 ;
        RECT 73.600 101.660 73.770 101.840 ;
        RECT 74.080 101.660 74.250 101.840 ;
        RECT 74.560 101.660 74.730 101.840 ;
        RECT 75.040 101.660 75.210 101.840 ;
        RECT 75.520 101.660 75.690 101.840 ;
        RECT 76.000 101.660 76.170 101.840 ;
        RECT 76.480 101.660 76.650 101.840 ;
        RECT 76.960 101.660 77.130 101.840 ;
        RECT 77.440 101.660 77.610 101.840 ;
        RECT 77.920 101.660 78.090 101.840 ;
        RECT 78.400 101.660 78.570 101.840 ;
        RECT 78.880 101.660 79.050 101.840 ;
        RECT 79.360 101.660 79.530 101.840 ;
        RECT 79.840 101.660 80.010 101.840 ;
        RECT 80.320 101.660 80.490 101.840 ;
        RECT 80.800 101.660 80.970 101.840 ;
        RECT 81.280 101.660 81.450 101.840 ;
        RECT 81.760 101.660 81.930 101.840 ;
        RECT 82.240 101.660 82.410 101.840 ;
        RECT 82.720 101.660 82.890 101.840 ;
        RECT 83.200 101.660 83.370 101.840 ;
        RECT 83.680 101.660 83.850 101.840 ;
        RECT 84.160 101.660 84.330 101.840 ;
        RECT 84.640 101.660 84.810 101.840 ;
        RECT 85.120 101.660 85.290 101.840 ;
        RECT 85.600 101.660 85.770 101.840 ;
        RECT 86.080 101.660 86.250 101.840 ;
        RECT 86.560 101.660 86.730 101.840 ;
        RECT 87.040 101.660 87.210 101.840 ;
        RECT 87.520 101.660 87.690 101.840 ;
        RECT 88.000 101.660 88.170 101.840 ;
        RECT 88.480 101.660 88.650 101.840 ;
        RECT 88.960 101.660 89.130 101.840 ;
        RECT 89.440 101.660 89.610 101.840 ;
        RECT 89.920 101.660 90.090 101.840 ;
        RECT 90.400 101.660 90.570 101.840 ;
        RECT 90.880 101.660 91.050 101.840 ;
        RECT 91.360 101.660 91.530 101.840 ;
        RECT 91.840 101.660 92.010 101.840 ;
        RECT 92.320 101.660 92.490 101.840 ;
        RECT 92.800 101.660 92.970 101.840 ;
        RECT 93.280 101.660 93.450 101.840 ;
        RECT 93.760 101.660 93.930 101.840 ;
        RECT 94.240 101.660 94.410 101.840 ;
        RECT 94.720 101.660 94.890 101.840 ;
        RECT 95.200 101.660 95.370 101.840 ;
        RECT 95.680 101.660 95.850 101.840 ;
        RECT 96.160 101.660 96.330 101.840 ;
        RECT 96.640 101.660 96.810 101.840 ;
        RECT 97.120 101.660 97.290 101.840 ;
        RECT 97.600 101.660 97.770 101.840 ;
        RECT 98.080 101.660 98.250 101.840 ;
        RECT 98.560 101.660 98.730 101.840 ;
        RECT 99.040 101.660 99.210 101.840 ;
        RECT 99.520 101.660 99.690 101.840 ;
        RECT 100.000 101.660 100.170 101.840 ;
        RECT 100.480 101.660 100.650 101.840 ;
        RECT 100.960 101.660 101.130 101.840 ;
        RECT 101.440 101.660 101.610 101.840 ;
        RECT 101.920 101.660 102.090 101.840 ;
        RECT 102.400 101.660 102.570 101.840 ;
        RECT 102.880 101.660 103.050 101.840 ;
        RECT 103.360 101.660 103.530 101.840 ;
        RECT 103.840 101.660 104.010 101.840 ;
        RECT 104.320 101.660 104.490 101.840 ;
        RECT 104.800 101.660 104.970 101.840 ;
        RECT 105.280 101.660 105.450 101.840 ;
        RECT 105.760 101.660 105.930 101.840 ;
        RECT 106.240 101.660 106.410 101.840 ;
        RECT 106.720 101.660 106.890 101.840 ;
        RECT 107.200 101.660 107.370 101.840 ;
        RECT 107.680 101.660 107.850 101.840 ;
        RECT 108.160 101.660 108.330 101.840 ;
        RECT 108.640 101.660 108.810 101.840 ;
        RECT 109.120 101.660 109.290 101.840 ;
        RECT 109.600 101.660 109.770 101.840 ;
        RECT 110.080 101.660 110.250 101.840 ;
        RECT 110.560 101.660 110.730 101.840 ;
        RECT 111.040 101.660 111.210 101.840 ;
        RECT 111.520 101.660 111.690 101.840 ;
        RECT 112.000 101.660 112.170 101.840 ;
        RECT 112.480 101.660 112.650 101.840 ;
        RECT 112.960 101.660 113.130 101.840 ;
        RECT 113.440 101.660 113.610 101.840 ;
        RECT 113.920 101.660 114.090 101.840 ;
        RECT 114.400 101.660 114.570 101.840 ;
        RECT 114.880 101.660 115.050 101.840 ;
        RECT 115.360 101.660 115.530 101.840 ;
        RECT 115.840 101.660 116.010 101.840 ;
        RECT 116.320 101.660 116.490 101.840 ;
        RECT 116.800 101.660 116.970 101.840 ;
        RECT 117.280 101.660 117.450 101.840 ;
        RECT 117.760 101.660 117.930 101.840 ;
        RECT 118.240 101.660 118.410 101.840 ;
        RECT 118.720 101.660 118.890 101.840 ;
        RECT 119.200 101.660 119.370 101.840 ;
        RECT 119.680 101.660 119.850 101.840 ;
        RECT 120.160 101.660 120.330 101.840 ;
        RECT 120.640 101.660 120.810 101.840 ;
      LAYER li1 ;
        RECT 120.960 101.660 121.440 101.840 ;
      LAYER li1 ;
        RECT 121.600 101.660 121.770 101.840 ;
        RECT 122.080 101.660 122.250 101.840 ;
        RECT 122.560 101.660 122.730 101.840 ;
        RECT 123.040 101.660 123.210 101.840 ;
        RECT 123.520 101.660 123.690 101.840 ;
        RECT 124.000 101.660 124.170 101.840 ;
        RECT 124.480 101.660 124.650 101.840 ;
        RECT 124.960 101.660 125.130 101.840 ;
        RECT 125.440 101.660 125.610 101.840 ;
        RECT 125.920 101.660 126.090 101.840 ;
        RECT 126.400 101.660 126.570 101.840 ;
        RECT 126.880 101.660 127.050 101.840 ;
        RECT 127.360 101.660 127.530 101.840 ;
        RECT 127.840 101.660 128.010 101.840 ;
        RECT 128.320 101.660 128.490 101.840 ;
        RECT 128.800 101.660 128.970 101.840 ;
        RECT 129.280 101.660 129.450 101.840 ;
        RECT 129.760 101.660 129.930 101.840 ;
        RECT 130.240 101.660 130.410 101.840 ;
        RECT 130.720 101.660 130.890 101.840 ;
        RECT 131.200 101.660 131.370 101.840 ;
        RECT 131.680 101.660 131.850 101.840 ;
        RECT 132.160 101.660 132.330 101.840 ;
        RECT 132.640 101.660 132.810 101.840 ;
        RECT 133.120 101.660 133.290 101.840 ;
        RECT 133.600 101.660 133.770 101.840 ;
        RECT 134.080 101.660 134.250 101.840 ;
        RECT 134.560 101.660 134.730 101.840 ;
        RECT 135.040 101.660 135.210 101.840 ;
        RECT 135.520 101.660 135.690 101.840 ;
        RECT 136.000 101.660 136.170 101.840 ;
        RECT 136.480 101.660 136.650 101.840 ;
        RECT 136.960 101.660 137.130 101.840 ;
        RECT 137.440 101.660 137.610 101.840 ;
        RECT 137.920 101.660 138.090 101.840 ;
        RECT 138.400 101.660 138.570 101.840 ;
        RECT 138.880 101.660 139.050 101.840 ;
        RECT 139.360 101.660 139.530 101.840 ;
        RECT 139.840 101.660 140.010 101.840 ;
        RECT 140.320 101.660 140.490 101.840 ;
        RECT 140.800 101.660 140.970 101.840 ;
        RECT 141.280 101.660 141.450 101.840 ;
        RECT 141.760 101.660 141.930 101.840 ;
        RECT 6.510 101.190 6.680 101.360 ;
        RECT 6.950 101.190 7.120 101.360 ;
        RECT 7.360 101.190 7.530 101.360 ;
        RECT 7.790 101.190 7.960 101.360 ;
        RECT 8.230 101.190 8.400 101.360 ;
        RECT 8.640 101.190 8.810 101.360 ;
        RECT 10.350 101.190 10.520 101.360 ;
        RECT 10.790 101.190 10.960 101.360 ;
        RECT 11.200 101.190 11.370 101.360 ;
        RECT 11.630 101.190 11.800 101.360 ;
        RECT 12.070 101.190 12.240 101.360 ;
        RECT 12.480 101.190 12.650 101.360 ;
        RECT 13.660 101.180 13.830 101.350 ;
        RECT 14.100 101.180 14.270 101.350 ;
        RECT 14.540 101.180 14.710 101.350 ;
        RECT 14.950 101.180 15.120 101.350 ;
        RECT 16.870 101.180 17.040 101.350 ;
        RECT 17.230 101.180 17.400 101.350 ;
        RECT 17.590 101.180 17.760 101.350 ;
        RECT 17.950 101.180 18.120 101.350 ;
        RECT 18.940 101.180 19.110 101.350 ;
        RECT 19.380 101.180 19.550 101.350 ;
        RECT 19.820 101.180 19.990 101.350 ;
        RECT 20.230 101.180 20.400 101.350 ;
        RECT 22.200 101.180 22.370 101.350 ;
        RECT 22.560 101.180 22.730 101.350 ;
        RECT 24.270 101.190 24.440 101.360 ;
        RECT 24.710 101.190 24.880 101.360 ;
        RECT 25.120 101.190 25.290 101.360 ;
        RECT 25.550 101.190 25.720 101.360 ;
        RECT 25.990 101.190 26.160 101.360 ;
        RECT 26.400 101.190 26.570 101.360 ;
        RECT 28.920 101.180 29.090 101.350 ;
        RECT 29.280 101.180 29.450 101.350 ;
        RECT 30.460 101.180 30.630 101.350 ;
        RECT 30.900 101.180 31.070 101.350 ;
        RECT 31.340 101.180 31.510 101.350 ;
        RECT 31.750 101.180 31.920 101.350 ;
        RECT 32.710 101.180 32.880 101.350 ;
        RECT 33.070 101.180 33.240 101.350 ;
        RECT 33.430 101.180 33.600 101.350 ;
        RECT 33.790 101.180 33.960 101.350 ;
        RECT 34.780 101.180 34.950 101.350 ;
        RECT 35.220 101.180 35.390 101.350 ;
        RECT 35.660 101.180 35.830 101.350 ;
        RECT 36.070 101.180 36.240 101.350 ;
        RECT 37.030 101.180 37.200 101.350 ;
        RECT 37.390 101.180 37.560 101.350 ;
        RECT 37.750 101.180 37.920 101.350 ;
        RECT 38.110 101.180 38.280 101.350 ;
        RECT 39.100 101.180 39.270 101.350 ;
        RECT 39.540 101.180 39.710 101.350 ;
        RECT 39.980 101.180 40.150 101.350 ;
        RECT 40.390 101.180 40.560 101.350 ;
        RECT 40.920 101.180 41.090 101.350 ;
        RECT 41.280 101.180 41.450 101.350 ;
        RECT 41.640 101.180 41.810 101.350 ;
        RECT 42.480 101.180 42.650 101.350 ;
        RECT 42.840 101.180 43.010 101.350 ;
        RECT 43.200 101.180 43.370 101.350 ;
        RECT 44.040 101.180 44.210 101.350 ;
        RECT 44.400 101.180 44.570 101.350 ;
        RECT 44.760 101.180 44.930 101.350 ;
        RECT 45.820 101.180 45.990 101.350 ;
        RECT 46.260 101.180 46.430 101.350 ;
        RECT 46.700 101.180 46.870 101.350 ;
        RECT 47.110 101.180 47.280 101.350 ;
        RECT 47.640 101.180 47.810 101.350 ;
        RECT 48.000 101.180 48.170 101.350 ;
        RECT 48.360 101.180 48.530 101.350 ;
        RECT 49.200 101.180 49.370 101.350 ;
        RECT 49.560 101.180 49.730 101.350 ;
        RECT 49.920 101.180 50.090 101.350 ;
        RECT 50.760 101.180 50.930 101.350 ;
        RECT 51.120 101.180 51.290 101.350 ;
        RECT 51.480 101.180 51.650 101.350 ;
        RECT 52.540 101.180 52.710 101.350 ;
        RECT 52.980 101.180 53.150 101.350 ;
        RECT 53.420 101.180 53.590 101.350 ;
        RECT 53.830 101.180 54.000 101.350 ;
        RECT 54.360 101.180 54.530 101.350 ;
        RECT 54.720 101.180 54.890 101.350 ;
        RECT 55.080 101.180 55.250 101.350 ;
        RECT 55.920 101.180 56.090 101.350 ;
        RECT 56.280 101.180 56.450 101.350 ;
        RECT 56.640 101.180 56.810 101.350 ;
        RECT 57.480 101.180 57.650 101.350 ;
        RECT 57.840 101.180 58.010 101.350 ;
        RECT 58.200 101.180 58.370 101.350 ;
        RECT 59.260 101.180 59.430 101.350 ;
        RECT 59.700 101.180 59.870 101.350 ;
        RECT 60.140 101.180 60.310 101.350 ;
        RECT 60.550 101.180 60.720 101.350 ;
        RECT 63.160 101.180 63.330 101.350 ;
        RECT 63.520 101.180 63.690 101.350 ;
        RECT 63.880 101.180 64.050 101.350 ;
        RECT 65.020 101.180 65.190 101.350 ;
        RECT 65.460 101.180 65.630 101.350 ;
        RECT 65.900 101.180 66.070 101.350 ;
        RECT 66.310 101.180 66.480 101.350 ;
        RECT 67.270 101.180 67.440 101.350 ;
        RECT 67.630 101.180 67.800 101.350 ;
        RECT 67.990 101.180 68.160 101.350 ;
        RECT 68.350 101.180 68.520 101.350 ;
        RECT 69.340 101.180 69.510 101.350 ;
        RECT 69.780 101.180 69.950 101.350 ;
        RECT 70.220 101.180 70.390 101.350 ;
        RECT 70.630 101.180 70.800 101.350 ;
        RECT 72.600 101.180 72.770 101.350 ;
        RECT 72.960 101.180 73.130 101.350 ;
        RECT 73.870 101.180 74.040 101.350 ;
        RECT 74.230 101.180 74.400 101.350 ;
        RECT 74.590 101.180 74.760 101.350 ;
        RECT 76.060 101.180 76.230 101.350 ;
        RECT 76.500 101.180 76.670 101.350 ;
        RECT 76.940 101.180 77.110 101.350 ;
        RECT 77.350 101.180 77.520 101.350 ;
        RECT 77.880 101.180 78.050 101.350 ;
        RECT 78.240 101.180 78.410 101.350 ;
        RECT 78.600 101.180 78.770 101.350 ;
        RECT 79.440 101.180 79.610 101.350 ;
        RECT 79.800 101.180 79.970 101.350 ;
        RECT 80.160 101.180 80.330 101.350 ;
        RECT 81.000 101.180 81.170 101.350 ;
        RECT 81.360 101.180 81.530 101.350 ;
        RECT 81.720 101.180 81.890 101.350 ;
        RECT 82.780 101.180 82.950 101.350 ;
        RECT 83.220 101.180 83.390 101.350 ;
        RECT 83.660 101.180 83.830 101.350 ;
        RECT 84.070 101.180 84.240 101.350 ;
        RECT 84.600 101.180 84.770 101.350 ;
        RECT 84.960 101.180 85.130 101.350 ;
        RECT 85.320 101.180 85.490 101.350 ;
        RECT 86.160 101.180 86.330 101.350 ;
        RECT 86.520 101.180 86.690 101.350 ;
        RECT 86.880 101.180 87.050 101.350 ;
        RECT 87.720 101.180 87.890 101.350 ;
        RECT 88.080 101.180 88.250 101.350 ;
        RECT 88.440 101.180 88.610 101.350 ;
        RECT 90.030 101.190 90.200 101.360 ;
        RECT 90.470 101.190 90.640 101.360 ;
        RECT 90.880 101.190 91.050 101.360 ;
        RECT 91.310 101.190 91.480 101.360 ;
        RECT 91.750 101.190 91.920 101.360 ;
        RECT 92.160 101.190 92.330 101.360 ;
        RECT 93.240 101.180 93.410 101.350 ;
        RECT 93.600 101.180 93.770 101.350 ;
        RECT 93.960 101.180 94.130 101.350 ;
        RECT 94.800 101.180 94.970 101.350 ;
        RECT 95.160 101.180 95.330 101.350 ;
        RECT 95.520 101.180 95.690 101.350 ;
        RECT 96.360 101.180 96.530 101.350 ;
        RECT 96.720 101.180 96.890 101.350 ;
        RECT 97.080 101.180 97.250 101.350 ;
        RECT 98.140 101.180 98.310 101.350 ;
        RECT 98.580 101.180 98.750 101.350 ;
        RECT 99.020 101.180 99.190 101.350 ;
        RECT 99.430 101.180 99.600 101.350 ;
        RECT 100.400 101.180 100.570 101.350 ;
        RECT 100.760 101.180 100.930 101.350 ;
        RECT 101.120 101.180 101.290 101.350 ;
        RECT 103.760 101.180 103.930 101.350 ;
        RECT 104.120 101.180 104.290 101.350 ;
        RECT 104.480 101.180 104.650 101.350 ;
        RECT 104.840 101.180 105.010 101.350 ;
        RECT 105.340 101.180 105.510 101.350 ;
        RECT 105.780 101.180 105.950 101.350 ;
        RECT 106.220 101.180 106.390 101.350 ;
        RECT 106.630 101.180 106.800 101.350 ;
        RECT 107.590 101.180 107.760 101.350 ;
        RECT 107.950 101.180 108.120 101.350 ;
        RECT 108.310 101.180 108.480 101.350 ;
        RECT 108.670 101.180 108.840 101.350 ;
        RECT 109.660 101.180 109.830 101.350 ;
        RECT 110.100 101.180 110.270 101.350 ;
        RECT 110.540 101.180 110.710 101.350 ;
        RECT 110.950 101.180 111.120 101.350 ;
        RECT 111.960 101.180 112.130 101.350 ;
        RECT 112.320 101.180 112.490 101.350 ;
        RECT 113.830 101.180 114.000 101.350 ;
        RECT 114.190 101.180 114.360 101.350 ;
        RECT 116.250 101.180 116.420 101.350 ;
        RECT 116.610 101.180 116.780 101.350 ;
        RECT 116.970 101.180 117.140 101.350 ;
        RECT 118.190 101.180 118.360 101.350 ;
        RECT 118.550 101.180 118.720 101.350 ;
        RECT 118.910 101.180 119.080 101.350 ;
        RECT 122.730 101.180 122.900 101.350 ;
        RECT 123.090 101.180 123.260 101.350 ;
        RECT 124.650 101.180 124.820 101.350 ;
        RECT 125.010 101.180 125.180 101.350 ;
        RECT 125.370 101.180 125.540 101.350 ;
        RECT 126.460 101.180 126.630 101.350 ;
        RECT 126.900 101.180 127.070 101.350 ;
        RECT 127.340 101.180 127.510 101.350 ;
        RECT 127.750 101.180 127.920 101.350 ;
        RECT 128.280 101.180 128.450 101.350 ;
        RECT 128.640 101.180 128.810 101.350 ;
        RECT 129.000 101.180 129.170 101.350 ;
        RECT 129.840 101.180 130.010 101.350 ;
        RECT 130.200 101.180 130.370 101.350 ;
        RECT 130.560 101.180 130.730 101.350 ;
        RECT 131.400 101.180 131.570 101.350 ;
        RECT 131.760 101.180 131.930 101.350 ;
        RECT 132.120 101.180 132.290 101.350 ;
        RECT 133.710 101.190 133.880 101.360 ;
        RECT 134.150 101.190 134.320 101.360 ;
        RECT 134.560 101.190 134.730 101.360 ;
        RECT 134.990 101.190 135.160 101.360 ;
        RECT 135.430 101.190 135.600 101.360 ;
        RECT 135.840 101.190 136.010 101.360 ;
        RECT 137.550 101.190 137.720 101.360 ;
        RECT 137.990 101.190 138.160 101.360 ;
        RECT 138.400 101.190 138.570 101.360 ;
        RECT 138.830 101.190 139.000 101.360 ;
        RECT 139.270 101.190 139.440 101.360 ;
        RECT 139.680 101.190 139.850 101.360 ;
        RECT 5.920 93.520 6.090 93.700 ;
        RECT 6.400 93.520 6.570 93.700 ;
        RECT 6.880 93.520 7.050 93.700 ;
        RECT 7.360 93.520 7.530 93.700 ;
        RECT 7.840 93.520 8.010 93.700 ;
        RECT 8.320 93.520 8.490 93.700 ;
        RECT 8.800 93.520 8.970 93.700 ;
        RECT 9.280 93.520 9.450 93.700 ;
        RECT 9.760 93.520 9.930 93.700 ;
        RECT 10.240 93.520 10.410 93.700 ;
        RECT 10.720 93.520 10.890 93.700 ;
        RECT 11.200 93.520 11.370 93.700 ;
        RECT 11.680 93.520 11.850 93.700 ;
        RECT 12.160 93.520 12.330 93.700 ;
        RECT 12.640 93.520 12.810 93.700 ;
        RECT 13.120 93.520 13.290 93.700 ;
        RECT 13.600 93.520 13.770 93.700 ;
        RECT 14.080 93.520 14.250 93.700 ;
        RECT 14.560 93.520 14.730 93.700 ;
        RECT 15.040 93.520 15.210 93.700 ;
        RECT 15.520 93.520 15.690 93.700 ;
        RECT 16.000 93.520 16.170 93.700 ;
        RECT 16.480 93.520 16.650 93.700 ;
        RECT 16.960 93.520 17.130 93.700 ;
        RECT 17.440 93.520 17.610 93.700 ;
        RECT 17.920 93.520 18.090 93.700 ;
        RECT 18.400 93.520 18.570 93.700 ;
        RECT 18.880 93.520 19.050 93.700 ;
        RECT 19.360 93.520 19.530 93.700 ;
        RECT 19.840 93.520 20.010 93.700 ;
        RECT 20.320 93.520 20.490 93.700 ;
        RECT 20.800 93.520 20.970 93.700 ;
        RECT 21.280 93.520 21.450 93.700 ;
        RECT 21.760 93.520 21.930 93.700 ;
        RECT 22.240 93.520 22.410 93.700 ;
        RECT 22.720 93.520 22.890 93.700 ;
        RECT 23.200 93.520 23.370 93.700 ;
        RECT 23.680 93.520 23.850 93.700 ;
        RECT 24.160 93.520 24.330 93.700 ;
        RECT 24.640 93.520 24.810 93.700 ;
        RECT 25.120 93.520 25.290 93.700 ;
        RECT 25.600 93.520 25.770 93.700 ;
        RECT 26.080 93.520 26.250 93.700 ;
        RECT 26.560 93.520 26.730 93.700 ;
        RECT 27.040 93.520 27.210 93.700 ;
        RECT 27.520 93.520 27.690 93.700 ;
        RECT 28.000 93.520 28.170 93.700 ;
        RECT 28.480 93.520 28.650 93.700 ;
        RECT 28.960 93.520 29.130 93.700 ;
        RECT 29.440 93.520 29.610 93.700 ;
        RECT 29.920 93.520 30.090 93.700 ;
        RECT 30.400 93.520 30.570 93.700 ;
        RECT 30.880 93.520 31.050 93.700 ;
        RECT 31.360 93.520 31.530 93.700 ;
        RECT 31.840 93.520 32.010 93.700 ;
        RECT 32.320 93.520 32.490 93.700 ;
      LAYER li1 ;
        RECT 32.640 93.520 33.120 93.700 ;
      LAYER li1 ;
        RECT 33.280 93.520 33.450 93.700 ;
        RECT 33.760 93.520 33.930 93.700 ;
        RECT 34.240 93.520 34.410 93.700 ;
        RECT 34.720 93.520 34.890 93.700 ;
        RECT 35.200 93.520 35.370 93.700 ;
        RECT 35.680 93.520 35.850 93.700 ;
        RECT 36.160 93.520 36.330 93.700 ;
        RECT 36.640 93.520 36.810 93.700 ;
        RECT 37.120 93.520 37.290 93.700 ;
        RECT 37.600 93.520 37.770 93.700 ;
        RECT 38.080 93.520 38.250 93.700 ;
        RECT 38.560 93.520 38.730 93.700 ;
        RECT 39.040 93.520 39.210 93.700 ;
        RECT 39.520 93.520 39.690 93.700 ;
        RECT 40.000 93.520 40.170 93.700 ;
        RECT 40.480 93.520 40.650 93.700 ;
        RECT 40.960 93.520 41.130 93.700 ;
        RECT 41.440 93.520 41.610 93.700 ;
        RECT 41.920 93.520 42.090 93.700 ;
        RECT 42.400 93.520 42.570 93.700 ;
        RECT 42.880 93.520 43.050 93.700 ;
        RECT 43.360 93.520 43.530 93.700 ;
        RECT 43.840 93.520 44.010 93.700 ;
        RECT 44.320 93.520 44.490 93.700 ;
        RECT 44.800 93.520 44.970 93.700 ;
        RECT 45.280 93.520 45.450 93.700 ;
        RECT 45.760 93.520 45.930 93.700 ;
        RECT 46.240 93.520 46.410 93.700 ;
        RECT 46.720 93.520 46.890 93.700 ;
        RECT 47.200 93.520 47.370 93.700 ;
        RECT 47.680 93.520 47.850 93.700 ;
        RECT 48.160 93.520 48.330 93.700 ;
        RECT 48.640 93.520 48.810 93.700 ;
        RECT 49.120 93.520 49.290 93.700 ;
        RECT 49.600 93.520 49.770 93.700 ;
        RECT 50.080 93.520 50.250 93.700 ;
        RECT 50.560 93.520 50.730 93.700 ;
        RECT 51.040 93.520 51.210 93.700 ;
        RECT 51.520 93.520 51.690 93.700 ;
        RECT 52.000 93.520 52.170 93.700 ;
        RECT 52.480 93.520 52.650 93.700 ;
        RECT 52.960 93.520 53.130 93.700 ;
        RECT 53.440 93.520 53.610 93.700 ;
        RECT 53.920 93.520 54.090 93.700 ;
        RECT 54.400 93.520 54.570 93.700 ;
        RECT 54.880 93.520 55.050 93.700 ;
        RECT 55.360 93.520 55.530 93.700 ;
        RECT 55.840 93.520 56.010 93.700 ;
        RECT 56.320 93.520 56.490 93.700 ;
        RECT 56.800 93.520 56.970 93.700 ;
        RECT 57.280 93.520 57.450 93.700 ;
        RECT 57.760 93.520 57.930 93.700 ;
        RECT 58.240 93.520 58.410 93.700 ;
        RECT 58.720 93.520 58.890 93.700 ;
        RECT 59.200 93.520 59.370 93.700 ;
        RECT 59.680 93.520 59.850 93.700 ;
        RECT 60.160 93.520 60.330 93.700 ;
        RECT 60.640 93.520 60.810 93.700 ;
        RECT 61.120 93.520 61.290 93.700 ;
        RECT 61.600 93.520 61.770 93.700 ;
        RECT 62.080 93.520 62.250 93.700 ;
        RECT 62.560 93.520 62.730 93.700 ;
        RECT 63.040 93.520 63.210 93.700 ;
        RECT 63.520 93.520 63.690 93.700 ;
        RECT 64.000 93.520 64.170 93.700 ;
        RECT 64.480 93.520 64.650 93.700 ;
        RECT 64.960 93.520 65.130 93.700 ;
        RECT 65.440 93.520 65.610 93.700 ;
        RECT 65.920 93.520 66.090 93.700 ;
        RECT 66.400 93.520 66.570 93.700 ;
        RECT 66.880 93.520 67.050 93.700 ;
        RECT 67.360 93.520 67.530 93.700 ;
        RECT 67.840 93.520 68.010 93.700 ;
        RECT 68.320 93.520 68.490 93.700 ;
        RECT 68.800 93.520 68.970 93.700 ;
        RECT 69.280 93.520 69.450 93.700 ;
        RECT 69.760 93.520 69.930 93.700 ;
        RECT 70.240 93.520 70.410 93.700 ;
        RECT 70.720 93.520 70.890 93.700 ;
        RECT 71.200 93.520 71.370 93.700 ;
        RECT 71.680 93.520 71.850 93.700 ;
        RECT 72.160 93.520 72.330 93.700 ;
        RECT 72.640 93.520 72.810 93.700 ;
        RECT 73.120 93.520 73.290 93.700 ;
        RECT 73.600 93.520 73.770 93.700 ;
      LAYER li1 ;
        RECT 73.920 93.520 74.400 93.700 ;
      LAYER li1 ;
        RECT 74.560 93.520 74.730 93.700 ;
        RECT 75.040 93.520 75.210 93.700 ;
        RECT 75.520 93.520 75.690 93.700 ;
        RECT 76.000 93.520 76.170 93.700 ;
        RECT 76.480 93.520 76.650 93.700 ;
        RECT 76.960 93.520 77.130 93.700 ;
        RECT 77.440 93.520 77.610 93.700 ;
        RECT 77.920 93.520 78.090 93.700 ;
        RECT 78.400 93.520 78.570 93.700 ;
        RECT 78.880 93.520 79.050 93.700 ;
        RECT 79.360 93.520 79.530 93.700 ;
        RECT 79.840 93.520 80.010 93.700 ;
        RECT 80.320 93.520 80.490 93.700 ;
        RECT 80.800 93.520 80.970 93.700 ;
        RECT 81.280 93.520 81.450 93.700 ;
        RECT 81.760 93.520 81.930 93.700 ;
        RECT 82.240 93.520 82.410 93.700 ;
        RECT 82.720 93.520 82.890 93.700 ;
        RECT 83.200 93.520 83.370 93.700 ;
        RECT 83.680 93.520 83.850 93.700 ;
        RECT 84.160 93.520 84.330 93.700 ;
        RECT 84.640 93.520 84.810 93.700 ;
        RECT 85.120 93.520 85.290 93.700 ;
        RECT 85.600 93.520 85.770 93.700 ;
        RECT 86.080 93.520 86.250 93.700 ;
        RECT 86.560 93.520 86.730 93.700 ;
        RECT 87.040 93.520 87.210 93.700 ;
        RECT 87.520 93.520 87.690 93.700 ;
        RECT 88.000 93.520 88.170 93.700 ;
        RECT 88.480 93.520 88.650 93.700 ;
        RECT 88.960 93.520 89.130 93.700 ;
        RECT 89.440 93.520 89.610 93.700 ;
        RECT 89.920 93.520 90.090 93.700 ;
        RECT 90.400 93.520 90.570 93.700 ;
        RECT 90.880 93.520 91.050 93.700 ;
        RECT 91.360 93.520 91.530 93.700 ;
        RECT 91.840 93.520 92.010 93.700 ;
        RECT 92.320 93.520 92.490 93.700 ;
        RECT 92.800 93.520 92.970 93.700 ;
        RECT 93.280 93.520 93.450 93.700 ;
        RECT 93.760 93.520 93.930 93.700 ;
        RECT 94.240 93.520 94.410 93.700 ;
        RECT 94.720 93.520 94.890 93.700 ;
        RECT 95.200 93.520 95.370 93.700 ;
        RECT 95.680 93.520 95.850 93.700 ;
        RECT 96.160 93.520 96.330 93.700 ;
        RECT 96.640 93.520 96.810 93.700 ;
        RECT 97.120 93.520 97.290 93.700 ;
        RECT 97.600 93.520 97.770 93.700 ;
        RECT 98.080 93.520 98.250 93.700 ;
      LAYER li1 ;
        RECT 98.400 93.520 98.880 93.700 ;
      LAYER li1 ;
        RECT 99.040 93.520 99.210 93.700 ;
        RECT 99.520 93.520 99.690 93.700 ;
        RECT 100.000 93.520 100.170 93.700 ;
        RECT 100.480 93.520 100.650 93.700 ;
        RECT 100.960 93.520 101.130 93.700 ;
        RECT 101.440 93.520 101.610 93.700 ;
        RECT 101.920 93.520 102.090 93.700 ;
        RECT 102.400 93.520 102.570 93.700 ;
        RECT 102.880 93.520 103.050 93.700 ;
        RECT 103.360 93.520 103.530 93.700 ;
        RECT 103.840 93.520 104.010 93.700 ;
        RECT 104.320 93.520 104.490 93.700 ;
        RECT 104.800 93.520 104.970 93.700 ;
        RECT 105.280 93.520 105.450 93.700 ;
        RECT 105.760 93.520 105.930 93.700 ;
        RECT 106.240 93.520 106.410 93.700 ;
        RECT 106.720 93.520 106.890 93.700 ;
        RECT 107.200 93.520 107.370 93.700 ;
        RECT 107.680 93.520 107.850 93.700 ;
        RECT 108.160 93.520 108.330 93.700 ;
        RECT 108.640 93.520 108.810 93.700 ;
        RECT 109.120 93.520 109.290 93.700 ;
        RECT 109.600 93.520 109.770 93.700 ;
        RECT 110.080 93.520 110.250 93.700 ;
        RECT 110.560 93.520 110.730 93.700 ;
        RECT 111.040 93.520 111.210 93.700 ;
        RECT 111.520 93.520 111.690 93.700 ;
        RECT 112.000 93.520 112.170 93.700 ;
        RECT 112.480 93.520 112.650 93.700 ;
        RECT 112.960 93.520 113.130 93.700 ;
        RECT 113.440 93.520 113.610 93.700 ;
        RECT 113.920 93.520 114.090 93.700 ;
        RECT 114.400 93.520 114.570 93.700 ;
        RECT 114.880 93.520 115.050 93.700 ;
        RECT 115.360 93.520 115.530 93.700 ;
        RECT 115.840 93.520 116.010 93.700 ;
        RECT 116.320 93.520 116.490 93.700 ;
        RECT 116.800 93.520 116.970 93.700 ;
        RECT 117.280 93.520 117.450 93.700 ;
        RECT 117.760 93.520 117.930 93.700 ;
        RECT 118.240 93.520 118.410 93.700 ;
        RECT 118.720 93.520 118.890 93.700 ;
        RECT 119.200 93.520 119.370 93.700 ;
        RECT 119.680 93.520 119.850 93.700 ;
        RECT 120.160 93.520 120.330 93.700 ;
        RECT 120.640 93.520 120.810 93.700 ;
      LAYER li1 ;
        RECT 120.960 93.520 121.440 93.700 ;
      LAYER li1 ;
        RECT 121.600 93.520 121.770 93.700 ;
        RECT 122.080 93.520 122.250 93.700 ;
        RECT 122.560 93.520 122.730 93.700 ;
        RECT 123.040 93.520 123.210 93.700 ;
        RECT 123.520 93.520 123.690 93.700 ;
        RECT 124.000 93.520 124.170 93.700 ;
        RECT 124.480 93.520 124.650 93.700 ;
        RECT 124.960 93.520 125.130 93.700 ;
        RECT 125.440 93.520 125.610 93.700 ;
        RECT 125.920 93.520 126.090 93.700 ;
        RECT 126.400 93.520 126.570 93.700 ;
        RECT 126.880 93.520 127.050 93.700 ;
        RECT 127.360 93.520 127.530 93.700 ;
        RECT 127.840 93.520 128.010 93.700 ;
        RECT 128.320 93.520 128.490 93.700 ;
        RECT 128.800 93.520 128.970 93.700 ;
        RECT 129.280 93.520 129.450 93.700 ;
        RECT 129.760 93.520 129.930 93.700 ;
        RECT 130.240 93.520 130.410 93.700 ;
        RECT 130.720 93.520 130.890 93.700 ;
        RECT 131.200 93.520 131.370 93.700 ;
        RECT 131.680 93.520 131.850 93.700 ;
        RECT 132.160 93.520 132.330 93.700 ;
        RECT 132.640 93.520 132.810 93.700 ;
        RECT 133.120 93.520 133.290 93.700 ;
        RECT 133.600 93.520 133.770 93.700 ;
        RECT 134.080 93.520 134.250 93.700 ;
        RECT 134.560 93.520 134.730 93.700 ;
        RECT 135.040 93.520 135.210 93.700 ;
        RECT 135.520 93.520 135.690 93.700 ;
        RECT 136.000 93.520 136.170 93.700 ;
        RECT 136.480 93.520 136.650 93.700 ;
        RECT 136.960 93.520 137.130 93.700 ;
        RECT 137.440 93.520 137.610 93.700 ;
        RECT 137.920 93.520 138.090 93.700 ;
        RECT 138.400 93.520 138.570 93.700 ;
        RECT 138.880 93.520 139.050 93.700 ;
        RECT 139.360 93.520 139.530 93.700 ;
        RECT 139.840 93.520 140.010 93.700 ;
        RECT 140.320 93.520 140.490 93.700 ;
        RECT 140.800 93.520 140.970 93.700 ;
        RECT 141.280 93.520 141.450 93.700 ;
        RECT 141.760 93.520 141.930 93.700 ;
        RECT 6.510 93.050 6.680 93.220 ;
        RECT 6.950 93.050 7.120 93.220 ;
        RECT 7.360 93.050 7.530 93.220 ;
        RECT 7.790 93.050 7.960 93.220 ;
        RECT 8.230 93.050 8.400 93.220 ;
        RECT 8.640 93.050 8.810 93.220 ;
        RECT 9.820 93.040 9.990 93.210 ;
        RECT 10.260 93.040 10.430 93.210 ;
        RECT 10.700 93.040 10.870 93.210 ;
        RECT 11.110 93.040 11.280 93.210 ;
        RECT 13.510 93.040 13.680 93.210 ;
        RECT 13.870 93.040 14.040 93.210 ;
        RECT 14.230 93.040 14.400 93.210 ;
        RECT 14.590 93.040 14.760 93.210 ;
        RECT 16.110 93.050 16.280 93.220 ;
        RECT 16.550 93.050 16.720 93.220 ;
        RECT 16.960 93.050 17.130 93.220 ;
        RECT 17.390 93.050 17.560 93.220 ;
        RECT 17.830 93.050 18.000 93.220 ;
        RECT 18.240 93.050 18.410 93.220 ;
        RECT 19.950 93.050 20.120 93.220 ;
        RECT 20.390 93.050 20.560 93.220 ;
        RECT 20.800 93.050 20.970 93.220 ;
        RECT 21.230 93.050 21.400 93.220 ;
        RECT 21.670 93.050 21.840 93.220 ;
        RECT 22.080 93.050 22.250 93.220 ;
        RECT 24.120 93.040 24.290 93.210 ;
        RECT 24.480 93.040 24.650 93.210 ;
        RECT 25.660 93.040 25.830 93.210 ;
        RECT 26.100 93.040 26.270 93.210 ;
        RECT 26.540 93.040 26.710 93.210 ;
        RECT 26.950 93.040 27.120 93.210 ;
        RECT 29.560 93.040 29.730 93.210 ;
        RECT 29.920 93.040 30.090 93.210 ;
        RECT 30.280 93.040 30.450 93.210 ;
        RECT 31.420 93.040 31.590 93.210 ;
        RECT 31.860 93.040 32.030 93.210 ;
        RECT 32.300 93.040 32.470 93.210 ;
        RECT 32.710 93.040 32.880 93.210 ;
        RECT 33.670 93.040 33.840 93.210 ;
        RECT 34.030 93.040 34.200 93.210 ;
        RECT 34.390 93.040 34.560 93.210 ;
        RECT 34.750 93.040 34.920 93.210 ;
        RECT 35.740 93.040 35.910 93.210 ;
        RECT 36.180 93.040 36.350 93.210 ;
        RECT 36.620 93.040 36.790 93.210 ;
        RECT 37.030 93.040 37.200 93.210 ;
        RECT 38.040 93.040 38.210 93.210 ;
        RECT 38.400 93.040 38.570 93.210 ;
        RECT 39.910 93.040 40.080 93.210 ;
        RECT 40.270 93.040 40.440 93.210 ;
        RECT 42.330 93.040 42.500 93.210 ;
        RECT 42.690 93.040 42.860 93.210 ;
        RECT 43.050 93.040 43.220 93.210 ;
        RECT 44.270 93.040 44.440 93.210 ;
        RECT 44.630 93.040 44.800 93.210 ;
        RECT 44.990 93.040 45.160 93.210 ;
        RECT 48.810 93.040 48.980 93.210 ;
        RECT 49.170 93.040 49.340 93.210 ;
        RECT 50.730 93.040 50.900 93.210 ;
        RECT 51.090 93.040 51.260 93.210 ;
        RECT 51.450 93.040 51.620 93.210 ;
        RECT 53.070 93.050 53.240 93.220 ;
        RECT 53.510 93.050 53.680 93.220 ;
        RECT 53.920 93.050 54.090 93.220 ;
        RECT 54.350 93.050 54.520 93.220 ;
        RECT 54.790 93.050 54.960 93.220 ;
        RECT 55.200 93.050 55.370 93.220 ;
        RECT 57.230 93.040 57.400 93.210 ;
        RECT 57.590 93.040 57.760 93.210 ;
        RECT 57.950 93.040 58.120 93.210 ;
        RECT 58.870 93.040 59.040 93.210 ;
        RECT 59.230 93.040 59.400 93.210 ;
        RECT 63.830 93.040 64.000 93.210 ;
        RECT 64.190 93.040 64.360 93.210 ;
        RECT 64.550 93.040 64.720 93.210 ;
        RECT 67.800 93.040 67.970 93.210 ;
        RECT 68.160 93.040 68.330 93.210 ;
        RECT 68.520 93.040 68.690 93.210 ;
        RECT 70.410 93.040 70.580 93.210 ;
        RECT 70.770 93.040 70.940 93.210 ;
        RECT 71.130 93.040 71.300 93.210 ;
        RECT 72.220 93.040 72.390 93.210 ;
        RECT 72.660 93.040 72.830 93.210 ;
        RECT 73.100 93.040 73.270 93.210 ;
        RECT 73.510 93.040 73.680 93.210 ;
        RECT 75.000 93.040 75.170 93.210 ;
        RECT 75.360 93.040 75.530 93.210 ;
        RECT 75.720 93.040 75.890 93.210 ;
        RECT 76.560 93.040 76.730 93.210 ;
        RECT 76.920 93.040 77.090 93.210 ;
        RECT 77.280 93.040 77.450 93.210 ;
        RECT 78.120 93.040 78.290 93.210 ;
        RECT 78.480 93.040 78.650 93.210 ;
        RECT 78.840 93.040 79.010 93.210 ;
        RECT 79.900 93.040 80.070 93.210 ;
        RECT 80.340 93.040 80.510 93.210 ;
        RECT 80.780 93.040 80.950 93.210 ;
        RECT 81.190 93.040 81.360 93.210 ;
        RECT 81.720 93.040 81.890 93.210 ;
        RECT 82.080 93.040 82.250 93.210 ;
        RECT 82.440 93.040 82.610 93.210 ;
        RECT 83.280 93.040 83.450 93.210 ;
        RECT 83.640 93.040 83.810 93.210 ;
        RECT 84.000 93.040 84.170 93.210 ;
        RECT 84.840 93.040 85.010 93.210 ;
        RECT 85.200 93.040 85.370 93.210 ;
        RECT 85.560 93.040 85.730 93.210 ;
        RECT 86.620 93.040 86.790 93.210 ;
        RECT 87.060 93.040 87.230 93.210 ;
        RECT 87.500 93.040 87.670 93.210 ;
        RECT 87.910 93.040 88.080 93.210 ;
        RECT 88.440 93.040 88.610 93.210 ;
        RECT 88.800 93.040 88.970 93.210 ;
        RECT 89.160 93.040 89.330 93.210 ;
        RECT 90.000 93.040 90.170 93.210 ;
        RECT 90.360 93.040 90.530 93.210 ;
        RECT 90.720 93.040 90.890 93.210 ;
        RECT 91.560 93.040 91.730 93.210 ;
        RECT 91.920 93.040 92.090 93.210 ;
        RECT 92.280 93.040 92.450 93.210 ;
        RECT 93.340 93.040 93.510 93.210 ;
        RECT 93.780 93.040 93.950 93.210 ;
        RECT 94.220 93.040 94.390 93.210 ;
        RECT 94.630 93.040 94.800 93.210 ;
        RECT 95.160 93.040 95.330 93.210 ;
        RECT 95.520 93.040 95.690 93.210 ;
        RECT 95.880 93.040 96.050 93.210 ;
        RECT 96.720 93.040 96.890 93.210 ;
        RECT 97.080 93.040 97.250 93.210 ;
        RECT 97.440 93.040 97.610 93.210 ;
        RECT 98.280 93.040 98.450 93.210 ;
        RECT 98.640 93.040 98.810 93.210 ;
        RECT 99.000 93.040 99.170 93.210 ;
        RECT 100.060 93.040 100.230 93.210 ;
        RECT 100.500 93.040 100.670 93.210 ;
        RECT 100.940 93.040 101.110 93.210 ;
        RECT 101.350 93.040 101.520 93.210 ;
        RECT 101.880 93.040 102.050 93.210 ;
        RECT 102.240 93.040 102.410 93.210 ;
        RECT 102.600 93.040 102.770 93.210 ;
        RECT 103.440 93.040 103.610 93.210 ;
        RECT 103.800 93.040 103.970 93.210 ;
        RECT 104.160 93.040 104.330 93.210 ;
        RECT 105.000 93.040 105.170 93.210 ;
        RECT 105.360 93.040 105.530 93.210 ;
        RECT 105.720 93.040 105.890 93.210 ;
        RECT 106.780 93.040 106.950 93.210 ;
        RECT 107.220 93.040 107.390 93.210 ;
        RECT 107.660 93.040 107.830 93.210 ;
        RECT 108.070 93.040 108.240 93.210 ;
        RECT 109.120 93.040 109.290 93.210 ;
        RECT 109.480 93.040 109.650 93.210 ;
        RECT 109.840 93.040 110.010 93.210 ;
        RECT 112.060 93.040 112.230 93.210 ;
        RECT 112.500 93.040 112.670 93.210 ;
        RECT 112.940 93.040 113.110 93.210 ;
        RECT 113.350 93.040 113.520 93.210 ;
        RECT 113.880 93.040 114.050 93.210 ;
        RECT 114.240 93.040 114.410 93.210 ;
        RECT 115.420 93.040 115.590 93.210 ;
        RECT 115.860 93.040 116.030 93.210 ;
        RECT 116.300 93.040 116.470 93.210 ;
        RECT 116.710 93.040 116.880 93.210 ;
        RECT 117.670 93.040 117.840 93.210 ;
        RECT 118.030 93.040 118.200 93.210 ;
        RECT 118.390 93.040 118.560 93.210 ;
        RECT 118.750 93.040 118.920 93.210 ;
        RECT 119.740 93.040 119.910 93.210 ;
        RECT 120.180 93.040 120.350 93.210 ;
        RECT 120.620 93.040 120.790 93.210 ;
        RECT 121.030 93.040 121.200 93.210 ;
        RECT 121.560 93.040 121.730 93.210 ;
        RECT 121.920 93.040 122.090 93.210 ;
        RECT 122.280 93.040 122.450 93.210 ;
        RECT 123.120 93.040 123.290 93.210 ;
        RECT 123.480 93.040 123.650 93.210 ;
        RECT 123.840 93.040 124.010 93.210 ;
        RECT 124.680 93.040 124.850 93.210 ;
        RECT 125.040 93.040 125.210 93.210 ;
        RECT 125.400 93.040 125.570 93.210 ;
        RECT 126.990 93.050 127.160 93.220 ;
        RECT 127.430 93.050 127.600 93.220 ;
        RECT 127.840 93.050 128.010 93.220 ;
        RECT 128.270 93.050 128.440 93.220 ;
        RECT 128.710 93.050 128.880 93.220 ;
        RECT 129.120 93.050 129.290 93.220 ;
        RECT 130.830 93.050 131.000 93.220 ;
        RECT 131.270 93.050 131.440 93.220 ;
        RECT 131.680 93.050 131.850 93.220 ;
        RECT 132.110 93.050 132.280 93.220 ;
        RECT 132.550 93.050 132.720 93.220 ;
        RECT 132.960 93.050 133.130 93.220 ;
        RECT 134.670 93.050 134.840 93.220 ;
        RECT 135.110 93.050 135.280 93.220 ;
        RECT 135.520 93.050 135.690 93.220 ;
        RECT 135.950 93.050 136.120 93.220 ;
        RECT 136.390 93.050 136.560 93.220 ;
        RECT 136.800 93.050 136.970 93.220 ;
        RECT 138.510 93.050 138.680 93.220 ;
        RECT 138.950 93.050 139.120 93.220 ;
        RECT 139.360 93.050 139.530 93.220 ;
        RECT 139.790 93.050 139.960 93.220 ;
        RECT 140.230 93.050 140.400 93.220 ;
        RECT 140.640 93.050 140.810 93.220 ;
        RECT 5.920 85.380 6.090 85.560 ;
        RECT 6.400 85.380 6.570 85.560 ;
        RECT 6.880 85.380 7.050 85.560 ;
        RECT 7.360 85.380 7.530 85.560 ;
        RECT 7.840 85.380 8.010 85.560 ;
        RECT 8.320 85.380 8.490 85.560 ;
        RECT 8.800 85.380 8.970 85.560 ;
        RECT 9.280 85.380 9.450 85.560 ;
        RECT 9.760 85.380 9.930 85.560 ;
        RECT 10.240 85.380 10.410 85.560 ;
        RECT 10.720 85.380 10.890 85.560 ;
        RECT 11.200 85.380 11.370 85.560 ;
        RECT 11.680 85.380 11.850 85.560 ;
        RECT 12.160 85.380 12.330 85.560 ;
        RECT 12.640 85.380 12.810 85.560 ;
        RECT 13.120 85.380 13.290 85.560 ;
        RECT 13.600 85.380 13.770 85.560 ;
        RECT 14.080 85.380 14.250 85.560 ;
        RECT 14.560 85.380 14.730 85.560 ;
        RECT 15.040 85.380 15.210 85.560 ;
        RECT 15.520 85.380 15.690 85.560 ;
        RECT 16.000 85.380 16.170 85.560 ;
        RECT 16.480 85.380 16.650 85.560 ;
        RECT 16.960 85.380 17.130 85.560 ;
        RECT 17.440 85.380 17.610 85.560 ;
        RECT 17.920 85.380 18.090 85.560 ;
        RECT 18.400 85.380 18.570 85.560 ;
        RECT 18.880 85.380 19.050 85.560 ;
        RECT 19.360 85.380 19.530 85.560 ;
        RECT 19.840 85.380 20.010 85.560 ;
      LAYER li1 ;
        RECT 20.160 85.380 20.640 85.560 ;
      LAYER li1 ;
        RECT 20.800 85.380 20.970 85.560 ;
        RECT 21.280 85.380 21.450 85.560 ;
        RECT 21.760 85.380 21.930 85.560 ;
        RECT 22.240 85.380 22.410 85.560 ;
        RECT 22.720 85.380 22.890 85.560 ;
        RECT 23.200 85.380 23.370 85.560 ;
        RECT 23.680 85.380 23.850 85.560 ;
        RECT 24.160 85.380 24.330 85.560 ;
        RECT 24.640 85.380 24.810 85.560 ;
        RECT 25.120 85.380 25.290 85.560 ;
        RECT 25.600 85.380 25.770 85.560 ;
        RECT 26.080 85.380 26.250 85.560 ;
        RECT 26.560 85.380 26.730 85.560 ;
        RECT 27.040 85.380 27.210 85.560 ;
        RECT 27.520 85.380 27.690 85.560 ;
        RECT 28.000 85.380 28.170 85.560 ;
        RECT 28.480 85.380 28.650 85.560 ;
        RECT 28.960 85.380 29.130 85.560 ;
        RECT 29.440 85.380 29.610 85.560 ;
        RECT 29.920 85.380 30.090 85.560 ;
        RECT 30.400 85.380 30.570 85.560 ;
        RECT 30.880 85.380 31.050 85.560 ;
        RECT 31.360 85.380 31.530 85.560 ;
        RECT 31.840 85.380 32.010 85.560 ;
        RECT 32.320 85.380 32.490 85.560 ;
        RECT 32.800 85.380 32.970 85.560 ;
        RECT 33.280 85.380 33.450 85.560 ;
        RECT 33.760 85.380 33.930 85.560 ;
        RECT 34.240 85.380 34.410 85.560 ;
        RECT 34.720 85.380 34.890 85.560 ;
        RECT 35.200 85.380 35.370 85.560 ;
        RECT 35.680 85.380 35.850 85.560 ;
        RECT 36.160 85.380 36.330 85.560 ;
        RECT 36.640 85.380 36.810 85.560 ;
        RECT 37.120 85.380 37.290 85.560 ;
        RECT 37.600 85.380 37.770 85.560 ;
        RECT 38.080 85.380 38.250 85.560 ;
        RECT 38.560 85.380 38.730 85.560 ;
        RECT 39.040 85.380 39.210 85.560 ;
        RECT 39.520 85.380 39.690 85.560 ;
        RECT 40.000 85.380 40.170 85.560 ;
        RECT 40.480 85.380 40.650 85.560 ;
        RECT 40.960 85.380 41.130 85.560 ;
        RECT 41.440 85.380 41.610 85.560 ;
        RECT 41.920 85.380 42.090 85.560 ;
        RECT 42.400 85.380 42.570 85.560 ;
        RECT 42.880 85.380 43.050 85.560 ;
        RECT 43.360 85.380 43.530 85.560 ;
        RECT 43.840 85.380 44.010 85.560 ;
        RECT 44.320 85.380 44.490 85.560 ;
        RECT 44.800 85.380 44.970 85.560 ;
        RECT 45.280 85.380 45.450 85.560 ;
        RECT 45.760 85.380 45.930 85.560 ;
        RECT 46.240 85.380 46.410 85.560 ;
        RECT 46.720 85.380 46.890 85.560 ;
        RECT 47.200 85.380 47.370 85.560 ;
        RECT 47.680 85.380 47.850 85.560 ;
        RECT 48.160 85.380 48.330 85.560 ;
        RECT 48.640 85.380 48.810 85.560 ;
        RECT 49.120 85.380 49.290 85.560 ;
        RECT 49.600 85.380 49.770 85.560 ;
        RECT 50.080 85.380 50.250 85.560 ;
        RECT 50.560 85.380 50.730 85.560 ;
        RECT 51.040 85.380 51.210 85.560 ;
        RECT 51.520 85.380 51.690 85.560 ;
        RECT 52.000 85.380 52.170 85.560 ;
        RECT 52.480 85.380 52.650 85.560 ;
        RECT 52.960 85.380 53.130 85.560 ;
        RECT 53.440 85.380 53.610 85.560 ;
        RECT 53.920 85.380 54.090 85.560 ;
        RECT 54.400 85.380 54.570 85.560 ;
        RECT 54.880 85.380 55.050 85.560 ;
        RECT 55.360 85.380 55.530 85.560 ;
        RECT 55.840 85.380 56.010 85.560 ;
        RECT 56.320 85.380 56.490 85.560 ;
        RECT 56.800 85.380 56.970 85.560 ;
        RECT 57.280 85.380 57.450 85.560 ;
        RECT 57.760 85.380 57.930 85.560 ;
        RECT 58.240 85.380 58.410 85.560 ;
        RECT 58.720 85.380 58.890 85.560 ;
        RECT 59.200 85.380 59.370 85.560 ;
        RECT 59.680 85.380 59.850 85.560 ;
        RECT 60.160 85.380 60.330 85.560 ;
        RECT 60.640 85.380 60.810 85.560 ;
        RECT 61.120 85.380 61.290 85.560 ;
        RECT 61.600 85.380 61.770 85.560 ;
        RECT 62.080 85.380 62.250 85.560 ;
        RECT 62.560 85.380 62.730 85.560 ;
        RECT 63.040 85.380 63.210 85.560 ;
        RECT 63.520 85.380 63.690 85.560 ;
        RECT 64.000 85.380 64.170 85.560 ;
        RECT 64.480 85.380 64.650 85.560 ;
        RECT 64.960 85.380 65.130 85.560 ;
        RECT 65.440 85.380 65.610 85.560 ;
        RECT 65.920 85.380 66.090 85.560 ;
        RECT 66.400 85.380 66.570 85.560 ;
        RECT 66.880 85.380 67.050 85.560 ;
        RECT 67.360 85.380 67.530 85.560 ;
        RECT 67.840 85.380 68.010 85.560 ;
      LAYER li1 ;
        RECT 68.160 85.380 68.640 85.560 ;
      LAYER li1 ;
        RECT 68.800 85.380 68.970 85.560 ;
        RECT 69.280 85.380 69.450 85.560 ;
        RECT 69.760 85.380 69.930 85.560 ;
        RECT 70.240 85.380 70.410 85.560 ;
        RECT 70.720 85.380 70.890 85.560 ;
        RECT 71.200 85.380 71.370 85.560 ;
        RECT 71.680 85.380 71.850 85.560 ;
        RECT 72.160 85.380 72.330 85.560 ;
        RECT 72.640 85.380 72.810 85.560 ;
        RECT 73.120 85.380 73.290 85.560 ;
        RECT 73.600 85.380 73.770 85.560 ;
        RECT 74.080 85.380 74.250 85.560 ;
        RECT 74.560 85.380 74.730 85.560 ;
        RECT 75.040 85.380 75.210 85.560 ;
        RECT 75.520 85.380 75.690 85.560 ;
        RECT 76.000 85.380 76.170 85.560 ;
        RECT 76.480 85.380 76.650 85.560 ;
        RECT 76.960 85.380 77.130 85.560 ;
        RECT 77.440 85.380 77.610 85.560 ;
        RECT 77.920 85.380 78.090 85.560 ;
        RECT 78.400 85.380 78.570 85.560 ;
        RECT 78.880 85.380 79.050 85.560 ;
        RECT 79.360 85.380 79.530 85.560 ;
        RECT 79.840 85.380 80.010 85.560 ;
        RECT 80.320 85.380 80.490 85.560 ;
        RECT 80.800 85.380 80.970 85.560 ;
        RECT 81.280 85.380 81.450 85.560 ;
        RECT 81.760 85.380 81.930 85.560 ;
        RECT 82.240 85.380 82.410 85.560 ;
        RECT 82.720 85.380 82.890 85.560 ;
        RECT 83.200 85.380 83.370 85.560 ;
        RECT 83.680 85.380 83.850 85.560 ;
        RECT 84.160 85.380 84.330 85.560 ;
        RECT 84.640 85.380 84.810 85.560 ;
        RECT 85.120 85.380 85.290 85.560 ;
        RECT 85.600 85.380 85.770 85.560 ;
        RECT 86.080 85.380 86.250 85.560 ;
        RECT 86.560 85.380 86.730 85.560 ;
        RECT 87.040 85.380 87.210 85.560 ;
        RECT 87.520 85.380 87.690 85.560 ;
        RECT 88.000 85.380 88.170 85.560 ;
        RECT 88.480 85.380 88.650 85.560 ;
        RECT 88.960 85.380 89.130 85.560 ;
        RECT 89.440 85.380 89.610 85.560 ;
        RECT 89.920 85.380 90.090 85.560 ;
        RECT 90.400 85.380 90.570 85.560 ;
        RECT 90.880 85.380 91.050 85.560 ;
        RECT 91.360 85.380 91.530 85.560 ;
        RECT 91.840 85.380 92.010 85.560 ;
        RECT 92.320 85.380 92.490 85.560 ;
        RECT 92.800 85.380 92.970 85.560 ;
        RECT 93.280 85.380 93.450 85.560 ;
        RECT 93.760 85.380 93.930 85.560 ;
        RECT 94.240 85.380 94.410 85.560 ;
        RECT 94.720 85.380 94.890 85.560 ;
        RECT 95.200 85.380 95.370 85.560 ;
        RECT 95.680 85.380 95.850 85.560 ;
        RECT 96.160 85.380 96.330 85.560 ;
        RECT 96.640 85.380 96.810 85.560 ;
        RECT 97.120 85.380 97.290 85.560 ;
        RECT 97.600 85.380 97.770 85.560 ;
        RECT 98.080 85.380 98.250 85.560 ;
        RECT 98.560 85.380 98.730 85.560 ;
        RECT 99.040 85.380 99.210 85.560 ;
        RECT 99.520 85.380 99.690 85.560 ;
        RECT 100.000 85.380 100.170 85.560 ;
        RECT 100.480 85.380 100.650 85.560 ;
        RECT 100.960 85.380 101.130 85.560 ;
      LAYER li1 ;
        RECT 101.280 85.380 101.760 85.560 ;
      LAYER li1 ;
        RECT 101.920 85.380 102.090 85.560 ;
        RECT 102.400 85.380 102.570 85.560 ;
        RECT 102.880 85.380 103.050 85.560 ;
        RECT 103.360 85.380 103.530 85.560 ;
        RECT 103.840 85.380 104.010 85.560 ;
        RECT 104.320 85.380 104.490 85.560 ;
        RECT 104.800 85.380 104.970 85.560 ;
        RECT 105.280 85.380 105.450 85.560 ;
        RECT 105.760 85.380 105.930 85.560 ;
        RECT 106.240 85.380 106.410 85.560 ;
        RECT 106.720 85.380 106.890 85.560 ;
        RECT 107.200 85.380 107.370 85.560 ;
        RECT 107.680 85.380 107.850 85.560 ;
        RECT 108.160 85.380 108.330 85.560 ;
        RECT 108.640 85.380 108.810 85.560 ;
        RECT 109.120 85.380 109.290 85.560 ;
        RECT 109.600 85.380 109.770 85.560 ;
        RECT 110.080 85.380 110.250 85.560 ;
        RECT 110.560 85.380 110.730 85.560 ;
        RECT 111.040 85.380 111.210 85.560 ;
        RECT 111.520 85.380 111.690 85.560 ;
        RECT 112.000 85.380 112.170 85.560 ;
        RECT 112.480 85.380 112.650 85.560 ;
        RECT 112.960 85.380 113.130 85.560 ;
        RECT 113.440 85.380 113.610 85.560 ;
        RECT 113.920 85.380 114.090 85.560 ;
        RECT 114.400 85.380 114.570 85.560 ;
        RECT 114.880 85.380 115.050 85.560 ;
        RECT 115.360 85.380 115.530 85.560 ;
        RECT 115.840 85.380 116.010 85.560 ;
        RECT 116.320 85.380 116.490 85.560 ;
        RECT 116.800 85.380 116.970 85.560 ;
        RECT 117.280 85.380 117.450 85.560 ;
      LAYER li1 ;
        RECT 117.600 85.380 118.080 85.560 ;
      LAYER li1 ;
        RECT 118.240 85.380 118.410 85.560 ;
        RECT 118.720 85.380 118.890 85.560 ;
        RECT 119.200 85.380 119.370 85.560 ;
        RECT 119.680 85.380 119.850 85.560 ;
        RECT 120.160 85.380 120.330 85.560 ;
        RECT 120.640 85.380 120.810 85.560 ;
        RECT 121.120 85.380 121.290 85.560 ;
        RECT 121.600 85.380 121.770 85.560 ;
        RECT 122.080 85.380 122.250 85.560 ;
        RECT 122.560 85.380 122.730 85.560 ;
        RECT 123.040 85.380 123.210 85.560 ;
        RECT 123.520 85.380 123.690 85.560 ;
        RECT 124.000 85.380 124.170 85.560 ;
        RECT 124.480 85.380 124.650 85.560 ;
        RECT 124.960 85.380 125.130 85.560 ;
        RECT 125.440 85.380 125.610 85.560 ;
        RECT 125.920 85.380 126.090 85.560 ;
        RECT 126.400 85.380 126.570 85.560 ;
        RECT 126.880 85.380 127.050 85.560 ;
        RECT 127.360 85.380 127.530 85.560 ;
        RECT 127.840 85.380 128.010 85.560 ;
        RECT 128.320 85.380 128.490 85.560 ;
        RECT 128.800 85.380 128.970 85.560 ;
        RECT 129.280 85.380 129.450 85.560 ;
        RECT 129.760 85.380 129.930 85.560 ;
        RECT 130.240 85.380 130.410 85.560 ;
        RECT 130.720 85.380 130.890 85.560 ;
        RECT 131.200 85.380 131.370 85.560 ;
        RECT 131.680 85.380 131.850 85.560 ;
        RECT 132.160 85.380 132.330 85.560 ;
        RECT 132.640 85.380 132.810 85.560 ;
        RECT 133.120 85.380 133.290 85.560 ;
        RECT 133.600 85.380 133.770 85.560 ;
      LAYER li1 ;
        RECT 133.920 85.380 134.400 85.560 ;
      LAYER li1 ;
        RECT 134.560 85.380 134.730 85.560 ;
        RECT 135.040 85.380 135.210 85.560 ;
        RECT 135.520 85.380 135.690 85.560 ;
        RECT 136.000 85.380 136.170 85.560 ;
        RECT 136.480 85.380 136.650 85.560 ;
        RECT 136.960 85.380 137.130 85.560 ;
        RECT 137.440 85.380 137.610 85.560 ;
        RECT 137.920 85.380 138.090 85.560 ;
        RECT 138.400 85.380 138.570 85.560 ;
        RECT 138.880 85.380 139.050 85.560 ;
        RECT 139.360 85.380 139.530 85.560 ;
        RECT 139.840 85.380 140.010 85.560 ;
        RECT 140.320 85.380 140.490 85.560 ;
        RECT 140.800 85.380 140.970 85.560 ;
        RECT 141.280 85.380 141.450 85.560 ;
      LAYER li1 ;
        RECT 141.600 85.380 142.080 85.560 ;
      LAYER li1 ;
        RECT 5.980 84.900 6.150 85.070 ;
        RECT 6.420 84.900 6.590 85.070 ;
        RECT 6.860 84.900 7.030 85.070 ;
        RECT 7.270 84.900 7.440 85.070 ;
        RECT 8.270 84.900 8.440 85.070 ;
        RECT 8.630 84.900 8.800 85.070 ;
        RECT 8.990 84.900 9.160 85.070 ;
        RECT 9.910 84.900 10.080 85.070 ;
        RECT 10.270 84.900 10.440 85.070 ;
        RECT 14.870 84.900 15.040 85.070 ;
        RECT 15.230 84.900 15.400 85.070 ;
        RECT 15.590 84.900 15.760 85.070 ;
        RECT 18.840 84.900 19.010 85.070 ;
        RECT 19.200 84.900 19.370 85.070 ;
        RECT 19.560 84.900 19.730 85.070 ;
        RECT 21.450 84.900 21.620 85.070 ;
        RECT 21.810 84.900 21.980 85.070 ;
        RECT 22.170 84.900 22.340 85.070 ;
        RECT 23.260 84.900 23.430 85.070 ;
        RECT 23.700 84.900 23.870 85.070 ;
        RECT 24.140 84.900 24.310 85.070 ;
        RECT 24.550 84.900 24.720 85.070 ;
        RECT 25.510 84.900 25.680 85.070 ;
        RECT 25.870 84.900 26.040 85.070 ;
        RECT 26.230 84.900 26.400 85.070 ;
        RECT 26.590 84.900 26.760 85.070 ;
        RECT 27.580 84.900 27.750 85.070 ;
        RECT 28.020 84.900 28.190 85.070 ;
        RECT 28.460 84.900 28.630 85.070 ;
        RECT 28.870 84.900 29.040 85.070 ;
        RECT 31.480 84.900 31.650 85.070 ;
        RECT 31.840 84.900 32.010 85.070 ;
        RECT 32.200 84.900 32.370 85.070 ;
        RECT 33.340 84.900 33.510 85.070 ;
        RECT 33.780 84.900 33.950 85.070 ;
        RECT 34.220 84.900 34.390 85.070 ;
        RECT 34.630 84.900 34.800 85.070 ;
        RECT 35.590 84.900 35.760 85.070 ;
        RECT 35.950 84.900 36.120 85.070 ;
        RECT 36.310 84.900 36.480 85.070 ;
        RECT 36.670 84.900 36.840 85.070 ;
        RECT 37.660 84.900 37.830 85.070 ;
        RECT 38.100 84.900 38.270 85.070 ;
        RECT 38.540 84.900 38.710 85.070 ;
        RECT 38.950 84.900 39.120 85.070 ;
        RECT 39.480 84.900 39.650 85.070 ;
        RECT 39.840 84.900 40.010 85.070 ;
        RECT 40.200 84.900 40.370 85.070 ;
        RECT 41.040 84.900 41.210 85.070 ;
        RECT 41.400 84.900 41.570 85.070 ;
        RECT 41.760 84.900 41.930 85.070 ;
        RECT 42.600 84.900 42.770 85.070 ;
        RECT 42.960 84.900 43.130 85.070 ;
        RECT 43.320 84.900 43.490 85.070 ;
        RECT 44.910 84.910 45.080 85.080 ;
        RECT 45.350 84.910 45.520 85.080 ;
        RECT 45.760 84.910 45.930 85.080 ;
        RECT 46.190 84.910 46.360 85.080 ;
        RECT 46.630 84.910 46.800 85.080 ;
        RECT 47.040 84.910 47.210 85.080 ;
        RECT 49.080 84.900 49.250 85.070 ;
        RECT 49.440 84.900 49.610 85.070 ;
        RECT 49.800 84.900 49.970 85.070 ;
        RECT 50.640 84.900 50.810 85.070 ;
        RECT 51.000 84.900 51.170 85.070 ;
        RECT 51.360 84.900 51.530 85.070 ;
        RECT 52.200 84.900 52.370 85.070 ;
        RECT 52.560 84.900 52.730 85.070 ;
        RECT 52.920 84.900 53.090 85.070 ;
        RECT 53.980 84.900 54.150 85.070 ;
        RECT 54.420 84.900 54.590 85.070 ;
        RECT 54.860 84.900 55.030 85.070 ;
        RECT 55.270 84.900 55.440 85.070 ;
        RECT 55.800 84.900 55.970 85.070 ;
        RECT 56.160 84.900 56.330 85.070 ;
        RECT 56.520 84.900 56.690 85.070 ;
        RECT 57.360 84.900 57.530 85.070 ;
        RECT 57.720 84.900 57.890 85.070 ;
        RECT 58.080 84.900 58.250 85.070 ;
        RECT 58.920 84.900 59.090 85.070 ;
        RECT 59.280 84.900 59.450 85.070 ;
        RECT 59.640 84.900 59.810 85.070 ;
        RECT 61.230 84.910 61.400 85.080 ;
        RECT 61.670 84.910 61.840 85.080 ;
        RECT 62.080 84.910 62.250 85.080 ;
        RECT 62.510 84.910 62.680 85.080 ;
        RECT 62.950 84.910 63.120 85.080 ;
        RECT 63.360 84.910 63.530 85.080 ;
        RECT 65.350 84.900 65.520 85.070 ;
        RECT 65.710 84.900 65.880 85.070 ;
        RECT 66.070 84.900 66.240 85.070 ;
        RECT 66.430 84.900 66.600 85.070 ;
        RECT 67.950 84.910 68.120 85.080 ;
        RECT 68.390 84.910 68.560 85.080 ;
        RECT 68.800 84.910 68.970 85.080 ;
        RECT 69.230 84.910 69.400 85.080 ;
        RECT 69.670 84.910 69.840 85.080 ;
        RECT 70.080 84.910 70.250 85.080 ;
        RECT 72.120 84.900 72.290 85.070 ;
        RECT 72.480 84.900 72.650 85.070 ;
        RECT 72.840 84.900 73.010 85.070 ;
        RECT 73.200 84.900 73.370 85.070 ;
        RECT 74.620 84.900 74.790 85.070 ;
        RECT 75.060 84.900 75.230 85.070 ;
        RECT 75.500 84.900 75.670 85.070 ;
        RECT 75.910 84.900 76.080 85.070 ;
        RECT 76.900 84.900 77.070 85.070 ;
        RECT 77.490 84.900 77.660 85.070 ;
        RECT 79.010 84.900 79.180 85.070 ;
        RECT 79.370 84.900 79.540 85.070 ;
        RECT 80.380 84.900 80.550 85.070 ;
        RECT 80.820 84.900 80.990 85.070 ;
        RECT 81.260 84.900 81.430 85.070 ;
        RECT 81.670 84.900 81.840 85.070 ;
        RECT 82.200 84.900 82.370 85.070 ;
        RECT 82.560 84.900 82.730 85.070 ;
        RECT 84.220 84.900 84.390 85.070 ;
        RECT 84.580 84.900 84.750 85.070 ;
        RECT 84.940 84.900 85.110 85.070 ;
        RECT 85.300 84.900 85.470 85.070 ;
        RECT 85.660 84.900 85.830 85.070 ;
        RECT 86.140 84.900 86.310 85.070 ;
        RECT 86.580 84.900 86.750 85.070 ;
        RECT 87.020 84.900 87.190 85.070 ;
        RECT 87.430 84.900 87.600 85.070 ;
        RECT 87.960 84.900 88.130 85.070 ;
        RECT 88.320 84.900 88.490 85.070 ;
        RECT 88.680 84.900 88.850 85.070 ;
        RECT 89.520 84.900 89.690 85.070 ;
        RECT 89.880 84.900 90.050 85.070 ;
        RECT 90.240 84.900 90.410 85.070 ;
        RECT 91.080 84.900 91.250 85.070 ;
        RECT 91.440 84.900 91.610 85.070 ;
        RECT 91.800 84.900 91.970 85.070 ;
        RECT 92.860 84.900 93.030 85.070 ;
        RECT 93.300 84.900 93.470 85.070 ;
        RECT 93.740 84.900 93.910 85.070 ;
        RECT 94.150 84.900 94.320 85.070 ;
        RECT 94.680 84.900 94.850 85.070 ;
        RECT 95.040 84.900 95.210 85.070 ;
        RECT 95.400 84.900 95.570 85.070 ;
        RECT 96.240 84.900 96.410 85.070 ;
        RECT 96.600 84.900 96.770 85.070 ;
        RECT 96.960 84.900 97.130 85.070 ;
        RECT 97.800 84.900 97.970 85.070 ;
        RECT 98.160 84.900 98.330 85.070 ;
        RECT 98.520 84.900 98.690 85.070 ;
        RECT 99.580 84.900 99.750 85.070 ;
        RECT 100.020 84.900 100.190 85.070 ;
        RECT 100.460 84.900 100.630 85.070 ;
        RECT 100.870 84.900 101.040 85.070 ;
        RECT 101.400 84.900 101.570 85.070 ;
        RECT 101.760 84.900 101.930 85.070 ;
        RECT 102.940 84.900 103.110 85.070 ;
        RECT 103.380 84.900 103.550 85.070 ;
        RECT 103.820 84.900 103.990 85.070 ;
        RECT 104.230 84.900 104.400 85.070 ;
        RECT 105.710 84.900 105.880 85.070 ;
        RECT 106.070 84.900 106.240 85.070 ;
        RECT 106.430 84.900 106.600 85.070 ;
        RECT 107.350 84.900 107.520 85.070 ;
        RECT 107.710 84.900 107.880 85.070 ;
        RECT 112.310 84.900 112.480 85.070 ;
        RECT 112.670 84.900 112.840 85.070 ;
        RECT 113.030 84.900 113.200 85.070 ;
        RECT 116.280 84.900 116.450 85.070 ;
        RECT 116.640 84.900 116.810 85.070 ;
        RECT 117.000 84.900 117.170 85.070 ;
        RECT 118.890 84.900 119.060 85.070 ;
        RECT 119.250 84.900 119.420 85.070 ;
        RECT 119.610 84.900 119.780 85.070 ;
        RECT 121.230 84.910 121.400 85.080 ;
        RECT 121.670 84.910 121.840 85.080 ;
        RECT 122.080 84.910 122.250 85.080 ;
        RECT 122.510 84.910 122.680 85.080 ;
        RECT 122.950 84.910 123.120 85.080 ;
        RECT 123.360 84.910 123.530 85.080 ;
        RECT 125.070 84.910 125.240 85.080 ;
        RECT 125.510 84.910 125.680 85.080 ;
        RECT 125.920 84.910 126.090 85.080 ;
        RECT 126.350 84.910 126.520 85.080 ;
        RECT 126.790 84.910 126.960 85.080 ;
        RECT 127.200 84.910 127.370 85.080 ;
        RECT 128.910 84.910 129.080 85.080 ;
        RECT 129.350 84.910 129.520 85.080 ;
        RECT 129.760 84.910 129.930 85.080 ;
        RECT 130.190 84.910 130.360 85.080 ;
        RECT 130.630 84.910 130.800 85.080 ;
        RECT 131.040 84.910 131.210 85.080 ;
        RECT 132.750 84.910 132.920 85.080 ;
        RECT 133.190 84.910 133.360 85.080 ;
        RECT 133.600 84.910 133.770 85.080 ;
        RECT 134.030 84.910 134.200 85.080 ;
        RECT 134.470 84.910 134.640 85.080 ;
        RECT 134.880 84.910 135.050 85.080 ;
        RECT 136.590 84.910 136.760 85.080 ;
        RECT 137.030 84.910 137.200 85.080 ;
        RECT 137.440 84.910 137.610 85.080 ;
        RECT 137.870 84.910 138.040 85.080 ;
        RECT 138.310 84.910 138.480 85.080 ;
        RECT 138.720 84.910 138.890 85.080 ;
        RECT 139.900 84.900 140.070 85.070 ;
        RECT 140.340 84.900 140.510 85.070 ;
        RECT 140.780 84.900 140.950 85.070 ;
        RECT 141.190 84.900 141.360 85.070 ;
        RECT 5.920 77.240 6.090 77.420 ;
        RECT 6.400 77.240 6.570 77.420 ;
        RECT 6.880 77.240 7.050 77.420 ;
        RECT 7.360 77.240 7.530 77.420 ;
        RECT 7.840 77.240 8.010 77.420 ;
        RECT 8.320 77.240 8.490 77.420 ;
        RECT 8.800 77.240 8.970 77.420 ;
        RECT 9.280 77.240 9.450 77.420 ;
        RECT 9.760 77.240 9.930 77.420 ;
        RECT 10.240 77.240 10.410 77.420 ;
        RECT 10.720 77.240 10.890 77.420 ;
        RECT 11.200 77.240 11.370 77.420 ;
        RECT 11.680 77.240 11.850 77.420 ;
        RECT 12.160 77.240 12.330 77.420 ;
        RECT 12.640 77.240 12.810 77.420 ;
        RECT 13.120 77.240 13.290 77.420 ;
        RECT 13.600 77.240 13.770 77.420 ;
        RECT 14.080 77.240 14.250 77.420 ;
      LAYER li1 ;
        RECT 14.400 77.240 14.880 77.420 ;
      LAYER li1 ;
        RECT 15.040 77.240 15.210 77.420 ;
        RECT 15.520 77.240 15.690 77.420 ;
        RECT 16.000 77.240 16.170 77.420 ;
        RECT 16.480 77.240 16.650 77.420 ;
        RECT 16.960 77.240 17.130 77.420 ;
        RECT 17.440 77.240 17.610 77.420 ;
        RECT 17.920 77.240 18.090 77.420 ;
        RECT 18.400 77.240 18.570 77.420 ;
        RECT 18.880 77.240 19.050 77.420 ;
        RECT 19.360 77.240 19.530 77.420 ;
        RECT 19.840 77.240 20.010 77.420 ;
        RECT 20.320 77.240 20.490 77.420 ;
        RECT 20.800 77.240 20.970 77.420 ;
        RECT 21.280 77.240 21.450 77.420 ;
        RECT 21.760 77.240 21.930 77.420 ;
        RECT 22.240 77.240 22.410 77.420 ;
        RECT 22.720 77.240 22.890 77.420 ;
        RECT 23.200 77.240 23.370 77.420 ;
        RECT 23.680 77.240 23.850 77.420 ;
        RECT 24.160 77.240 24.330 77.420 ;
        RECT 24.640 77.240 24.810 77.420 ;
        RECT 25.120 77.240 25.290 77.420 ;
        RECT 25.600 77.240 25.770 77.420 ;
        RECT 26.080 77.240 26.250 77.420 ;
        RECT 26.560 77.240 26.730 77.420 ;
        RECT 27.040 77.240 27.210 77.420 ;
        RECT 27.520 77.240 27.690 77.420 ;
        RECT 28.000 77.240 28.170 77.420 ;
        RECT 28.480 77.240 28.650 77.420 ;
        RECT 28.960 77.240 29.130 77.420 ;
        RECT 29.440 77.240 29.610 77.420 ;
        RECT 29.920 77.240 30.090 77.420 ;
        RECT 30.400 77.240 30.570 77.420 ;
        RECT 30.880 77.240 31.050 77.420 ;
        RECT 31.360 77.240 31.530 77.420 ;
        RECT 31.840 77.240 32.010 77.420 ;
        RECT 32.320 77.240 32.490 77.420 ;
        RECT 32.800 77.240 32.970 77.420 ;
        RECT 33.280 77.240 33.450 77.420 ;
        RECT 33.760 77.240 33.930 77.420 ;
        RECT 34.240 77.240 34.410 77.420 ;
        RECT 34.720 77.240 34.890 77.420 ;
        RECT 35.200 77.240 35.370 77.420 ;
        RECT 35.680 77.240 35.850 77.420 ;
        RECT 36.160 77.240 36.330 77.420 ;
        RECT 36.640 77.240 36.810 77.420 ;
        RECT 37.120 77.240 37.290 77.420 ;
        RECT 37.600 77.240 37.770 77.420 ;
        RECT 38.080 77.240 38.250 77.420 ;
        RECT 38.560 77.240 38.730 77.420 ;
        RECT 39.040 77.240 39.210 77.420 ;
        RECT 39.520 77.240 39.690 77.420 ;
        RECT 40.000 77.240 40.170 77.420 ;
        RECT 40.480 77.240 40.650 77.420 ;
        RECT 40.960 77.240 41.130 77.420 ;
        RECT 41.440 77.240 41.610 77.420 ;
        RECT 41.920 77.240 42.090 77.420 ;
        RECT 42.400 77.240 42.570 77.420 ;
        RECT 42.880 77.240 43.050 77.420 ;
        RECT 43.360 77.240 43.530 77.420 ;
        RECT 43.840 77.240 44.010 77.420 ;
        RECT 44.320 77.240 44.490 77.420 ;
        RECT 44.800 77.240 44.970 77.420 ;
        RECT 45.280 77.240 45.450 77.420 ;
        RECT 45.760 77.240 45.930 77.420 ;
        RECT 46.240 77.240 46.410 77.420 ;
        RECT 46.720 77.240 46.890 77.420 ;
        RECT 47.200 77.240 47.370 77.420 ;
        RECT 47.680 77.240 47.850 77.420 ;
        RECT 48.160 77.240 48.330 77.420 ;
        RECT 48.640 77.240 48.810 77.420 ;
        RECT 49.120 77.240 49.290 77.420 ;
        RECT 49.600 77.240 49.770 77.420 ;
        RECT 50.080 77.240 50.250 77.420 ;
        RECT 50.560 77.240 50.730 77.420 ;
        RECT 51.040 77.240 51.210 77.420 ;
        RECT 51.520 77.240 51.690 77.420 ;
        RECT 52.000 77.240 52.170 77.420 ;
        RECT 52.480 77.240 52.650 77.420 ;
        RECT 52.960 77.240 53.130 77.420 ;
        RECT 53.440 77.240 53.610 77.420 ;
        RECT 53.920 77.240 54.090 77.420 ;
        RECT 54.400 77.240 54.570 77.420 ;
        RECT 54.880 77.240 55.050 77.420 ;
        RECT 55.360 77.240 55.530 77.420 ;
        RECT 55.840 77.240 56.010 77.420 ;
        RECT 56.320 77.240 56.490 77.420 ;
        RECT 56.800 77.240 56.970 77.420 ;
        RECT 57.280 77.240 57.450 77.420 ;
        RECT 57.760 77.240 57.930 77.420 ;
        RECT 58.240 77.240 58.410 77.420 ;
        RECT 58.720 77.240 58.890 77.420 ;
        RECT 59.200 77.240 59.370 77.420 ;
        RECT 59.680 77.240 59.850 77.420 ;
        RECT 60.160 77.240 60.330 77.420 ;
        RECT 60.640 77.240 60.810 77.420 ;
        RECT 61.120 77.240 61.290 77.420 ;
        RECT 61.600 77.240 61.770 77.420 ;
        RECT 62.080 77.240 62.250 77.420 ;
        RECT 62.560 77.240 62.730 77.420 ;
        RECT 63.040 77.240 63.210 77.420 ;
        RECT 63.520 77.240 63.690 77.420 ;
        RECT 64.000 77.240 64.170 77.420 ;
        RECT 64.480 77.240 64.650 77.420 ;
        RECT 64.960 77.240 65.130 77.420 ;
        RECT 65.440 77.240 65.610 77.420 ;
        RECT 65.920 77.240 66.090 77.420 ;
        RECT 66.400 77.240 66.570 77.420 ;
        RECT 66.880 77.240 67.050 77.420 ;
        RECT 67.360 77.240 67.530 77.420 ;
        RECT 67.840 77.240 68.010 77.420 ;
        RECT 68.320 77.240 68.490 77.420 ;
        RECT 68.800 77.240 68.970 77.420 ;
        RECT 69.280 77.240 69.450 77.420 ;
        RECT 69.760 77.240 69.930 77.420 ;
        RECT 70.240 77.240 70.410 77.420 ;
        RECT 70.720 77.240 70.890 77.420 ;
      LAYER li1 ;
        RECT 71.040 77.240 71.520 77.420 ;
      LAYER li1 ;
        RECT 71.680 77.240 71.850 77.420 ;
        RECT 72.160 77.240 72.330 77.420 ;
        RECT 72.640 77.240 72.810 77.420 ;
        RECT 73.120 77.240 73.290 77.420 ;
        RECT 73.600 77.240 73.770 77.420 ;
        RECT 74.080 77.240 74.250 77.420 ;
        RECT 74.560 77.240 74.730 77.420 ;
        RECT 75.040 77.240 75.210 77.420 ;
        RECT 75.520 77.240 75.690 77.420 ;
        RECT 76.000 77.240 76.170 77.420 ;
        RECT 76.480 77.240 76.650 77.420 ;
        RECT 76.960 77.240 77.130 77.420 ;
        RECT 77.440 77.240 77.610 77.420 ;
        RECT 77.920 77.240 78.090 77.420 ;
        RECT 78.400 77.240 78.570 77.420 ;
        RECT 78.880 77.240 79.050 77.420 ;
        RECT 79.360 77.240 79.530 77.420 ;
        RECT 79.840 77.240 80.010 77.420 ;
        RECT 80.320 77.240 80.490 77.420 ;
      LAYER li1 ;
        RECT 80.640 77.240 81.120 77.420 ;
      LAYER li1 ;
        RECT 81.280 77.240 81.450 77.420 ;
        RECT 81.760 77.240 81.930 77.420 ;
        RECT 82.240 77.240 82.410 77.420 ;
        RECT 82.720 77.240 82.890 77.420 ;
        RECT 83.200 77.240 83.370 77.420 ;
        RECT 83.680 77.240 83.850 77.420 ;
        RECT 84.160 77.240 84.330 77.420 ;
        RECT 84.640 77.240 84.810 77.420 ;
        RECT 85.120 77.240 85.290 77.420 ;
        RECT 85.600 77.240 85.770 77.420 ;
        RECT 86.080 77.240 86.250 77.420 ;
        RECT 86.560 77.240 86.730 77.420 ;
        RECT 87.040 77.240 87.210 77.420 ;
        RECT 87.520 77.240 87.690 77.420 ;
        RECT 88.000 77.240 88.170 77.420 ;
        RECT 88.480 77.240 88.650 77.420 ;
        RECT 88.960 77.240 89.130 77.420 ;
        RECT 89.440 77.240 89.610 77.420 ;
        RECT 89.920 77.240 90.090 77.420 ;
        RECT 90.400 77.240 90.570 77.420 ;
        RECT 90.880 77.240 91.050 77.420 ;
        RECT 91.360 77.240 91.530 77.420 ;
        RECT 91.840 77.240 92.010 77.420 ;
        RECT 92.320 77.240 92.490 77.420 ;
        RECT 92.800 77.240 92.970 77.420 ;
        RECT 93.280 77.240 93.450 77.420 ;
        RECT 93.760 77.240 93.930 77.420 ;
        RECT 94.240 77.240 94.410 77.420 ;
        RECT 94.720 77.240 94.890 77.420 ;
        RECT 95.200 77.240 95.370 77.420 ;
        RECT 95.680 77.240 95.850 77.420 ;
        RECT 96.160 77.240 96.330 77.420 ;
        RECT 96.640 77.240 96.810 77.420 ;
        RECT 97.120 77.240 97.290 77.420 ;
        RECT 97.600 77.240 97.770 77.420 ;
        RECT 98.080 77.240 98.250 77.420 ;
        RECT 98.560 77.240 98.730 77.420 ;
        RECT 99.040 77.240 99.210 77.420 ;
        RECT 99.520 77.240 99.690 77.420 ;
        RECT 100.000 77.240 100.170 77.420 ;
        RECT 100.480 77.240 100.650 77.420 ;
        RECT 100.960 77.240 101.130 77.420 ;
        RECT 101.440 77.240 101.610 77.420 ;
        RECT 101.920 77.240 102.090 77.420 ;
        RECT 102.400 77.240 102.570 77.420 ;
        RECT 102.880 77.240 103.050 77.420 ;
        RECT 103.360 77.240 103.530 77.420 ;
        RECT 103.840 77.240 104.010 77.420 ;
        RECT 104.320 77.240 104.490 77.420 ;
        RECT 104.800 77.240 104.970 77.420 ;
        RECT 105.280 77.240 105.450 77.420 ;
        RECT 105.760 77.240 105.930 77.420 ;
        RECT 106.240 77.240 106.410 77.420 ;
        RECT 106.720 77.240 106.890 77.420 ;
        RECT 107.200 77.240 107.370 77.420 ;
        RECT 107.680 77.240 107.850 77.420 ;
        RECT 108.160 77.240 108.330 77.420 ;
        RECT 108.640 77.240 108.810 77.420 ;
        RECT 109.120 77.240 109.290 77.420 ;
        RECT 109.600 77.240 109.770 77.420 ;
        RECT 110.080 77.240 110.250 77.420 ;
        RECT 110.560 77.240 110.730 77.420 ;
        RECT 111.040 77.240 111.210 77.420 ;
        RECT 111.520 77.240 111.690 77.420 ;
        RECT 112.000 77.240 112.170 77.420 ;
        RECT 112.480 77.240 112.650 77.420 ;
        RECT 112.960 77.240 113.130 77.420 ;
        RECT 113.440 77.240 113.610 77.420 ;
        RECT 113.920 77.240 114.090 77.420 ;
        RECT 114.400 77.240 114.570 77.420 ;
        RECT 114.880 77.240 115.050 77.420 ;
        RECT 115.360 77.240 115.530 77.420 ;
        RECT 115.840 77.240 116.010 77.420 ;
        RECT 116.320 77.240 116.490 77.420 ;
        RECT 116.800 77.240 116.970 77.420 ;
        RECT 117.280 77.240 117.450 77.420 ;
        RECT 117.760 77.240 117.930 77.420 ;
        RECT 118.240 77.240 118.410 77.420 ;
        RECT 118.720 77.240 118.890 77.420 ;
        RECT 119.200 77.240 119.370 77.420 ;
        RECT 119.680 77.240 119.850 77.420 ;
        RECT 120.160 77.240 120.330 77.420 ;
        RECT 120.640 77.240 120.810 77.420 ;
        RECT 121.120 77.240 121.290 77.420 ;
        RECT 121.600 77.240 121.770 77.420 ;
        RECT 122.080 77.240 122.250 77.420 ;
        RECT 122.560 77.240 122.730 77.420 ;
        RECT 123.040 77.240 123.210 77.420 ;
        RECT 123.520 77.240 123.690 77.420 ;
        RECT 124.000 77.240 124.170 77.420 ;
        RECT 124.480 77.240 124.650 77.420 ;
        RECT 124.960 77.240 125.130 77.420 ;
        RECT 125.440 77.240 125.610 77.420 ;
        RECT 125.920 77.240 126.090 77.420 ;
        RECT 126.400 77.240 126.570 77.420 ;
        RECT 126.880 77.240 127.050 77.420 ;
        RECT 127.360 77.240 127.530 77.420 ;
        RECT 127.840 77.240 128.010 77.420 ;
        RECT 128.320 77.240 128.490 77.420 ;
        RECT 128.800 77.240 128.970 77.420 ;
        RECT 129.280 77.240 129.450 77.420 ;
        RECT 129.760 77.240 129.930 77.420 ;
        RECT 130.240 77.240 130.410 77.420 ;
        RECT 130.720 77.240 130.890 77.420 ;
        RECT 131.200 77.240 131.370 77.420 ;
        RECT 131.680 77.240 131.850 77.420 ;
        RECT 132.160 77.240 132.330 77.420 ;
        RECT 132.640 77.240 132.810 77.420 ;
        RECT 133.120 77.240 133.290 77.420 ;
        RECT 133.600 77.240 133.770 77.420 ;
        RECT 134.080 77.240 134.250 77.420 ;
        RECT 134.560 77.240 134.730 77.420 ;
        RECT 135.040 77.240 135.210 77.420 ;
        RECT 135.520 77.240 135.690 77.420 ;
        RECT 136.000 77.240 136.170 77.420 ;
        RECT 136.480 77.240 136.650 77.420 ;
        RECT 136.960 77.240 137.130 77.420 ;
        RECT 137.440 77.240 137.610 77.420 ;
        RECT 137.920 77.240 138.090 77.420 ;
        RECT 138.400 77.240 138.570 77.420 ;
        RECT 138.880 77.240 139.050 77.420 ;
        RECT 139.360 77.240 139.530 77.420 ;
        RECT 139.840 77.240 140.010 77.420 ;
        RECT 140.320 77.240 140.490 77.420 ;
        RECT 140.800 77.240 140.970 77.420 ;
        RECT 141.280 77.240 141.450 77.420 ;
        RECT 141.760 77.240 141.930 77.420 ;
        RECT 6.510 76.770 6.680 76.940 ;
        RECT 6.950 76.770 7.120 76.940 ;
        RECT 7.360 76.770 7.530 76.940 ;
        RECT 7.790 76.770 7.960 76.940 ;
        RECT 8.230 76.770 8.400 76.940 ;
        RECT 8.640 76.770 8.810 76.940 ;
        RECT 10.350 76.770 10.520 76.940 ;
        RECT 10.790 76.770 10.960 76.940 ;
        RECT 11.200 76.770 11.370 76.940 ;
        RECT 11.630 76.770 11.800 76.940 ;
        RECT 12.070 76.770 12.240 76.940 ;
        RECT 12.480 76.770 12.650 76.940 ;
        RECT 14.190 76.770 14.360 76.940 ;
        RECT 14.630 76.770 14.800 76.940 ;
        RECT 15.040 76.770 15.210 76.940 ;
        RECT 15.470 76.770 15.640 76.940 ;
        RECT 15.910 76.770 16.080 76.940 ;
        RECT 16.320 76.770 16.490 76.940 ;
        RECT 17.830 76.760 18.000 76.930 ;
        RECT 18.190 76.760 18.360 76.930 ;
        RECT 18.550 76.760 18.720 76.930 ;
        RECT 18.910 76.760 19.080 76.930 ;
        RECT 19.900 76.760 20.070 76.930 ;
        RECT 20.340 76.760 20.510 76.930 ;
        RECT 20.780 76.760 20.950 76.930 ;
        RECT 21.190 76.760 21.360 76.930 ;
        RECT 22.150 76.760 22.320 76.930 ;
        RECT 22.510 76.760 22.680 76.930 ;
        RECT 22.870 76.760 23.040 76.930 ;
        RECT 23.230 76.760 23.400 76.930 ;
        RECT 24.220 76.760 24.390 76.930 ;
        RECT 24.660 76.760 24.830 76.930 ;
        RECT 25.100 76.760 25.270 76.930 ;
        RECT 25.510 76.760 25.680 76.930 ;
        RECT 26.040 76.760 26.210 76.930 ;
        RECT 26.400 76.760 26.570 76.930 ;
        RECT 26.760 76.760 26.930 76.930 ;
        RECT 27.600 76.760 27.770 76.930 ;
        RECT 27.960 76.760 28.130 76.930 ;
        RECT 28.320 76.760 28.490 76.930 ;
        RECT 29.160 76.760 29.330 76.930 ;
        RECT 29.520 76.760 29.690 76.930 ;
        RECT 29.880 76.760 30.050 76.930 ;
        RECT 30.940 76.760 31.110 76.930 ;
        RECT 31.380 76.760 31.550 76.930 ;
        RECT 31.820 76.760 31.990 76.930 ;
        RECT 32.230 76.760 32.400 76.930 ;
        RECT 32.760 76.760 32.930 76.930 ;
        RECT 33.120 76.760 33.290 76.930 ;
        RECT 33.480 76.760 33.650 76.930 ;
        RECT 34.320 76.760 34.490 76.930 ;
        RECT 34.680 76.760 34.850 76.930 ;
        RECT 35.040 76.760 35.210 76.930 ;
        RECT 35.880 76.760 36.050 76.930 ;
        RECT 36.240 76.760 36.410 76.930 ;
        RECT 36.600 76.760 36.770 76.930 ;
        RECT 37.660 76.760 37.830 76.930 ;
        RECT 38.100 76.760 38.270 76.930 ;
        RECT 38.540 76.760 38.710 76.930 ;
        RECT 38.950 76.760 39.120 76.930 ;
        RECT 39.480 76.760 39.650 76.930 ;
        RECT 39.840 76.760 40.010 76.930 ;
        RECT 40.200 76.760 40.370 76.930 ;
        RECT 41.040 76.760 41.210 76.930 ;
        RECT 41.400 76.760 41.570 76.930 ;
        RECT 41.760 76.760 41.930 76.930 ;
        RECT 42.600 76.760 42.770 76.930 ;
        RECT 42.960 76.760 43.130 76.930 ;
        RECT 43.320 76.760 43.490 76.930 ;
        RECT 44.380 76.760 44.550 76.930 ;
        RECT 44.820 76.760 44.990 76.930 ;
        RECT 45.260 76.760 45.430 76.930 ;
        RECT 45.670 76.760 45.840 76.930 ;
        RECT 47.640 76.760 47.810 76.930 ;
        RECT 48.000 76.760 48.170 76.930 ;
        RECT 48.360 76.760 48.530 76.930 ;
        RECT 49.200 76.760 49.370 76.930 ;
        RECT 49.560 76.760 49.730 76.930 ;
        RECT 49.920 76.760 50.090 76.930 ;
        RECT 50.760 76.760 50.930 76.930 ;
        RECT 51.120 76.760 51.290 76.930 ;
        RECT 51.480 76.760 51.650 76.930 ;
        RECT 52.540 76.760 52.710 76.930 ;
        RECT 52.980 76.760 53.150 76.930 ;
        RECT 53.420 76.760 53.590 76.930 ;
        RECT 53.830 76.760 54.000 76.930 ;
        RECT 54.840 76.760 55.010 76.930 ;
        RECT 55.200 76.760 55.370 76.930 ;
        RECT 55.560 76.760 55.730 76.930 ;
        RECT 55.920 76.760 56.090 76.930 ;
        RECT 56.280 76.760 56.450 76.930 ;
        RECT 57.330 76.760 57.500 76.930 ;
        RECT 57.690 76.760 57.860 76.930 ;
        RECT 58.050 76.760 58.220 76.930 ;
        RECT 58.410 76.760 58.580 76.930 ;
        RECT 58.770 76.760 58.940 76.930 ;
        RECT 59.740 76.760 59.910 76.930 ;
        RECT 60.180 76.760 60.350 76.930 ;
        RECT 60.620 76.760 60.790 76.930 ;
        RECT 61.030 76.760 61.200 76.930 ;
        RECT 62.030 76.760 62.200 76.930 ;
        RECT 62.390 76.760 62.560 76.930 ;
        RECT 62.750 76.760 62.920 76.930 ;
        RECT 63.670 76.760 63.840 76.930 ;
        RECT 64.030 76.760 64.200 76.930 ;
        RECT 68.630 76.760 68.800 76.930 ;
        RECT 68.990 76.760 69.160 76.930 ;
        RECT 69.350 76.760 69.520 76.930 ;
        RECT 72.600 76.760 72.770 76.930 ;
        RECT 72.960 76.760 73.130 76.930 ;
        RECT 73.320 76.760 73.490 76.930 ;
        RECT 75.210 76.760 75.380 76.930 ;
        RECT 75.570 76.760 75.740 76.930 ;
        RECT 75.930 76.760 76.100 76.930 ;
        RECT 77.020 76.760 77.190 76.930 ;
        RECT 77.460 76.760 77.630 76.930 ;
        RECT 77.900 76.760 78.070 76.930 ;
        RECT 78.310 76.760 78.480 76.930 ;
        RECT 79.320 76.760 79.490 76.930 ;
        RECT 79.680 76.760 79.850 76.930 ;
        RECT 80.860 76.760 81.030 76.930 ;
        RECT 81.300 76.760 81.470 76.930 ;
        RECT 81.740 76.760 81.910 76.930 ;
        RECT 82.150 76.760 82.320 76.930 ;
        RECT 83.120 76.760 83.290 76.930 ;
        RECT 83.480 76.760 83.650 76.930 ;
        RECT 83.840 76.760 84.010 76.930 ;
        RECT 86.480 76.760 86.650 76.930 ;
        RECT 86.840 76.760 87.010 76.930 ;
        RECT 87.200 76.760 87.370 76.930 ;
        RECT 87.560 76.760 87.730 76.930 ;
        RECT 88.060 76.760 88.230 76.930 ;
        RECT 88.500 76.760 88.670 76.930 ;
        RECT 88.940 76.760 89.110 76.930 ;
        RECT 89.350 76.760 89.520 76.930 ;
        RECT 90.360 76.760 90.530 76.930 ;
        RECT 90.870 76.760 91.040 76.930 ;
        RECT 92.550 76.760 92.720 76.930 ;
        RECT 92.910 76.760 93.080 76.930 ;
        RECT 93.270 76.760 93.440 76.930 ;
        RECT 94.300 76.760 94.470 76.930 ;
        RECT 94.740 76.760 94.910 76.930 ;
        RECT 95.180 76.760 95.350 76.930 ;
        RECT 95.590 76.760 95.760 76.930 ;
        RECT 96.640 76.760 96.810 76.930 ;
        RECT 97.000 76.760 97.170 76.930 ;
        RECT 97.360 76.760 97.530 76.930 ;
        RECT 99.580 76.760 99.750 76.930 ;
        RECT 100.020 76.760 100.190 76.930 ;
        RECT 100.460 76.760 100.630 76.930 ;
        RECT 100.870 76.760 101.040 76.930 ;
        RECT 101.880 76.760 102.050 76.930 ;
        RECT 102.240 76.760 102.410 76.930 ;
        RECT 102.600 76.760 102.770 76.930 ;
        RECT 102.960 76.760 103.130 76.930 ;
        RECT 103.320 76.760 103.490 76.930 ;
        RECT 104.370 76.760 104.540 76.930 ;
        RECT 104.730 76.760 104.900 76.930 ;
        RECT 105.090 76.760 105.260 76.930 ;
        RECT 105.450 76.760 105.620 76.930 ;
        RECT 105.810 76.760 105.980 76.930 ;
        RECT 106.780 76.760 106.950 76.930 ;
        RECT 107.220 76.760 107.390 76.930 ;
        RECT 107.660 76.760 107.830 76.930 ;
        RECT 108.070 76.760 108.240 76.930 ;
        RECT 109.560 76.760 109.730 76.930 ;
        RECT 109.920 76.760 110.090 76.930 ;
        RECT 110.280 76.760 110.450 76.930 ;
        RECT 110.640 76.760 110.810 76.930 ;
        RECT 112.060 76.760 112.230 76.930 ;
        RECT 112.500 76.760 112.670 76.930 ;
        RECT 112.940 76.760 113.110 76.930 ;
        RECT 113.350 76.760 113.520 76.930 ;
        RECT 114.350 76.760 114.520 76.930 ;
        RECT 114.710 76.760 114.880 76.930 ;
        RECT 115.070 76.760 115.240 76.930 ;
        RECT 115.990 76.760 116.160 76.930 ;
        RECT 116.350 76.760 116.520 76.930 ;
        RECT 120.950 76.760 121.120 76.930 ;
        RECT 121.310 76.760 121.480 76.930 ;
        RECT 121.670 76.760 121.840 76.930 ;
        RECT 124.920 76.760 125.090 76.930 ;
        RECT 125.280 76.760 125.450 76.930 ;
        RECT 125.640 76.760 125.810 76.930 ;
        RECT 127.530 76.760 127.700 76.930 ;
        RECT 127.890 76.760 128.060 76.930 ;
        RECT 128.250 76.760 128.420 76.930 ;
        RECT 129.870 76.770 130.040 76.940 ;
        RECT 130.310 76.770 130.480 76.940 ;
        RECT 130.720 76.770 130.890 76.940 ;
        RECT 131.150 76.770 131.320 76.940 ;
        RECT 131.590 76.770 131.760 76.940 ;
        RECT 132.000 76.770 132.170 76.940 ;
        RECT 136.000 76.760 136.170 76.930 ;
        RECT 136.360 76.760 136.530 76.930 ;
        RECT 137.550 76.770 137.720 76.940 ;
        RECT 137.990 76.770 138.160 76.940 ;
        RECT 138.400 76.770 138.570 76.940 ;
        RECT 138.830 76.770 139.000 76.940 ;
        RECT 139.270 76.770 139.440 76.940 ;
        RECT 139.680 76.770 139.850 76.940 ;
        RECT 5.920 69.100 6.090 69.280 ;
        RECT 6.400 69.100 6.570 69.280 ;
        RECT 6.880 69.100 7.050 69.280 ;
        RECT 7.360 69.100 7.530 69.280 ;
        RECT 7.840 69.100 8.010 69.280 ;
        RECT 8.320 69.100 8.490 69.280 ;
        RECT 8.800 69.100 8.970 69.280 ;
        RECT 9.280 69.100 9.450 69.280 ;
        RECT 9.760 69.100 9.930 69.280 ;
        RECT 10.240 69.100 10.410 69.280 ;
        RECT 10.720 69.100 10.890 69.280 ;
        RECT 11.200 69.100 11.370 69.280 ;
        RECT 11.680 69.100 11.850 69.280 ;
        RECT 12.160 69.100 12.330 69.280 ;
        RECT 12.640 69.100 12.810 69.280 ;
        RECT 13.120 69.100 13.290 69.280 ;
        RECT 13.600 69.100 13.770 69.280 ;
        RECT 14.080 69.100 14.250 69.280 ;
        RECT 14.560 69.100 14.730 69.280 ;
        RECT 15.040 69.100 15.210 69.280 ;
        RECT 15.520 69.100 15.690 69.280 ;
        RECT 16.000 69.100 16.170 69.280 ;
        RECT 16.480 69.100 16.650 69.280 ;
        RECT 16.960 69.100 17.130 69.280 ;
        RECT 17.440 69.100 17.610 69.280 ;
        RECT 17.920 69.100 18.090 69.280 ;
        RECT 18.400 69.100 18.570 69.280 ;
        RECT 18.880 69.100 19.050 69.280 ;
        RECT 19.360 69.100 19.530 69.280 ;
        RECT 19.840 69.100 20.010 69.280 ;
        RECT 20.320 69.100 20.490 69.280 ;
        RECT 20.800 69.100 20.970 69.280 ;
        RECT 21.280 69.100 21.450 69.280 ;
        RECT 21.760 69.100 21.930 69.280 ;
        RECT 22.240 69.100 22.410 69.280 ;
        RECT 22.720 69.100 22.890 69.280 ;
        RECT 23.200 69.100 23.370 69.280 ;
        RECT 23.680 69.100 23.850 69.280 ;
        RECT 24.160 69.100 24.330 69.280 ;
        RECT 24.640 69.100 24.810 69.280 ;
        RECT 25.120 69.100 25.290 69.280 ;
        RECT 25.600 69.100 25.770 69.280 ;
        RECT 26.080 69.100 26.250 69.280 ;
        RECT 26.560 69.100 26.730 69.280 ;
        RECT 27.040 69.100 27.210 69.280 ;
        RECT 27.520 69.100 27.690 69.280 ;
        RECT 28.000 69.100 28.170 69.280 ;
        RECT 28.480 69.100 28.650 69.280 ;
        RECT 28.960 69.100 29.130 69.280 ;
        RECT 29.440 69.100 29.610 69.280 ;
        RECT 29.920 69.100 30.090 69.280 ;
        RECT 30.400 69.100 30.570 69.280 ;
        RECT 30.880 69.100 31.050 69.280 ;
        RECT 31.360 69.100 31.530 69.280 ;
        RECT 31.840 69.100 32.010 69.280 ;
        RECT 32.320 69.100 32.490 69.280 ;
        RECT 32.800 69.100 32.970 69.280 ;
        RECT 33.280 69.100 33.450 69.280 ;
        RECT 33.760 69.100 33.930 69.280 ;
        RECT 34.240 69.100 34.410 69.280 ;
        RECT 34.720 69.100 34.890 69.280 ;
        RECT 35.200 69.100 35.370 69.280 ;
        RECT 35.680 69.100 35.850 69.280 ;
        RECT 36.160 69.100 36.330 69.280 ;
        RECT 36.640 69.100 36.810 69.280 ;
        RECT 37.120 69.100 37.290 69.280 ;
        RECT 37.600 69.100 37.770 69.280 ;
        RECT 38.080 69.100 38.250 69.280 ;
        RECT 38.560 69.100 38.730 69.280 ;
        RECT 39.040 69.100 39.210 69.280 ;
        RECT 39.520 69.100 39.690 69.280 ;
        RECT 40.000 69.100 40.170 69.280 ;
        RECT 40.480 69.100 40.650 69.280 ;
        RECT 40.960 69.100 41.130 69.280 ;
        RECT 41.440 69.100 41.610 69.280 ;
        RECT 41.920 69.100 42.090 69.280 ;
        RECT 42.400 69.100 42.570 69.280 ;
        RECT 42.880 69.100 43.050 69.280 ;
        RECT 43.360 69.100 43.530 69.280 ;
        RECT 43.840 69.100 44.010 69.280 ;
        RECT 44.320 69.100 44.490 69.280 ;
        RECT 44.800 69.100 44.970 69.280 ;
        RECT 45.280 69.100 45.450 69.280 ;
        RECT 45.760 69.100 45.930 69.280 ;
        RECT 46.240 69.100 46.410 69.280 ;
        RECT 46.720 69.100 46.890 69.280 ;
        RECT 47.200 69.100 47.370 69.280 ;
      LAYER li1 ;
        RECT 47.520 69.100 48.000 69.280 ;
      LAYER li1 ;
        RECT 48.160 69.100 48.330 69.280 ;
        RECT 48.640 69.100 48.810 69.280 ;
        RECT 49.120 69.100 49.290 69.280 ;
        RECT 49.600 69.100 49.770 69.280 ;
        RECT 50.080 69.100 50.250 69.280 ;
        RECT 50.560 69.100 50.730 69.280 ;
        RECT 51.040 69.100 51.210 69.280 ;
        RECT 51.520 69.100 51.690 69.280 ;
        RECT 52.000 69.100 52.170 69.280 ;
        RECT 52.480 69.100 52.650 69.280 ;
        RECT 52.960 69.100 53.130 69.280 ;
        RECT 53.440 69.100 53.610 69.280 ;
        RECT 53.920 69.100 54.090 69.280 ;
        RECT 54.400 69.100 54.570 69.280 ;
        RECT 54.880 69.100 55.050 69.280 ;
        RECT 55.360 69.100 55.530 69.280 ;
        RECT 55.840 69.100 56.010 69.280 ;
        RECT 56.320 69.100 56.490 69.280 ;
        RECT 56.800 69.100 56.970 69.280 ;
        RECT 57.280 69.100 57.450 69.280 ;
        RECT 57.760 69.100 57.930 69.280 ;
        RECT 58.240 69.100 58.410 69.280 ;
        RECT 58.720 69.100 58.890 69.280 ;
      LAYER li1 ;
        RECT 59.040 69.100 59.520 69.280 ;
      LAYER li1 ;
        RECT 59.680 69.100 59.850 69.280 ;
        RECT 60.160 69.100 60.330 69.280 ;
        RECT 60.640 69.100 60.810 69.280 ;
        RECT 61.120 69.100 61.290 69.280 ;
        RECT 61.600 69.100 61.770 69.280 ;
        RECT 62.080 69.100 62.250 69.280 ;
        RECT 62.560 69.100 62.730 69.280 ;
        RECT 63.040 69.100 63.210 69.280 ;
        RECT 63.520 69.100 63.690 69.280 ;
        RECT 64.000 69.100 64.170 69.280 ;
        RECT 64.480 69.100 64.650 69.280 ;
        RECT 64.960 69.100 65.130 69.280 ;
        RECT 65.440 69.100 65.610 69.280 ;
        RECT 65.920 69.100 66.090 69.280 ;
        RECT 66.400 69.100 66.570 69.280 ;
        RECT 66.880 69.100 67.050 69.280 ;
        RECT 67.360 69.100 67.530 69.280 ;
        RECT 67.840 69.100 68.010 69.280 ;
        RECT 68.320 69.100 68.490 69.280 ;
        RECT 68.800 69.100 68.970 69.280 ;
        RECT 69.280 69.100 69.450 69.280 ;
        RECT 69.760 69.100 69.930 69.280 ;
        RECT 70.240 69.100 70.410 69.280 ;
        RECT 70.720 69.100 70.890 69.280 ;
        RECT 71.200 69.100 71.370 69.280 ;
        RECT 71.680 69.100 71.850 69.280 ;
        RECT 72.160 69.100 72.330 69.280 ;
        RECT 72.640 69.100 72.810 69.280 ;
        RECT 73.120 69.100 73.290 69.280 ;
        RECT 73.600 69.100 73.770 69.280 ;
        RECT 74.080 69.100 74.250 69.280 ;
        RECT 74.560 69.100 74.730 69.280 ;
        RECT 75.040 69.100 75.210 69.280 ;
        RECT 75.520 69.100 75.690 69.280 ;
        RECT 76.000 69.100 76.170 69.280 ;
      LAYER li1 ;
        RECT 76.320 69.100 76.800 69.280 ;
      LAYER li1 ;
        RECT 76.960 69.100 77.130 69.280 ;
        RECT 77.440 69.100 77.610 69.280 ;
        RECT 77.920 69.100 78.090 69.280 ;
        RECT 78.400 69.100 78.570 69.280 ;
        RECT 78.880 69.100 79.050 69.280 ;
        RECT 79.360 69.100 79.530 69.280 ;
        RECT 79.840 69.100 80.010 69.280 ;
        RECT 80.320 69.100 80.490 69.280 ;
        RECT 80.800 69.100 80.970 69.280 ;
        RECT 81.280 69.100 81.450 69.280 ;
        RECT 81.760 69.100 81.930 69.280 ;
        RECT 82.240 69.100 82.410 69.280 ;
        RECT 82.720 69.100 82.890 69.280 ;
        RECT 83.200 69.100 83.370 69.280 ;
        RECT 83.680 69.100 83.850 69.280 ;
        RECT 84.160 69.100 84.330 69.280 ;
        RECT 84.640 69.100 84.810 69.280 ;
        RECT 85.120 69.100 85.290 69.280 ;
        RECT 85.600 69.100 85.770 69.280 ;
        RECT 86.080 69.100 86.250 69.280 ;
        RECT 86.560 69.100 86.730 69.280 ;
        RECT 87.040 69.100 87.210 69.280 ;
        RECT 87.520 69.100 87.690 69.280 ;
        RECT 88.000 69.100 88.170 69.280 ;
        RECT 88.480 69.100 88.650 69.280 ;
        RECT 88.960 69.100 89.130 69.280 ;
        RECT 89.440 69.100 89.610 69.280 ;
        RECT 89.920 69.100 90.090 69.280 ;
        RECT 90.400 69.100 90.570 69.280 ;
        RECT 90.880 69.100 91.050 69.280 ;
        RECT 91.360 69.100 91.530 69.280 ;
        RECT 91.840 69.100 92.010 69.280 ;
        RECT 92.320 69.100 92.490 69.280 ;
        RECT 92.800 69.100 92.970 69.280 ;
        RECT 93.280 69.100 93.450 69.280 ;
        RECT 93.760 69.100 93.930 69.280 ;
        RECT 94.240 69.100 94.410 69.280 ;
        RECT 94.720 69.100 94.890 69.280 ;
        RECT 95.200 69.100 95.370 69.280 ;
        RECT 95.680 69.100 95.850 69.280 ;
        RECT 96.160 69.100 96.330 69.280 ;
        RECT 96.640 69.100 96.810 69.280 ;
        RECT 97.120 69.100 97.290 69.280 ;
        RECT 97.600 69.100 97.770 69.280 ;
        RECT 98.080 69.100 98.250 69.280 ;
        RECT 98.560 69.100 98.730 69.280 ;
        RECT 99.040 69.100 99.210 69.280 ;
        RECT 99.520 69.100 99.690 69.280 ;
        RECT 100.000 69.100 100.170 69.280 ;
        RECT 100.480 69.100 100.650 69.280 ;
        RECT 100.960 69.100 101.130 69.280 ;
        RECT 101.440 69.100 101.610 69.280 ;
        RECT 101.920 69.100 102.090 69.280 ;
        RECT 102.400 69.100 102.570 69.280 ;
        RECT 102.880 69.100 103.050 69.280 ;
        RECT 103.360 69.100 103.530 69.280 ;
        RECT 103.840 69.100 104.010 69.280 ;
        RECT 104.320 69.100 104.490 69.280 ;
        RECT 104.800 69.100 104.970 69.280 ;
        RECT 105.280 69.100 105.450 69.280 ;
        RECT 105.760 69.100 105.930 69.280 ;
        RECT 106.240 69.100 106.410 69.280 ;
        RECT 106.720 69.100 106.890 69.280 ;
        RECT 107.200 69.100 107.370 69.280 ;
        RECT 107.680 69.100 107.850 69.280 ;
        RECT 108.160 69.100 108.330 69.280 ;
        RECT 108.640 69.100 108.810 69.280 ;
        RECT 109.120 69.100 109.290 69.280 ;
        RECT 109.600 69.100 109.770 69.280 ;
        RECT 110.080 69.100 110.250 69.280 ;
        RECT 110.560 69.100 110.730 69.280 ;
        RECT 111.040 69.100 111.210 69.280 ;
        RECT 111.520 69.100 111.690 69.280 ;
        RECT 112.000 69.100 112.170 69.280 ;
        RECT 112.480 69.100 112.650 69.280 ;
        RECT 112.960 69.100 113.130 69.280 ;
        RECT 113.440 69.100 113.610 69.280 ;
        RECT 113.920 69.100 114.090 69.280 ;
        RECT 114.400 69.100 114.570 69.280 ;
        RECT 114.880 69.100 115.050 69.280 ;
        RECT 115.360 69.100 115.530 69.280 ;
        RECT 115.840 69.100 116.010 69.280 ;
        RECT 116.320 69.100 116.490 69.280 ;
        RECT 116.800 69.100 116.970 69.280 ;
        RECT 117.280 69.100 117.450 69.280 ;
        RECT 117.760 69.100 117.930 69.280 ;
        RECT 118.240 69.100 118.410 69.280 ;
        RECT 118.720 69.100 118.890 69.280 ;
        RECT 119.200 69.100 119.370 69.280 ;
        RECT 119.680 69.100 119.850 69.280 ;
        RECT 120.160 69.100 120.330 69.280 ;
        RECT 120.640 69.100 120.810 69.280 ;
        RECT 121.120 69.100 121.290 69.280 ;
        RECT 121.600 69.100 121.770 69.280 ;
        RECT 122.080 69.100 122.250 69.280 ;
        RECT 122.560 69.100 122.730 69.280 ;
        RECT 123.040 69.100 123.210 69.280 ;
        RECT 123.520 69.100 123.690 69.280 ;
        RECT 124.000 69.100 124.170 69.280 ;
        RECT 124.480 69.100 124.650 69.280 ;
        RECT 124.960 69.100 125.130 69.280 ;
        RECT 125.440 69.100 125.610 69.280 ;
        RECT 125.920 69.100 126.090 69.280 ;
        RECT 126.400 69.100 126.570 69.280 ;
        RECT 126.880 69.100 127.050 69.280 ;
        RECT 127.360 69.100 127.530 69.280 ;
        RECT 127.840 69.100 128.010 69.280 ;
        RECT 128.320 69.100 128.490 69.280 ;
        RECT 128.800 69.100 128.970 69.280 ;
        RECT 129.280 69.100 129.450 69.280 ;
        RECT 129.760 69.100 129.930 69.280 ;
        RECT 130.240 69.100 130.410 69.280 ;
        RECT 130.720 69.100 130.890 69.280 ;
        RECT 131.200 69.100 131.370 69.280 ;
        RECT 131.680 69.100 131.850 69.280 ;
        RECT 132.160 69.100 132.330 69.280 ;
        RECT 132.640 69.100 132.810 69.280 ;
        RECT 133.120 69.100 133.290 69.280 ;
        RECT 133.600 69.100 133.770 69.280 ;
        RECT 134.080 69.100 134.250 69.280 ;
        RECT 134.560 69.100 134.730 69.280 ;
        RECT 135.040 69.100 135.210 69.280 ;
        RECT 135.520 69.100 135.690 69.280 ;
        RECT 136.000 69.100 136.170 69.280 ;
        RECT 136.480 69.100 136.650 69.280 ;
        RECT 136.960 69.100 137.130 69.280 ;
        RECT 137.440 69.100 137.610 69.280 ;
        RECT 137.920 69.100 138.090 69.280 ;
        RECT 138.400 69.100 138.570 69.280 ;
        RECT 138.880 69.100 139.050 69.280 ;
        RECT 139.360 69.100 139.530 69.280 ;
        RECT 139.840 69.100 140.010 69.280 ;
        RECT 140.320 69.100 140.490 69.280 ;
        RECT 140.800 69.100 140.970 69.280 ;
        RECT 141.280 69.100 141.450 69.280 ;
        RECT 141.760 69.100 141.930 69.280 ;
        RECT 5.980 68.620 6.150 68.790 ;
        RECT 6.420 68.620 6.590 68.790 ;
        RECT 6.860 68.620 7.030 68.790 ;
        RECT 7.270 68.620 7.440 68.790 ;
        RECT 9.670 68.620 9.840 68.790 ;
        RECT 10.030 68.620 10.200 68.790 ;
        RECT 10.390 68.620 10.560 68.790 ;
        RECT 10.750 68.620 10.920 68.790 ;
        RECT 11.740 68.620 11.910 68.790 ;
        RECT 12.180 68.620 12.350 68.790 ;
        RECT 12.620 68.620 12.790 68.790 ;
        RECT 13.030 68.620 13.200 68.790 ;
        RECT 13.550 68.620 13.720 68.790 ;
        RECT 13.910 68.620 14.080 68.790 ;
        RECT 14.270 68.620 14.440 68.790 ;
        RECT 15.190 68.620 15.360 68.790 ;
        RECT 15.550 68.620 15.720 68.790 ;
        RECT 16.060 68.620 16.230 68.790 ;
        RECT 16.500 68.620 16.670 68.790 ;
        RECT 16.940 68.620 17.110 68.790 ;
        RECT 17.350 68.620 17.520 68.790 ;
        RECT 17.880 68.620 18.050 68.790 ;
        RECT 18.240 68.620 18.410 68.790 ;
        RECT 18.600 68.620 18.770 68.790 ;
        RECT 18.960 68.620 19.130 68.790 ;
        RECT 20.380 68.620 20.550 68.790 ;
        RECT 20.820 68.620 20.990 68.790 ;
        RECT 21.260 68.620 21.430 68.790 ;
        RECT 21.670 68.620 21.840 68.790 ;
        RECT 22.200 68.620 22.370 68.790 ;
        RECT 22.560 68.620 22.730 68.790 ;
        RECT 22.920 68.620 23.090 68.790 ;
        RECT 23.760 68.620 23.930 68.790 ;
        RECT 24.120 68.620 24.290 68.790 ;
        RECT 24.480 68.620 24.650 68.790 ;
        RECT 25.320 68.620 25.490 68.790 ;
        RECT 25.680 68.620 25.850 68.790 ;
        RECT 26.040 68.620 26.210 68.790 ;
        RECT 27.100 68.620 27.270 68.790 ;
        RECT 27.540 68.620 27.710 68.790 ;
        RECT 27.980 68.620 28.150 68.790 ;
        RECT 28.390 68.620 28.560 68.790 ;
        RECT 28.920 68.620 29.090 68.790 ;
        RECT 29.280 68.620 29.450 68.790 ;
        RECT 29.640 68.620 29.810 68.790 ;
        RECT 30.480 68.620 30.650 68.790 ;
        RECT 30.840 68.620 31.010 68.790 ;
        RECT 31.200 68.620 31.370 68.790 ;
        RECT 32.040 68.620 32.210 68.790 ;
        RECT 32.400 68.620 32.570 68.790 ;
        RECT 32.760 68.620 32.930 68.790 ;
        RECT 33.820 68.620 33.990 68.790 ;
        RECT 34.260 68.620 34.430 68.790 ;
        RECT 34.700 68.620 34.870 68.790 ;
        RECT 35.110 68.620 35.280 68.790 ;
        RECT 35.640 68.620 35.810 68.790 ;
        RECT 36.000 68.620 36.170 68.790 ;
        RECT 37.180 68.620 37.350 68.790 ;
        RECT 37.620 68.620 37.790 68.790 ;
        RECT 38.060 68.620 38.230 68.790 ;
        RECT 38.470 68.620 38.640 68.790 ;
        RECT 39.000 68.620 39.170 68.790 ;
        RECT 39.360 68.620 39.530 68.790 ;
        RECT 39.720 68.620 39.890 68.790 ;
        RECT 40.560 68.620 40.730 68.790 ;
        RECT 40.920 68.620 41.090 68.790 ;
        RECT 41.280 68.620 41.450 68.790 ;
        RECT 42.120 68.620 42.290 68.790 ;
        RECT 42.480 68.620 42.650 68.790 ;
        RECT 42.840 68.620 43.010 68.790 ;
        RECT 44.430 68.630 44.600 68.800 ;
        RECT 44.870 68.630 45.040 68.800 ;
        RECT 45.280 68.630 45.450 68.800 ;
        RECT 45.710 68.630 45.880 68.800 ;
        RECT 46.150 68.630 46.320 68.800 ;
        RECT 46.560 68.630 46.730 68.800 ;
        RECT 48.120 68.620 48.290 68.790 ;
        RECT 48.480 68.620 48.650 68.790 ;
        RECT 48.840 68.620 49.010 68.790 ;
        RECT 49.680 68.620 49.850 68.790 ;
        RECT 50.040 68.620 50.210 68.790 ;
        RECT 50.400 68.620 50.570 68.790 ;
        RECT 51.240 68.620 51.410 68.790 ;
        RECT 51.600 68.620 51.770 68.790 ;
        RECT 51.960 68.620 52.130 68.790 ;
        RECT 53.550 68.630 53.720 68.800 ;
        RECT 53.990 68.630 54.160 68.800 ;
        RECT 54.400 68.630 54.570 68.800 ;
        RECT 54.830 68.630 55.000 68.800 ;
        RECT 55.270 68.630 55.440 68.800 ;
        RECT 55.680 68.630 55.850 68.800 ;
        RECT 57.720 68.620 57.890 68.790 ;
        RECT 58.080 68.620 58.250 68.790 ;
        RECT 58.440 68.620 58.610 68.790 ;
        RECT 59.280 68.620 59.450 68.790 ;
        RECT 59.640 68.620 59.810 68.790 ;
        RECT 60.000 68.620 60.170 68.790 ;
        RECT 60.840 68.620 61.010 68.790 ;
        RECT 61.200 68.620 61.370 68.790 ;
        RECT 61.560 68.620 61.730 68.790 ;
        RECT 62.620 68.620 62.790 68.790 ;
        RECT 63.060 68.620 63.230 68.790 ;
        RECT 63.500 68.620 63.670 68.790 ;
        RECT 63.910 68.620 64.080 68.790 ;
        RECT 64.440 68.620 64.610 68.790 ;
        RECT 64.800 68.620 64.970 68.790 ;
        RECT 65.160 68.620 65.330 68.790 ;
        RECT 66.000 68.620 66.170 68.790 ;
        RECT 66.360 68.620 66.530 68.790 ;
        RECT 66.720 68.620 66.890 68.790 ;
        RECT 67.560 68.620 67.730 68.790 ;
        RECT 67.920 68.620 68.090 68.790 ;
        RECT 68.280 68.620 68.450 68.790 ;
        RECT 69.340 68.620 69.510 68.790 ;
        RECT 69.780 68.620 69.950 68.790 ;
        RECT 70.220 68.620 70.390 68.790 ;
        RECT 70.630 68.620 70.800 68.790 ;
        RECT 71.160 68.620 71.330 68.790 ;
        RECT 71.520 68.620 71.690 68.790 ;
        RECT 71.880 68.620 72.050 68.790 ;
        RECT 72.720 68.620 72.890 68.790 ;
        RECT 73.080 68.620 73.250 68.790 ;
        RECT 73.440 68.620 73.610 68.790 ;
        RECT 74.280 68.620 74.450 68.790 ;
        RECT 74.640 68.620 74.810 68.790 ;
        RECT 75.000 68.620 75.170 68.790 ;
        RECT 76.060 68.620 76.230 68.790 ;
        RECT 76.500 68.620 76.670 68.790 ;
        RECT 76.940 68.620 77.110 68.790 ;
        RECT 77.350 68.620 77.520 68.790 ;
        RECT 77.860 68.620 78.030 68.790 ;
        RECT 78.220 68.620 78.390 68.790 ;
        RECT 78.580 68.620 78.750 68.790 ;
        RECT 78.940 68.620 79.110 68.790 ;
        RECT 79.300 68.620 79.470 68.790 ;
        RECT 81.340 68.620 81.510 68.790 ;
        RECT 81.780 68.620 81.950 68.790 ;
        RECT 82.220 68.620 82.390 68.790 ;
        RECT 82.630 68.620 82.800 68.790 ;
        RECT 83.680 68.620 83.850 68.790 ;
        RECT 84.040 68.620 84.210 68.790 ;
        RECT 84.400 68.620 84.570 68.790 ;
        RECT 84.760 68.620 84.930 68.790 ;
        RECT 85.120 68.620 85.290 68.790 ;
        RECT 85.930 68.620 86.100 68.790 ;
        RECT 86.290 68.620 86.460 68.790 ;
        RECT 86.650 68.620 86.820 68.790 ;
        RECT 87.010 68.620 87.180 68.790 ;
        RECT 88.110 68.630 88.280 68.800 ;
        RECT 88.550 68.630 88.720 68.800 ;
        RECT 88.960 68.630 89.130 68.800 ;
        RECT 89.390 68.630 89.560 68.800 ;
        RECT 89.830 68.630 90.000 68.800 ;
        RECT 90.240 68.630 90.410 68.800 ;
        RECT 92.270 68.620 92.440 68.790 ;
        RECT 92.630 68.620 92.800 68.790 ;
        RECT 92.990 68.620 93.160 68.790 ;
        RECT 93.910 68.620 94.080 68.790 ;
        RECT 94.270 68.620 94.440 68.790 ;
        RECT 98.870 68.620 99.040 68.790 ;
        RECT 99.230 68.620 99.400 68.790 ;
        RECT 99.590 68.620 99.760 68.790 ;
        RECT 102.840 68.620 103.010 68.790 ;
        RECT 103.200 68.620 103.370 68.790 ;
        RECT 103.560 68.620 103.730 68.790 ;
        RECT 105.450 68.620 105.620 68.790 ;
        RECT 105.810 68.620 105.980 68.790 ;
        RECT 106.170 68.620 106.340 68.790 ;
        RECT 107.790 68.630 107.960 68.800 ;
        RECT 108.230 68.630 108.400 68.800 ;
        RECT 108.640 68.630 108.810 68.800 ;
        RECT 109.070 68.630 109.240 68.800 ;
        RECT 109.510 68.630 109.680 68.800 ;
        RECT 109.920 68.630 110.090 68.800 ;
        RECT 111.520 68.620 111.690 68.790 ;
        RECT 111.880 68.620 112.050 68.790 ;
        RECT 112.240 68.620 112.410 68.790 ;
        RECT 114.460 68.620 114.630 68.790 ;
        RECT 114.900 68.620 115.070 68.790 ;
        RECT 115.340 68.620 115.510 68.790 ;
        RECT 115.750 68.620 115.920 68.790 ;
        RECT 116.280 68.620 116.450 68.790 ;
        RECT 116.640 68.620 116.810 68.790 ;
        RECT 117.000 68.620 117.170 68.790 ;
        RECT 117.840 68.620 118.010 68.790 ;
        RECT 118.200 68.620 118.370 68.790 ;
        RECT 118.560 68.620 118.730 68.790 ;
        RECT 119.400 68.620 119.570 68.790 ;
        RECT 119.760 68.620 119.930 68.790 ;
        RECT 120.120 68.620 120.290 68.790 ;
        RECT 121.180 68.620 121.350 68.790 ;
        RECT 121.620 68.620 121.790 68.790 ;
        RECT 122.060 68.620 122.230 68.790 ;
        RECT 122.470 68.620 122.640 68.790 ;
        RECT 123.000 68.620 123.170 68.790 ;
        RECT 123.360 68.620 123.530 68.790 ;
        RECT 124.270 68.620 124.440 68.790 ;
        RECT 124.630 68.620 124.800 68.790 ;
        RECT 124.990 68.620 125.160 68.790 ;
        RECT 126.990 68.630 127.160 68.800 ;
        RECT 127.430 68.630 127.600 68.800 ;
        RECT 127.840 68.630 128.010 68.800 ;
        RECT 128.270 68.630 128.440 68.800 ;
        RECT 128.710 68.630 128.880 68.800 ;
        RECT 129.120 68.630 129.290 68.800 ;
        RECT 131.110 68.620 131.280 68.790 ;
        RECT 131.470 68.620 131.640 68.790 ;
        RECT 131.830 68.620 132.000 68.790 ;
        RECT 132.190 68.620 132.360 68.790 ;
        RECT 133.180 68.620 133.350 68.790 ;
        RECT 133.620 68.620 133.790 68.790 ;
        RECT 134.060 68.620 134.230 68.790 ;
        RECT 134.470 68.620 134.640 68.790 ;
        RECT 135.000 68.620 135.170 68.790 ;
        RECT 135.360 68.620 135.530 68.790 ;
        RECT 137.070 68.630 137.240 68.800 ;
        RECT 137.510 68.630 137.680 68.800 ;
        RECT 137.920 68.630 138.090 68.800 ;
        RECT 138.350 68.630 138.520 68.800 ;
        RECT 138.790 68.630 138.960 68.800 ;
        RECT 139.200 68.630 139.370 68.800 ;
        RECT 140.380 68.620 140.550 68.790 ;
        RECT 140.820 68.620 140.990 68.790 ;
        RECT 141.260 68.620 141.430 68.790 ;
        RECT 141.670 68.620 141.840 68.790 ;
        RECT 5.920 60.960 6.090 61.140 ;
        RECT 6.400 60.960 6.570 61.140 ;
        RECT 6.880 60.960 7.050 61.140 ;
        RECT 7.360 60.960 7.530 61.140 ;
        RECT 7.840 60.960 8.010 61.140 ;
        RECT 8.320 60.960 8.490 61.140 ;
        RECT 8.800 60.960 8.970 61.140 ;
        RECT 9.280 60.960 9.450 61.140 ;
        RECT 9.760 60.960 9.930 61.140 ;
        RECT 10.240 60.960 10.410 61.140 ;
        RECT 10.720 60.960 10.890 61.140 ;
        RECT 11.200 60.960 11.370 61.140 ;
        RECT 11.680 60.960 11.850 61.140 ;
        RECT 12.160 60.960 12.330 61.140 ;
        RECT 12.640 60.960 12.810 61.140 ;
        RECT 13.120 60.960 13.290 61.140 ;
        RECT 13.600 60.960 13.770 61.140 ;
        RECT 14.080 60.960 14.250 61.140 ;
        RECT 14.560 60.960 14.730 61.140 ;
        RECT 15.040 60.960 15.210 61.140 ;
        RECT 15.520 60.960 15.690 61.140 ;
        RECT 16.000 60.960 16.170 61.140 ;
        RECT 16.480 60.960 16.650 61.140 ;
        RECT 16.960 60.960 17.130 61.140 ;
        RECT 17.440 60.960 17.610 61.140 ;
        RECT 17.920 60.960 18.090 61.140 ;
        RECT 18.400 60.960 18.570 61.140 ;
        RECT 18.880 60.960 19.050 61.140 ;
        RECT 19.360 60.960 19.530 61.140 ;
        RECT 19.840 60.960 20.010 61.140 ;
        RECT 20.320 60.960 20.490 61.140 ;
        RECT 20.800 60.960 20.970 61.140 ;
        RECT 21.280 60.960 21.450 61.140 ;
        RECT 21.760 60.960 21.930 61.140 ;
        RECT 22.240 60.960 22.410 61.140 ;
        RECT 22.720 60.960 22.890 61.140 ;
        RECT 23.200 60.960 23.370 61.140 ;
        RECT 23.680 60.960 23.850 61.140 ;
        RECT 24.160 60.960 24.330 61.140 ;
        RECT 24.640 60.960 24.810 61.140 ;
        RECT 25.120 60.960 25.290 61.140 ;
        RECT 25.600 60.960 25.770 61.140 ;
        RECT 26.080 60.960 26.250 61.140 ;
        RECT 26.560 60.960 26.730 61.140 ;
        RECT 27.040 60.960 27.210 61.140 ;
        RECT 27.520 60.960 27.690 61.140 ;
        RECT 28.000 60.960 28.170 61.140 ;
        RECT 28.480 60.960 28.650 61.140 ;
        RECT 28.960 60.960 29.130 61.140 ;
        RECT 29.440 60.960 29.610 61.140 ;
        RECT 29.920 60.960 30.090 61.140 ;
        RECT 30.400 60.960 30.570 61.140 ;
        RECT 30.880 60.960 31.050 61.140 ;
        RECT 31.360 60.960 31.530 61.140 ;
        RECT 31.840 60.960 32.010 61.140 ;
        RECT 32.320 60.960 32.490 61.140 ;
        RECT 32.800 60.960 32.970 61.140 ;
        RECT 33.280 60.960 33.450 61.140 ;
        RECT 33.760 60.960 33.930 61.140 ;
        RECT 34.240 60.960 34.410 61.140 ;
        RECT 34.720 60.960 34.890 61.140 ;
        RECT 35.200 60.960 35.370 61.140 ;
        RECT 35.680 60.960 35.850 61.140 ;
        RECT 36.160 60.960 36.330 61.140 ;
        RECT 36.640 60.960 36.810 61.140 ;
        RECT 37.120 60.960 37.290 61.140 ;
        RECT 37.600 60.960 37.770 61.140 ;
        RECT 38.080 60.960 38.250 61.140 ;
        RECT 38.560 60.960 38.730 61.140 ;
        RECT 39.040 60.960 39.210 61.140 ;
        RECT 39.520 60.960 39.690 61.140 ;
        RECT 40.000 60.960 40.170 61.140 ;
        RECT 40.480 60.960 40.650 61.140 ;
        RECT 40.960 60.960 41.130 61.140 ;
        RECT 41.440 60.960 41.610 61.140 ;
        RECT 41.920 60.960 42.090 61.140 ;
        RECT 42.400 60.960 42.570 61.140 ;
        RECT 42.880 60.960 43.050 61.140 ;
        RECT 43.360 60.960 43.530 61.140 ;
        RECT 43.840 60.960 44.010 61.140 ;
        RECT 44.320 60.960 44.490 61.140 ;
        RECT 44.800 60.960 44.970 61.140 ;
        RECT 45.280 60.960 45.450 61.140 ;
        RECT 45.760 60.960 45.930 61.140 ;
        RECT 46.240 60.960 46.410 61.140 ;
        RECT 46.720 60.960 46.890 61.140 ;
        RECT 47.200 60.960 47.370 61.140 ;
        RECT 47.680 60.960 47.850 61.140 ;
        RECT 48.160 60.960 48.330 61.140 ;
        RECT 48.640 60.960 48.810 61.140 ;
        RECT 49.120 60.960 49.290 61.140 ;
        RECT 49.600 60.960 49.770 61.140 ;
        RECT 50.080 60.960 50.250 61.140 ;
        RECT 50.560 60.960 50.730 61.140 ;
        RECT 51.040 60.960 51.210 61.140 ;
        RECT 51.520 60.960 51.690 61.140 ;
        RECT 52.000 60.960 52.170 61.140 ;
        RECT 52.480 60.960 52.650 61.140 ;
        RECT 52.960 60.960 53.130 61.140 ;
        RECT 53.440 60.960 53.610 61.140 ;
        RECT 53.920 60.960 54.090 61.140 ;
        RECT 54.400 60.960 54.570 61.140 ;
        RECT 54.880 60.960 55.050 61.140 ;
        RECT 55.360 60.960 55.530 61.140 ;
        RECT 55.840 60.960 56.010 61.140 ;
        RECT 56.320 60.960 56.490 61.140 ;
        RECT 56.800 60.960 56.970 61.140 ;
        RECT 57.280 60.960 57.450 61.140 ;
        RECT 57.760 60.960 57.930 61.140 ;
        RECT 58.240 60.960 58.410 61.140 ;
        RECT 58.720 60.960 58.890 61.140 ;
        RECT 59.200 60.960 59.370 61.140 ;
        RECT 59.680 60.960 59.850 61.140 ;
        RECT 60.160 60.960 60.330 61.140 ;
        RECT 60.640 60.960 60.810 61.140 ;
        RECT 61.120 60.960 61.290 61.140 ;
        RECT 61.600 60.960 61.770 61.140 ;
        RECT 62.080 60.960 62.250 61.140 ;
        RECT 62.560 60.960 62.730 61.140 ;
        RECT 63.040 60.960 63.210 61.140 ;
        RECT 63.520 60.960 63.690 61.140 ;
        RECT 64.000 60.960 64.170 61.140 ;
        RECT 64.480 60.960 64.650 61.140 ;
        RECT 64.960 60.960 65.130 61.140 ;
        RECT 65.440 60.960 65.610 61.140 ;
        RECT 65.920 60.960 66.090 61.140 ;
        RECT 66.400 60.960 66.570 61.140 ;
        RECT 66.880 60.960 67.050 61.140 ;
        RECT 67.360 60.960 67.530 61.140 ;
        RECT 67.840 60.960 68.010 61.140 ;
        RECT 68.320 60.960 68.490 61.140 ;
        RECT 68.800 60.960 68.970 61.140 ;
        RECT 69.280 60.960 69.450 61.140 ;
        RECT 69.760 60.960 69.930 61.140 ;
        RECT 70.240 60.960 70.410 61.140 ;
        RECT 70.720 60.960 70.890 61.140 ;
        RECT 71.200 60.960 71.370 61.140 ;
        RECT 71.680 60.960 71.850 61.140 ;
        RECT 72.160 60.960 72.330 61.140 ;
        RECT 72.640 60.960 72.810 61.140 ;
        RECT 73.120 60.960 73.290 61.140 ;
        RECT 73.600 60.960 73.770 61.140 ;
        RECT 74.080 60.960 74.250 61.140 ;
        RECT 74.560 60.960 74.730 61.140 ;
        RECT 75.040 60.960 75.210 61.140 ;
        RECT 75.520 60.960 75.690 61.140 ;
        RECT 76.000 60.960 76.170 61.140 ;
        RECT 76.480 60.960 76.650 61.140 ;
        RECT 76.960 60.960 77.130 61.140 ;
        RECT 77.440 60.960 77.610 61.140 ;
        RECT 77.920 60.960 78.090 61.140 ;
        RECT 78.400 60.960 78.570 61.140 ;
        RECT 78.880 60.960 79.050 61.140 ;
        RECT 79.360 60.960 79.530 61.140 ;
        RECT 79.840 60.960 80.010 61.140 ;
        RECT 80.320 60.960 80.490 61.140 ;
        RECT 80.800 60.960 80.970 61.140 ;
        RECT 81.280 60.960 81.450 61.140 ;
        RECT 81.760 60.960 81.930 61.140 ;
        RECT 82.240 60.960 82.410 61.140 ;
        RECT 82.720 60.960 82.890 61.140 ;
        RECT 83.200 60.960 83.370 61.140 ;
        RECT 83.680 60.960 83.850 61.140 ;
        RECT 84.160 60.960 84.330 61.140 ;
        RECT 84.640 60.960 84.810 61.140 ;
        RECT 85.120 60.960 85.290 61.140 ;
        RECT 85.600 60.960 85.770 61.140 ;
        RECT 86.080 60.960 86.250 61.140 ;
        RECT 86.560 60.960 86.730 61.140 ;
        RECT 87.040 60.960 87.210 61.140 ;
        RECT 87.520 60.960 87.690 61.140 ;
        RECT 88.000 60.960 88.170 61.140 ;
        RECT 88.480 60.960 88.650 61.140 ;
        RECT 88.960 60.960 89.130 61.140 ;
        RECT 89.440 60.960 89.610 61.140 ;
        RECT 89.920 60.960 90.090 61.140 ;
        RECT 90.400 60.960 90.570 61.140 ;
        RECT 90.880 60.960 91.050 61.140 ;
      LAYER li1 ;
        RECT 91.200 60.960 91.680 61.140 ;
      LAYER li1 ;
        RECT 91.840 60.960 92.010 61.140 ;
        RECT 92.320 60.960 92.490 61.140 ;
        RECT 92.800 60.960 92.970 61.140 ;
        RECT 93.280 60.960 93.450 61.140 ;
        RECT 93.760 60.960 93.930 61.140 ;
        RECT 94.240 60.960 94.410 61.140 ;
        RECT 94.720 60.960 94.890 61.140 ;
        RECT 95.200 60.960 95.370 61.140 ;
        RECT 95.680 60.960 95.850 61.140 ;
        RECT 96.160 60.960 96.330 61.140 ;
        RECT 96.640 60.960 96.810 61.140 ;
        RECT 97.120 60.960 97.290 61.140 ;
        RECT 97.600 60.960 97.770 61.140 ;
        RECT 98.080 60.960 98.250 61.140 ;
        RECT 98.560 60.960 98.730 61.140 ;
        RECT 99.040 60.960 99.210 61.140 ;
        RECT 99.520 60.960 99.690 61.140 ;
        RECT 100.000 60.960 100.170 61.140 ;
        RECT 100.480 60.960 100.650 61.140 ;
        RECT 100.960 60.960 101.130 61.140 ;
        RECT 101.440 60.960 101.610 61.140 ;
        RECT 101.920 60.960 102.090 61.140 ;
        RECT 102.400 60.960 102.570 61.140 ;
        RECT 102.880 60.960 103.050 61.140 ;
        RECT 103.360 60.960 103.530 61.140 ;
        RECT 103.840 60.960 104.010 61.140 ;
        RECT 104.320 60.960 104.490 61.140 ;
        RECT 104.800 60.960 104.970 61.140 ;
        RECT 105.280 60.960 105.450 61.140 ;
      LAYER li1 ;
        RECT 105.600 60.960 106.080 61.140 ;
      LAYER li1 ;
        RECT 106.240 60.960 106.410 61.140 ;
        RECT 106.720 60.960 106.890 61.140 ;
        RECT 107.200 60.960 107.370 61.140 ;
        RECT 107.680 60.960 107.850 61.140 ;
        RECT 108.160 60.960 108.330 61.140 ;
        RECT 108.640 60.960 108.810 61.140 ;
        RECT 109.120 60.960 109.290 61.140 ;
        RECT 109.600 60.960 109.770 61.140 ;
        RECT 110.080 60.960 110.250 61.140 ;
        RECT 110.560 60.960 110.730 61.140 ;
        RECT 111.040 60.960 111.210 61.140 ;
        RECT 111.520 60.960 111.690 61.140 ;
        RECT 112.000 60.960 112.170 61.140 ;
        RECT 112.480 60.960 112.650 61.140 ;
        RECT 112.960 60.960 113.130 61.140 ;
        RECT 113.440 60.960 113.610 61.140 ;
        RECT 113.920 60.960 114.090 61.140 ;
        RECT 114.400 60.960 114.570 61.140 ;
        RECT 114.880 60.960 115.050 61.140 ;
        RECT 115.360 60.960 115.530 61.140 ;
        RECT 115.840 60.960 116.010 61.140 ;
        RECT 116.320 60.960 116.490 61.140 ;
        RECT 116.800 60.960 116.970 61.140 ;
        RECT 117.280 60.960 117.450 61.140 ;
        RECT 117.760 60.960 117.930 61.140 ;
        RECT 118.240 60.960 118.410 61.140 ;
        RECT 118.720 60.960 118.890 61.140 ;
        RECT 119.200 60.960 119.370 61.140 ;
        RECT 119.680 60.960 119.850 61.140 ;
        RECT 120.160 60.960 120.330 61.140 ;
        RECT 120.640 60.960 120.810 61.140 ;
        RECT 121.120 60.960 121.290 61.140 ;
        RECT 121.600 60.960 121.770 61.140 ;
        RECT 122.080 60.960 122.250 61.140 ;
        RECT 122.560 60.960 122.730 61.140 ;
        RECT 123.040 60.960 123.210 61.140 ;
        RECT 123.520 60.960 123.690 61.140 ;
        RECT 124.000 60.960 124.170 61.140 ;
        RECT 124.480 60.960 124.650 61.140 ;
        RECT 124.960 60.960 125.130 61.140 ;
        RECT 125.440 60.960 125.610 61.140 ;
        RECT 125.920 60.960 126.090 61.140 ;
        RECT 126.400 60.960 126.570 61.140 ;
        RECT 126.880 60.960 127.050 61.140 ;
        RECT 127.360 60.960 127.530 61.140 ;
        RECT 127.840 60.960 128.010 61.140 ;
        RECT 128.320 60.960 128.490 61.140 ;
        RECT 128.800 60.960 128.970 61.140 ;
        RECT 129.280 60.960 129.450 61.140 ;
        RECT 129.760 60.960 129.930 61.140 ;
        RECT 130.240 60.960 130.410 61.140 ;
        RECT 130.720 60.960 130.890 61.140 ;
        RECT 131.200 60.960 131.370 61.140 ;
        RECT 131.680 60.960 131.850 61.140 ;
        RECT 132.160 60.960 132.330 61.140 ;
        RECT 132.640 60.960 132.810 61.140 ;
        RECT 133.120 60.960 133.290 61.140 ;
        RECT 133.600 60.960 133.770 61.140 ;
        RECT 134.080 60.960 134.250 61.140 ;
        RECT 134.560 60.960 134.730 61.140 ;
        RECT 135.040 60.960 135.210 61.140 ;
        RECT 135.520 60.960 135.690 61.140 ;
        RECT 136.000 60.960 136.170 61.140 ;
        RECT 136.480 60.960 136.650 61.140 ;
        RECT 136.960 60.960 137.130 61.140 ;
        RECT 137.440 60.960 137.610 61.140 ;
        RECT 137.920 60.960 138.090 61.140 ;
        RECT 138.400 60.960 138.570 61.140 ;
        RECT 138.880 60.960 139.050 61.140 ;
        RECT 139.360 60.960 139.530 61.140 ;
        RECT 139.840 60.960 140.010 61.140 ;
        RECT 140.320 60.960 140.490 61.140 ;
        RECT 140.800 60.960 140.970 61.140 ;
        RECT 141.280 60.960 141.450 61.140 ;
      LAYER li1 ;
        RECT 141.600 60.960 142.080 61.140 ;
      LAYER li1 ;
        RECT 5.980 60.480 6.150 60.650 ;
        RECT 6.420 60.480 6.590 60.650 ;
        RECT 6.860 60.480 7.030 60.650 ;
        RECT 7.270 60.480 7.440 60.650 ;
        RECT 8.270 60.480 8.440 60.650 ;
        RECT 8.630 60.480 8.800 60.650 ;
        RECT 8.990 60.480 9.160 60.650 ;
        RECT 9.910 60.480 10.080 60.650 ;
        RECT 10.270 60.480 10.440 60.650 ;
        RECT 14.870 60.480 15.040 60.650 ;
        RECT 15.230 60.480 15.400 60.650 ;
        RECT 15.590 60.480 15.760 60.650 ;
        RECT 18.840 60.480 19.010 60.650 ;
        RECT 19.200 60.480 19.370 60.650 ;
        RECT 19.560 60.480 19.730 60.650 ;
        RECT 21.450 60.480 21.620 60.650 ;
        RECT 21.810 60.480 21.980 60.650 ;
        RECT 22.170 60.480 22.340 60.650 ;
        RECT 23.260 60.480 23.430 60.650 ;
        RECT 23.700 60.480 23.870 60.650 ;
        RECT 24.140 60.480 24.310 60.650 ;
        RECT 24.550 60.480 24.720 60.650 ;
        RECT 25.510 60.480 25.680 60.650 ;
        RECT 25.870 60.480 26.040 60.650 ;
        RECT 26.230 60.480 26.400 60.650 ;
        RECT 26.590 60.480 26.760 60.650 ;
        RECT 27.580 60.480 27.750 60.650 ;
        RECT 28.020 60.480 28.190 60.650 ;
        RECT 28.460 60.480 28.630 60.650 ;
        RECT 28.870 60.480 29.040 60.650 ;
        RECT 29.400 60.480 29.570 60.650 ;
        RECT 29.760 60.480 29.930 60.650 ;
        RECT 30.120 60.480 30.290 60.650 ;
        RECT 30.960 60.480 31.130 60.650 ;
        RECT 31.320 60.480 31.490 60.650 ;
        RECT 31.680 60.480 31.850 60.650 ;
        RECT 32.520 60.480 32.690 60.650 ;
        RECT 32.880 60.480 33.050 60.650 ;
        RECT 33.240 60.480 33.410 60.650 ;
        RECT 34.300 60.480 34.470 60.650 ;
        RECT 34.740 60.480 34.910 60.650 ;
        RECT 35.180 60.480 35.350 60.650 ;
        RECT 35.590 60.480 35.760 60.650 ;
        RECT 36.120 60.480 36.290 60.650 ;
        RECT 36.480 60.480 36.650 60.650 ;
        RECT 36.840 60.480 37.010 60.650 ;
        RECT 37.680 60.480 37.850 60.650 ;
        RECT 38.040 60.480 38.210 60.650 ;
        RECT 38.400 60.480 38.570 60.650 ;
        RECT 39.240 60.480 39.410 60.650 ;
        RECT 39.600 60.480 39.770 60.650 ;
        RECT 39.960 60.480 40.130 60.650 ;
        RECT 41.020 60.480 41.190 60.650 ;
        RECT 41.460 60.480 41.630 60.650 ;
        RECT 41.900 60.480 42.070 60.650 ;
        RECT 42.310 60.480 42.480 60.650 ;
        RECT 42.840 60.480 43.010 60.650 ;
        RECT 43.200 60.480 43.370 60.650 ;
        RECT 43.560 60.480 43.730 60.650 ;
        RECT 44.400 60.480 44.570 60.650 ;
        RECT 44.760 60.480 44.930 60.650 ;
        RECT 45.120 60.480 45.290 60.650 ;
        RECT 45.960 60.480 46.130 60.650 ;
        RECT 46.320 60.480 46.490 60.650 ;
        RECT 46.680 60.480 46.850 60.650 ;
        RECT 47.740 60.480 47.910 60.650 ;
        RECT 48.180 60.480 48.350 60.650 ;
        RECT 48.620 60.480 48.790 60.650 ;
        RECT 49.030 60.480 49.200 60.650 ;
        RECT 50.040 60.480 50.210 60.650 ;
        RECT 50.400 60.480 50.570 60.650 ;
        RECT 50.760 60.480 50.930 60.650 ;
        RECT 51.600 60.480 51.770 60.650 ;
        RECT 51.960 60.480 52.130 60.650 ;
        RECT 52.320 60.480 52.490 60.650 ;
        RECT 53.160 60.480 53.330 60.650 ;
        RECT 53.520 60.480 53.690 60.650 ;
        RECT 53.880 60.480 54.050 60.650 ;
        RECT 54.940 60.480 55.110 60.650 ;
        RECT 55.380 60.480 55.550 60.650 ;
        RECT 55.820 60.480 55.990 60.650 ;
        RECT 56.230 60.480 56.400 60.650 ;
        RECT 56.760 60.480 56.930 60.650 ;
        RECT 57.120 60.480 57.290 60.650 ;
        RECT 58.030 60.480 58.200 60.650 ;
        RECT 58.390 60.480 58.560 60.650 ;
        RECT 58.750 60.480 58.920 60.650 ;
        RECT 60.220 60.480 60.390 60.650 ;
        RECT 60.660 60.480 60.830 60.650 ;
        RECT 61.100 60.480 61.270 60.650 ;
        RECT 61.510 60.480 61.680 60.650 ;
        RECT 62.510 60.480 62.680 60.650 ;
        RECT 62.870 60.480 63.040 60.650 ;
        RECT 63.230 60.480 63.400 60.650 ;
        RECT 64.150 60.480 64.320 60.650 ;
        RECT 64.510 60.480 64.680 60.650 ;
        RECT 69.110 60.480 69.280 60.650 ;
        RECT 69.470 60.480 69.640 60.650 ;
        RECT 69.830 60.480 70.000 60.650 ;
        RECT 73.080 60.480 73.250 60.650 ;
        RECT 73.440 60.480 73.610 60.650 ;
        RECT 73.800 60.480 73.970 60.650 ;
        RECT 75.690 60.480 75.860 60.650 ;
        RECT 76.050 60.480 76.220 60.650 ;
        RECT 76.410 60.480 76.580 60.650 ;
        RECT 77.500 60.480 77.670 60.650 ;
        RECT 77.940 60.480 78.110 60.650 ;
        RECT 78.380 60.480 78.550 60.650 ;
        RECT 78.790 60.480 78.960 60.650 ;
        RECT 79.320 60.480 79.490 60.650 ;
        RECT 79.680 60.480 79.850 60.650 ;
        RECT 80.040 60.480 80.210 60.650 ;
        RECT 80.880 60.480 81.050 60.650 ;
        RECT 81.240 60.480 81.410 60.650 ;
        RECT 81.600 60.480 81.770 60.650 ;
        RECT 82.440 60.480 82.610 60.650 ;
        RECT 82.800 60.480 82.970 60.650 ;
        RECT 83.160 60.480 83.330 60.650 ;
        RECT 84.750 60.490 84.920 60.660 ;
        RECT 85.190 60.490 85.360 60.660 ;
        RECT 85.600 60.490 85.770 60.660 ;
        RECT 86.030 60.490 86.200 60.660 ;
        RECT 86.470 60.490 86.640 60.660 ;
        RECT 86.880 60.490 87.050 60.660 ;
        RECT 87.960 60.480 88.130 60.650 ;
        RECT 88.320 60.480 88.490 60.650 ;
        RECT 88.680 60.480 88.850 60.650 ;
        RECT 89.520 60.480 89.690 60.650 ;
        RECT 89.880 60.480 90.050 60.650 ;
        RECT 90.240 60.480 90.410 60.650 ;
        RECT 91.080 60.480 91.250 60.650 ;
        RECT 91.440 60.480 91.610 60.650 ;
        RECT 91.800 60.480 91.970 60.650 ;
        RECT 92.860 60.480 93.030 60.650 ;
        RECT 93.300 60.480 93.470 60.650 ;
        RECT 93.740 60.480 93.910 60.650 ;
        RECT 94.150 60.480 94.320 60.650 ;
        RECT 94.680 60.480 94.850 60.650 ;
        RECT 95.040 60.480 95.210 60.650 ;
        RECT 95.400 60.480 95.570 60.650 ;
        RECT 96.240 60.480 96.410 60.650 ;
        RECT 96.600 60.480 96.770 60.650 ;
        RECT 96.960 60.480 97.130 60.650 ;
        RECT 97.800 60.480 97.970 60.650 ;
        RECT 98.160 60.480 98.330 60.650 ;
        RECT 98.520 60.480 98.690 60.650 ;
        RECT 99.580 60.480 99.750 60.650 ;
        RECT 100.020 60.480 100.190 60.650 ;
        RECT 100.460 60.480 100.630 60.650 ;
        RECT 100.870 60.480 101.040 60.650 ;
        RECT 103.040 60.480 103.210 60.650 ;
        RECT 103.400 60.480 103.570 60.650 ;
        RECT 103.760 60.480 103.930 60.650 ;
        RECT 104.120 60.480 104.290 60.650 ;
        RECT 104.480 60.480 104.650 60.650 ;
        RECT 105.340 60.480 105.510 60.650 ;
        RECT 105.700 60.480 105.870 60.650 ;
        RECT 107.740 60.480 107.910 60.650 ;
        RECT 108.180 60.480 108.350 60.650 ;
        RECT 108.620 60.480 108.790 60.650 ;
        RECT 109.030 60.480 109.200 60.650 ;
        RECT 109.560 60.480 109.730 60.650 ;
        RECT 109.920 60.480 110.090 60.650 ;
        RECT 110.280 60.480 110.450 60.650 ;
        RECT 111.120 60.480 111.290 60.650 ;
        RECT 111.480 60.480 111.650 60.650 ;
        RECT 111.840 60.480 112.010 60.650 ;
        RECT 112.680 60.480 112.850 60.650 ;
        RECT 113.040 60.480 113.210 60.650 ;
        RECT 113.400 60.480 113.570 60.650 ;
        RECT 114.460 60.480 114.630 60.650 ;
        RECT 114.900 60.480 115.070 60.650 ;
        RECT 115.340 60.480 115.510 60.650 ;
        RECT 115.750 60.480 115.920 60.650 ;
        RECT 116.280 60.480 116.450 60.650 ;
        RECT 116.640 60.480 116.810 60.650 ;
        RECT 117.000 60.480 117.170 60.650 ;
        RECT 117.840 60.480 118.010 60.650 ;
        RECT 118.200 60.480 118.370 60.650 ;
        RECT 118.560 60.480 118.730 60.650 ;
        RECT 119.400 60.480 119.570 60.650 ;
        RECT 119.760 60.480 119.930 60.650 ;
        RECT 120.120 60.480 120.290 60.650 ;
        RECT 121.180 60.480 121.350 60.650 ;
        RECT 121.620 60.480 121.790 60.650 ;
        RECT 122.060 60.480 122.230 60.650 ;
        RECT 122.470 60.480 122.640 60.650 ;
        RECT 123.000 60.480 123.170 60.650 ;
        RECT 123.360 60.480 123.530 60.650 ;
        RECT 123.720 60.480 123.890 60.650 ;
        RECT 124.560 60.480 124.730 60.650 ;
        RECT 124.920 60.480 125.090 60.650 ;
        RECT 125.280 60.480 125.450 60.650 ;
        RECT 126.120 60.480 126.290 60.650 ;
        RECT 126.480 60.480 126.650 60.650 ;
        RECT 126.840 60.480 127.010 60.650 ;
        RECT 127.900 60.480 128.070 60.650 ;
        RECT 128.340 60.480 128.510 60.650 ;
        RECT 128.780 60.480 128.950 60.650 ;
        RECT 129.190 60.480 129.360 60.650 ;
        RECT 129.720 60.480 129.890 60.650 ;
        RECT 130.080 60.480 130.250 60.650 ;
        RECT 130.440 60.480 130.610 60.650 ;
        RECT 131.280 60.480 131.450 60.650 ;
        RECT 131.640 60.480 131.810 60.650 ;
        RECT 132.000 60.480 132.170 60.650 ;
        RECT 132.840 60.480 133.010 60.650 ;
        RECT 133.200 60.480 133.370 60.650 ;
        RECT 133.560 60.480 133.730 60.650 ;
        RECT 134.620 60.480 134.790 60.650 ;
        RECT 135.060 60.480 135.230 60.650 ;
        RECT 135.500 60.480 135.670 60.650 ;
        RECT 135.910 60.480 136.080 60.650 ;
        RECT 137.920 60.480 138.090 60.650 ;
        RECT 138.280 60.480 138.450 60.650 ;
        RECT 138.940 60.480 139.110 60.650 ;
        RECT 139.380 60.480 139.550 60.650 ;
        RECT 139.820 60.480 139.990 60.650 ;
        RECT 140.230 60.480 140.400 60.650 ;
        RECT 5.920 52.820 6.090 53.000 ;
        RECT 6.400 52.820 6.570 53.000 ;
        RECT 6.880 52.820 7.050 53.000 ;
        RECT 7.360 52.820 7.530 53.000 ;
      LAYER li1 ;
        RECT 7.680 52.820 8.160 53.000 ;
      LAYER li1 ;
        RECT 8.320 52.820 8.490 53.000 ;
        RECT 8.800 52.820 8.970 53.000 ;
        RECT 9.280 52.820 9.450 53.000 ;
        RECT 9.760 52.820 9.930 53.000 ;
        RECT 10.240 52.820 10.410 53.000 ;
        RECT 10.720 52.820 10.890 53.000 ;
        RECT 11.200 52.820 11.370 53.000 ;
        RECT 11.680 52.820 11.850 53.000 ;
        RECT 12.160 52.820 12.330 53.000 ;
        RECT 12.640 52.820 12.810 53.000 ;
        RECT 13.120 52.820 13.290 53.000 ;
        RECT 13.600 52.820 13.770 53.000 ;
        RECT 14.080 52.820 14.250 53.000 ;
        RECT 14.560 52.820 14.730 53.000 ;
        RECT 15.040 52.820 15.210 53.000 ;
        RECT 15.520 52.820 15.690 53.000 ;
        RECT 16.000 52.820 16.170 53.000 ;
        RECT 16.480 52.820 16.650 53.000 ;
        RECT 16.960 52.820 17.130 53.000 ;
        RECT 17.440 52.820 17.610 53.000 ;
        RECT 17.920 52.820 18.090 53.000 ;
        RECT 18.400 52.820 18.570 53.000 ;
        RECT 18.880 52.820 19.050 53.000 ;
        RECT 19.360 52.820 19.530 53.000 ;
        RECT 19.840 52.820 20.010 53.000 ;
        RECT 20.320 52.820 20.490 53.000 ;
        RECT 20.800 52.820 20.970 53.000 ;
        RECT 21.280 52.820 21.450 53.000 ;
        RECT 21.760 52.820 21.930 53.000 ;
        RECT 22.240 52.820 22.410 53.000 ;
        RECT 22.720 52.820 22.890 53.000 ;
        RECT 23.200 52.820 23.370 53.000 ;
        RECT 23.680 52.820 23.850 53.000 ;
        RECT 24.160 52.820 24.330 53.000 ;
        RECT 24.640 52.820 24.810 53.000 ;
        RECT 25.120 52.820 25.290 53.000 ;
        RECT 25.600 52.820 25.770 53.000 ;
        RECT 26.080 52.820 26.250 53.000 ;
        RECT 26.560 52.820 26.730 53.000 ;
        RECT 27.040 52.820 27.210 53.000 ;
        RECT 27.520 52.820 27.690 53.000 ;
        RECT 28.000 52.820 28.170 53.000 ;
        RECT 28.480 52.820 28.650 53.000 ;
        RECT 28.960 52.820 29.130 53.000 ;
        RECT 29.440 52.820 29.610 53.000 ;
        RECT 29.920 52.820 30.090 53.000 ;
        RECT 30.400 52.820 30.570 53.000 ;
        RECT 30.880 52.820 31.050 53.000 ;
        RECT 31.360 52.820 31.530 53.000 ;
        RECT 31.840 52.820 32.010 53.000 ;
        RECT 32.320 52.820 32.490 53.000 ;
        RECT 32.800 52.820 32.970 53.000 ;
        RECT 33.280 52.820 33.450 53.000 ;
        RECT 33.760 52.820 33.930 53.000 ;
        RECT 34.240 52.820 34.410 53.000 ;
        RECT 34.720 52.820 34.890 53.000 ;
        RECT 35.200 52.820 35.370 53.000 ;
        RECT 35.680 52.820 35.850 53.000 ;
        RECT 36.160 52.820 36.330 53.000 ;
        RECT 36.640 52.820 36.810 53.000 ;
        RECT 37.120 52.820 37.290 53.000 ;
        RECT 37.600 52.820 37.770 53.000 ;
        RECT 38.080 52.820 38.250 53.000 ;
        RECT 38.560 52.820 38.730 53.000 ;
        RECT 39.040 52.820 39.210 53.000 ;
        RECT 39.520 52.820 39.690 53.000 ;
        RECT 40.000 52.820 40.170 53.000 ;
        RECT 40.480 52.820 40.650 53.000 ;
        RECT 40.960 52.820 41.130 53.000 ;
        RECT 41.440 52.820 41.610 53.000 ;
        RECT 41.920 52.820 42.090 53.000 ;
        RECT 42.400 52.820 42.570 53.000 ;
        RECT 42.880 52.820 43.050 53.000 ;
        RECT 43.360 52.820 43.530 53.000 ;
        RECT 43.840 52.820 44.010 53.000 ;
        RECT 44.320 52.820 44.490 53.000 ;
        RECT 44.800 52.820 44.970 53.000 ;
        RECT 45.280 52.820 45.450 53.000 ;
        RECT 45.760 52.820 45.930 53.000 ;
        RECT 46.240 52.820 46.410 53.000 ;
        RECT 46.720 52.820 46.890 53.000 ;
        RECT 47.200 52.820 47.370 53.000 ;
      LAYER li1 ;
        RECT 47.520 52.820 48.000 53.000 ;
      LAYER li1 ;
        RECT 48.160 52.820 48.330 53.000 ;
        RECT 48.640 52.820 48.810 53.000 ;
        RECT 49.120 52.820 49.290 53.000 ;
        RECT 49.600 52.820 49.770 53.000 ;
        RECT 50.080 52.820 50.250 53.000 ;
        RECT 50.560 52.820 50.730 53.000 ;
        RECT 51.040 52.820 51.210 53.000 ;
        RECT 51.520 52.820 51.690 53.000 ;
        RECT 52.000 52.820 52.170 53.000 ;
        RECT 52.480 52.820 52.650 53.000 ;
        RECT 52.960 52.820 53.130 53.000 ;
        RECT 53.440 52.820 53.610 53.000 ;
        RECT 53.920 52.820 54.090 53.000 ;
        RECT 54.400 52.820 54.570 53.000 ;
        RECT 54.880 52.820 55.050 53.000 ;
        RECT 55.360 52.820 55.530 53.000 ;
        RECT 55.840 52.820 56.010 53.000 ;
        RECT 56.320 52.820 56.490 53.000 ;
        RECT 56.800 52.820 56.970 53.000 ;
        RECT 57.280 52.820 57.450 53.000 ;
        RECT 57.760 52.820 57.930 53.000 ;
        RECT 58.240 52.820 58.410 53.000 ;
        RECT 58.720 52.820 58.890 53.000 ;
        RECT 59.200 52.820 59.370 53.000 ;
        RECT 59.680 52.820 59.850 53.000 ;
        RECT 60.160 52.820 60.330 53.000 ;
        RECT 60.640 52.820 60.810 53.000 ;
        RECT 61.120 52.820 61.290 53.000 ;
        RECT 61.600 52.820 61.770 53.000 ;
        RECT 62.080 52.820 62.250 53.000 ;
        RECT 62.560 52.820 62.730 53.000 ;
        RECT 63.040 52.820 63.210 53.000 ;
        RECT 63.520 52.820 63.690 53.000 ;
        RECT 64.000 52.820 64.170 53.000 ;
        RECT 64.480 52.820 64.650 53.000 ;
        RECT 64.960 52.820 65.130 53.000 ;
        RECT 65.440 52.820 65.610 53.000 ;
        RECT 65.920 52.820 66.090 53.000 ;
        RECT 66.400 52.820 66.570 53.000 ;
        RECT 66.880 52.820 67.050 53.000 ;
        RECT 67.360 52.820 67.530 53.000 ;
        RECT 67.840 52.820 68.010 53.000 ;
        RECT 68.320 52.820 68.490 53.000 ;
        RECT 68.800 52.820 68.970 53.000 ;
        RECT 69.280 52.820 69.450 53.000 ;
        RECT 69.760 52.820 69.930 53.000 ;
        RECT 70.240 52.820 70.410 53.000 ;
        RECT 70.720 52.820 70.890 53.000 ;
        RECT 71.200 52.820 71.370 53.000 ;
        RECT 71.680 52.820 71.850 53.000 ;
        RECT 72.160 52.820 72.330 53.000 ;
        RECT 72.640 52.820 72.810 53.000 ;
        RECT 73.120 52.820 73.290 53.000 ;
        RECT 73.600 52.820 73.770 53.000 ;
        RECT 74.080 52.820 74.250 53.000 ;
        RECT 74.560 52.820 74.730 53.000 ;
        RECT 75.040 52.820 75.210 53.000 ;
        RECT 75.520 52.820 75.690 53.000 ;
        RECT 76.000 52.820 76.170 53.000 ;
        RECT 76.480 52.820 76.650 53.000 ;
        RECT 76.960 52.820 77.130 53.000 ;
        RECT 77.440 52.820 77.610 53.000 ;
        RECT 77.920 52.820 78.090 53.000 ;
        RECT 78.400 52.820 78.570 53.000 ;
        RECT 78.880 52.820 79.050 53.000 ;
        RECT 79.360 52.820 79.530 53.000 ;
        RECT 79.840 52.820 80.010 53.000 ;
        RECT 80.320 52.820 80.490 53.000 ;
        RECT 80.800 52.820 80.970 53.000 ;
      LAYER li1 ;
        RECT 81.120 52.820 81.600 53.000 ;
      LAYER li1 ;
        RECT 81.760 52.820 81.930 53.000 ;
        RECT 82.240 52.820 82.410 53.000 ;
        RECT 82.720 52.820 82.890 53.000 ;
        RECT 83.200 52.820 83.370 53.000 ;
        RECT 83.680 52.820 83.850 53.000 ;
        RECT 84.160 52.820 84.330 53.000 ;
        RECT 84.640 52.820 84.810 53.000 ;
        RECT 85.120 52.820 85.290 53.000 ;
        RECT 85.600 52.820 85.770 53.000 ;
        RECT 86.080 52.820 86.250 53.000 ;
        RECT 86.560 52.820 86.730 53.000 ;
        RECT 87.040 52.820 87.210 53.000 ;
        RECT 87.520 52.820 87.690 53.000 ;
        RECT 88.000 52.820 88.170 53.000 ;
        RECT 88.480 52.820 88.650 53.000 ;
        RECT 88.960 52.820 89.130 53.000 ;
        RECT 89.440 52.820 89.610 53.000 ;
        RECT 89.920 52.820 90.090 53.000 ;
        RECT 90.400 52.820 90.570 53.000 ;
        RECT 90.880 52.820 91.050 53.000 ;
        RECT 91.360 52.820 91.530 53.000 ;
        RECT 91.840 52.820 92.010 53.000 ;
        RECT 92.320 52.820 92.490 53.000 ;
        RECT 92.800 52.820 92.970 53.000 ;
        RECT 93.280 52.820 93.450 53.000 ;
        RECT 93.760 52.820 93.930 53.000 ;
        RECT 94.240 52.820 94.410 53.000 ;
        RECT 94.720 52.820 94.890 53.000 ;
        RECT 95.200 52.820 95.370 53.000 ;
        RECT 95.680 52.820 95.850 53.000 ;
        RECT 96.160 52.820 96.330 53.000 ;
        RECT 96.640 52.820 96.810 53.000 ;
        RECT 97.120 52.820 97.290 53.000 ;
        RECT 97.600 52.820 97.770 53.000 ;
        RECT 98.080 52.820 98.250 53.000 ;
        RECT 98.560 52.820 98.730 53.000 ;
        RECT 99.040 52.820 99.210 53.000 ;
        RECT 99.520 52.820 99.690 53.000 ;
        RECT 100.000 52.820 100.170 53.000 ;
        RECT 100.480 52.820 100.650 53.000 ;
        RECT 100.960 52.820 101.130 53.000 ;
        RECT 101.440 52.820 101.610 53.000 ;
        RECT 101.920 52.820 102.090 53.000 ;
        RECT 102.400 52.820 102.570 53.000 ;
        RECT 102.880 52.820 103.050 53.000 ;
        RECT 103.360 52.820 103.530 53.000 ;
        RECT 103.840 52.820 104.010 53.000 ;
        RECT 104.320 52.820 104.490 53.000 ;
        RECT 104.800 52.820 104.970 53.000 ;
        RECT 105.280 52.820 105.450 53.000 ;
        RECT 105.760 52.820 105.930 53.000 ;
        RECT 106.240 52.820 106.410 53.000 ;
        RECT 106.720 52.820 106.890 53.000 ;
      LAYER li1 ;
        RECT 107.040 52.820 107.520 53.000 ;
      LAYER li1 ;
        RECT 107.680 52.820 107.850 53.000 ;
        RECT 108.160 52.820 108.330 53.000 ;
        RECT 108.640 52.820 108.810 53.000 ;
        RECT 109.120 52.820 109.290 53.000 ;
        RECT 109.600 52.820 109.770 53.000 ;
        RECT 110.080 52.820 110.250 53.000 ;
        RECT 110.560 52.820 110.730 53.000 ;
        RECT 111.040 52.820 111.210 53.000 ;
        RECT 111.520 52.820 111.690 53.000 ;
        RECT 112.000 52.820 112.170 53.000 ;
        RECT 112.480 52.820 112.650 53.000 ;
        RECT 112.960 52.820 113.130 53.000 ;
        RECT 113.440 52.820 113.610 53.000 ;
        RECT 113.920 52.820 114.090 53.000 ;
        RECT 114.400 52.820 114.570 53.000 ;
        RECT 114.880 52.820 115.050 53.000 ;
        RECT 115.360 52.820 115.530 53.000 ;
        RECT 115.840 52.820 116.010 53.000 ;
        RECT 116.320 52.820 116.490 53.000 ;
        RECT 116.800 52.820 116.970 53.000 ;
        RECT 117.280 52.820 117.450 53.000 ;
        RECT 117.760 52.820 117.930 53.000 ;
        RECT 118.240 52.820 118.410 53.000 ;
        RECT 118.720 52.820 118.890 53.000 ;
        RECT 119.200 52.820 119.370 53.000 ;
        RECT 119.680 52.820 119.850 53.000 ;
        RECT 120.160 52.820 120.330 53.000 ;
        RECT 120.640 52.820 120.810 53.000 ;
        RECT 121.120 52.820 121.290 53.000 ;
        RECT 121.600 52.820 121.770 53.000 ;
        RECT 122.080 52.820 122.250 53.000 ;
        RECT 122.560 52.820 122.730 53.000 ;
      LAYER li1 ;
        RECT 122.880 52.820 123.360 53.000 ;
      LAYER li1 ;
        RECT 123.520 52.820 123.690 53.000 ;
        RECT 124.000 52.820 124.170 53.000 ;
        RECT 124.480 52.820 124.650 53.000 ;
        RECT 124.960 52.820 125.130 53.000 ;
        RECT 125.440 52.820 125.610 53.000 ;
        RECT 125.920 52.820 126.090 53.000 ;
        RECT 126.400 52.820 126.570 53.000 ;
        RECT 126.880 52.820 127.050 53.000 ;
        RECT 127.360 52.820 127.530 53.000 ;
        RECT 127.840 52.820 128.010 53.000 ;
        RECT 128.320 52.820 128.490 53.000 ;
        RECT 128.800 52.820 128.970 53.000 ;
        RECT 129.280 52.820 129.450 53.000 ;
        RECT 129.760 52.820 129.930 53.000 ;
        RECT 130.240 52.820 130.410 53.000 ;
        RECT 130.720 52.820 130.890 53.000 ;
        RECT 131.200 52.820 131.370 53.000 ;
        RECT 131.680 52.820 131.850 53.000 ;
        RECT 132.160 52.820 132.330 53.000 ;
        RECT 132.640 52.820 132.810 53.000 ;
        RECT 133.120 52.820 133.290 53.000 ;
        RECT 133.600 52.820 133.770 53.000 ;
        RECT 134.080 52.820 134.250 53.000 ;
        RECT 134.560 52.820 134.730 53.000 ;
        RECT 135.040 52.820 135.210 53.000 ;
        RECT 135.520 52.820 135.690 53.000 ;
        RECT 136.000 52.820 136.170 53.000 ;
        RECT 136.480 52.820 136.650 53.000 ;
        RECT 136.960 52.820 137.130 53.000 ;
        RECT 137.440 52.820 137.610 53.000 ;
        RECT 137.920 52.820 138.090 53.000 ;
        RECT 138.400 52.820 138.570 53.000 ;
        RECT 138.880 52.820 139.050 53.000 ;
        RECT 139.360 52.820 139.530 53.000 ;
        RECT 139.840 52.820 140.010 53.000 ;
        RECT 140.320 52.820 140.490 53.000 ;
        RECT 140.800 52.820 140.970 53.000 ;
        RECT 141.280 52.820 141.450 53.000 ;
        RECT 141.760 52.820 141.930 53.000 ;
        RECT 5.980 52.340 6.150 52.510 ;
        RECT 6.420 52.340 6.590 52.510 ;
        RECT 6.860 52.340 7.030 52.510 ;
        RECT 7.270 52.340 7.440 52.510 ;
        RECT 8.280 52.340 8.450 52.510 ;
        RECT 8.640 52.340 8.810 52.510 ;
        RECT 9.820 52.340 9.990 52.510 ;
        RECT 10.260 52.340 10.430 52.510 ;
        RECT 10.700 52.340 10.870 52.510 ;
        RECT 11.110 52.340 11.280 52.510 ;
        RECT 12.070 52.340 12.240 52.510 ;
        RECT 12.430 52.340 12.600 52.510 ;
        RECT 12.790 52.340 12.960 52.510 ;
        RECT 13.150 52.340 13.320 52.510 ;
        RECT 14.140 52.340 14.310 52.510 ;
        RECT 14.580 52.340 14.750 52.510 ;
        RECT 15.020 52.340 15.190 52.510 ;
        RECT 15.430 52.340 15.600 52.510 ;
        RECT 15.960 52.340 16.130 52.510 ;
        RECT 16.320 52.340 16.490 52.510 ;
        RECT 16.680 52.340 16.850 52.510 ;
        RECT 17.040 52.340 17.210 52.510 ;
        RECT 18.460 52.340 18.630 52.510 ;
        RECT 18.900 52.340 19.070 52.510 ;
        RECT 19.340 52.340 19.510 52.510 ;
        RECT 19.750 52.340 19.920 52.510 ;
        RECT 20.280 52.340 20.450 52.510 ;
        RECT 20.640 52.340 20.810 52.510 ;
        RECT 22.300 52.340 22.470 52.510 ;
        RECT 22.660 52.340 22.830 52.510 ;
        RECT 23.020 52.340 23.190 52.510 ;
        RECT 23.380 52.340 23.550 52.510 ;
        RECT 23.740 52.340 23.910 52.510 ;
        RECT 24.220 52.340 24.390 52.510 ;
        RECT 24.660 52.340 24.830 52.510 ;
        RECT 25.100 52.340 25.270 52.510 ;
        RECT 25.510 52.340 25.680 52.510 ;
        RECT 26.520 52.340 26.690 52.510 ;
        RECT 27.030 52.340 27.200 52.510 ;
        RECT 28.710 52.340 28.880 52.510 ;
        RECT 29.070 52.340 29.240 52.510 ;
        RECT 29.430 52.340 29.600 52.510 ;
        RECT 30.460 52.340 30.630 52.510 ;
        RECT 30.900 52.340 31.070 52.510 ;
        RECT 31.340 52.340 31.510 52.510 ;
        RECT 31.750 52.340 31.920 52.510 ;
        RECT 32.280 52.340 32.450 52.510 ;
        RECT 32.640 52.340 32.810 52.510 ;
        RECT 33.000 52.340 33.170 52.510 ;
        RECT 33.840 52.340 34.010 52.510 ;
        RECT 34.200 52.340 34.370 52.510 ;
        RECT 34.560 52.340 34.730 52.510 ;
        RECT 35.400 52.340 35.570 52.510 ;
        RECT 35.760 52.340 35.930 52.510 ;
        RECT 36.120 52.340 36.290 52.510 ;
        RECT 37.180 52.340 37.350 52.510 ;
        RECT 37.620 52.340 37.790 52.510 ;
        RECT 38.060 52.340 38.230 52.510 ;
        RECT 38.470 52.340 38.640 52.510 ;
        RECT 39.000 52.340 39.170 52.510 ;
        RECT 39.360 52.340 39.530 52.510 ;
        RECT 39.720 52.340 39.890 52.510 ;
        RECT 40.560 52.340 40.730 52.510 ;
        RECT 40.920 52.340 41.090 52.510 ;
        RECT 41.280 52.340 41.450 52.510 ;
        RECT 42.120 52.340 42.290 52.510 ;
        RECT 42.480 52.340 42.650 52.510 ;
        RECT 42.840 52.340 43.010 52.510 ;
        RECT 44.430 52.350 44.600 52.520 ;
        RECT 44.870 52.350 45.040 52.520 ;
        RECT 45.280 52.350 45.450 52.520 ;
        RECT 45.710 52.350 45.880 52.520 ;
        RECT 46.150 52.350 46.320 52.520 ;
        RECT 46.560 52.350 46.730 52.520 ;
        RECT 48.120 52.340 48.290 52.510 ;
        RECT 48.480 52.340 48.650 52.510 ;
        RECT 48.840 52.340 49.010 52.510 ;
        RECT 49.680 52.340 49.850 52.510 ;
        RECT 50.040 52.340 50.210 52.510 ;
        RECT 50.400 52.340 50.570 52.510 ;
        RECT 51.240 52.340 51.410 52.510 ;
        RECT 51.600 52.340 51.770 52.510 ;
        RECT 51.960 52.340 52.130 52.510 ;
        RECT 53.550 52.350 53.720 52.520 ;
        RECT 53.990 52.350 54.160 52.520 ;
        RECT 54.400 52.350 54.570 52.520 ;
        RECT 54.830 52.350 55.000 52.520 ;
        RECT 55.270 52.350 55.440 52.520 ;
        RECT 55.680 52.350 55.850 52.520 ;
        RECT 57.720 52.340 57.890 52.510 ;
        RECT 58.080 52.340 58.250 52.510 ;
        RECT 58.440 52.340 58.610 52.510 ;
        RECT 59.280 52.340 59.450 52.510 ;
        RECT 59.640 52.340 59.810 52.510 ;
        RECT 60.000 52.340 60.170 52.510 ;
        RECT 60.840 52.340 61.010 52.510 ;
        RECT 61.200 52.340 61.370 52.510 ;
        RECT 61.560 52.340 61.730 52.510 ;
        RECT 62.620 52.340 62.790 52.510 ;
        RECT 63.060 52.340 63.230 52.510 ;
        RECT 63.500 52.340 63.670 52.510 ;
        RECT 63.910 52.340 64.080 52.510 ;
        RECT 64.440 52.340 64.610 52.510 ;
        RECT 64.800 52.340 64.970 52.510 ;
        RECT 65.160 52.340 65.330 52.510 ;
        RECT 66.000 52.340 66.170 52.510 ;
        RECT 66.360 52.340 66.530 52.510 ;
        RECT 66.720 52.340 66.890 52.510 ;
        RECT 67.560 52.340 67.730 52.510 ;
        RECT 67.920 52.340 68.090 52.510 ;
        RECT 68.280 52.340 68.450 52.510 ;
        RECT 69.340 52.340 69.510 52.510 ;
        RECT 69.780 52.340 69.950 52.510 ;
        RECT 70.220 52.340 70.390 52.510 ;
        RECT 70.630 52.340 70.800 52.510 ;
        RECT 71.160 52.340 71.330 52.510 ;
        RECT 71.520 52.340 71.690 52.510 ;
        RECT 71.880 52.340 72.050 52.510 ;
        RECT 72.720 52.340 72.890 52.510 ;
        RECT 73.080 52.340 73.250 52.510 ;
        RECT 73.440 52.340 73.610 52.510 ;
        RECT 74.280 52.340 74.450 52.510 ;
        RECT 74.640 52.340 74.810 52.510 ;
        RECT 75.000 52.340 75.170 52.510 ;
        RECT 76.060 52.340 76.230 52.510 ;
        RECT 76.500 52.340 76.670 52.510 ;
        RECT 76.940 52.340 77.110 52.510 ;
        RECT 77.350 52.340 77.520 52.510 ;
        RECT 77.880 52.340 78.050 52.510 ;
        RECT 78.240 52.340 78.410 52.510 ;
        RECT 79.420 52.340 79.590 52.510 ;
        RECT 79.860 52.340 80.030 52.510 ;
        RECT 80.300 52.340 80.470 52.510 ;
        RECT 80.710 52.340 80.880 52.510 ;
        RECT 81.720 52.340 81.890 52.510 ;
        RECT 82.080 52.340 82.250 52.510 ;
        RECT 82.440 52.340 82.610 52.510 ;
        RECT 83.280 52.340 83.450 52.510 ;
        RECT 83.640 52.340 83.810 52.510 ;
        RECT 84.000 52.340 84.170 52.510 ;
        RECT 84.840 52.340 85.010 52.510 ;
        RECT 85.200 52.340 85.370 52.510 ;
        RECT 85.560 52.340 85.730 52.510 ;
        RECT 86.620 52.340 86.790 52.510 ;
        RECT 87.060 52.340 87.230 52.510 ;
        RECT 87.500 52.340 87.670 52.510 ;
        RECT 87.910 52.340 88.080 52.510 ;
        RECT 88.440 52.340 88.610 52.510 ;
        RECT 88.800 52.340 88.970 52.510 ;
        RECT 89.160 52.340 89.330 52.510 ;
        RECT 90.000 52.340 90.170 52.510 ;
        RECT 90.360 52.340 90.530 52.510 ;
        RECT 90.720 52.340 90.890 52.510 ;
        RECT 91.560 52.340 91.730 52.510 ;
        RECT 91.920 52.340 92.090 52.510 ;
        RECT 92.280 52.340 92.450 52.510 ;
        RECT 93.340 52.340 93.510 52.510 ;
        RECT 93.780 52.340 93.950 52.510 ;
        RECT 94.220 52.340 94.390 52.510 ;
        RECT 94.630 52.340 94.800 52.510 ;
        RECT 95.160 52.340 95.330 52.510 ;
        RECT 95.520 52.340 95.690 52.510 ;
        RECT 96.700 52.340 96.870 52.510 ;
        RECT 97.140 52.340 97.310 52.510 ;
        RECT 97.580 52.340 97.750 52.510 ;
        RECT 97.990 52.340 98.160 52.510 ;
        RECT 98.520 52.340 98.690 52.510 ;
        RECT 98.880 52.340 99.050 52.510 ;
        RECT 99.240 52.340 99.410 52.510 ;
        RECT 100.080 52.340 100.250 52.510 ;
        RECT 100.440 52.340 100.610 52.510 ;
        RECT 100.800 52.340 100.970 52.510 ;
        RECT 101.640 52.340 101.810 52.510 ;
        RECT 102.000 52.340 102.170 52.510 ;
        RECT 102.360 52.340 102.530 52.510 ;
        RECT 103.950 52.350 104.120 52.520 ;
        RECT 104.390 52.350 104.560 52.520 ;
        RECT 104.800 52.350 104.970 52.520 ;
        RECT 105.230 52.350 105.400 52.520 ;
        RECT 105.670 52.350 105.840 52.520 ;
        RECT 106.080 52.350 106.250 52.520 ;
        RECT 107.640 52.340 107.810 52.510 ;
        RECT 108.000 52.340 108.170 52.510 ;
        RECT 108.360 52.340 108.530 52.510 ;
        RECT 109.200 52.340 109.370 52.510 ;
        RECT 109.560 52.340 109.730 52.510 ;
        RECT 109.920 52.340 110.090 52.510 ;
        RECT 110.760 52.340 110.930 52.510 ;
        RECT 111.120 52.340 111.290 52.510 ;
        RECT 111.480 52.340 111.650 52.510 ;
        RECT 112.540 52.340 112.710 52.510 ;
        RECT 112.980 52.340 113.150 52.510 ;
        RECT 113.420 52.340 113.590 52.510 ;
        RECT 113.830 52.340 114.000 52.510 ;
        RECT 114.360 52.340 114.530 52.510 ;
        RECT 114.720 52.340 114.890 52.510 ;
        RECT 115.080 52.340 115.250 52.510 ;
        RECT 115.920 52.340 116.090 52.510 ;
        RECT 116.280 52.340 116.450 52.510 ;
        RECT 116.640 52.340 116.810 52.510 ;
        RECT 117.480 52.340 117.650 52.510 ;
        RECT 117.840 52.340 118.010 52.510 ;
        RECT 118.200 52.340 118.370 52.510 ;
        RECT 119.790 52.350 119.960 52.520 ;
        RECT 120.230 52.350 120.400 52.520 ;
        RECT 120.640 52.350 120.810 52.520 ;
        RECT 121.070 52.350 121.240 52.520 ;
        RECT 121.510 52.350 121.680 52.520 ;
        RECT 121.920 52.350 122.090 52.520 ;
        RECT 124.160 52.340 124.330 52.510 ;
        RECT 124.520 52.340 124.690 52.510 ;
        RECT 124.880 52.340 125.050 52.510 ;
        RECT 125.240 52.340 125.410 52.510 ;
        RECT 125.600 52.340 125.770 52.510 ;
        RECT 126.460 52.340 126.630 52.510 ;
        RECT 126.820 52.340 126.990 52.510 ;
        RECT 128.860 52.340 129.030 52.510 ;
        RECT 129.300 52.340 129.470 52.510 ;
        RECT 129.740 52.340 129.910 52.510 ;
        RECT 130.150 52.340 130.320 52.510 ;
        RECT 130.680 52.340 130.850 52.510 ;
        RECT 131.040 52.340 131.210 52.510 ;
        RECT 131.400 52.340 131.570 52.510 ;
        RECT 132.240 52.340 132.410 52.510 ;
        RECT 132.600 52.340 132.770 52.510 ;
        RECT 132.960 52.340 133.130 52.510 ;
        RECT 133.800 52.340 133.970 52.510 ;
        RECT 134.160 52.340 134.330 52.510 ;
        RECT 134.520 52.340 134.690 52.510 ;
        RECT 135.580 52.340 135.750 52.510 ;
        RECT 136.020 52.340 136.190 52.510 ;
        RECT 136.460 52.340 136.630 52.510 ;
        RECT 136.870 52.340 137.040 52.510 ;
        RECT 137.390 52.340 137.560 52.510 ;
        RECT 137.750 52.340 137.920 52.510 ;
        RECT 138.110 52.340 138.280 52.510 ;
        RECT 139.030 52.340 139.200 52.510 ;
        RECT 139.390 52.340 139.560 52.510 ;
        RECT 139.900 52.340 140.070 52.510 ;
        RECT 140.340 52.340 140.510 52.510 ;
        RECT 140.780 52.340 140.950 52.510 ;
        RECT 141.190 52.340 141.360 52.510 ;
        RECT 5.920 44.680 6.090 44.860 ;
        RECT 6.400 44.680 6.570 44.860 ;
        RECT 6.880 44.680 7.050 44.860 ;
        RECT 7.360 44.680 7.530 44.860 ;
        RECT 7.840 44.680 8.010 44.860 ;
        RECT 8.320 44.680 8.490 44.860 ;
        RECT 8.800 44.680 8.970 44.860 ;
        RECT 9.280 44.680 9.450 44.860 ;
        RECT 9.760 44.680 9.930 44.860 ;
        RECT 10.240 44.680 10.410 44.860 ;
        RECT 10.720 44.680 10.890 44.860 ;
        RECT 11.200 44.680 11.370 44.860 ;
        RECT 11.680 44.680 11.850 44.860 ;
        RECT 12.160 44.680 12.330 44.860 ;
        RECT 12.640 44.680 12.810 44.860 ;
        RECT 13.120 44.680 13.290 44.860 ;
        RECT 13.600 44.680 13.770 44.860 ;
        RECT 14.080 44.680 14.250 44.860 ;
        RECT 14.560 44.680 14.730 44.860 ;
        RECT 15.040 44.680 15.210 44.860 ;
        RECT 15.520 44.680 15.690 44.860 ;
        RECT 16.000 44.680 16.170 44.860 ;
        RECT 16.480 44.680 16.650 44.860 ;
        RECT 16.960 44.680 17.130 44.860 ;
        RECT 17.440 44.680 17.610 44.860 ;
        RECT 17.920 44.680 18.090 44.860 ;
        RECT 18.400 44.680 18.570 44.860 ;
        RECT 18.880 44.680 19.050 44.860 ;
        RECT 19.360 44.680 19.530 44.860 ;
        RECT 19.840 44.680 20.010 44.860 ;
        RECT 20.320 44.680 20.490 44.860 ;
        RECT 20.800 44.680 20.970 44.860 ;
        RECT 21.280 44.680 21.450 44.860 ;
        RECT 21.760 44.680 21.930 44.860 ;
        RECT 22.240 44.680 22.410 44.860 ;
        RECT 22.720 44.680 22.890 44.860 ;
        RECT 23.200 44.680 23.370 44.860 ;
        RECT 23.680 44.680 23.850 44.860 ;
        RECT 24.160 44.680 24.330 44.860 ;
        RECT 24.640 44.680 24.810 44.860 ;
        RECT 25.120 44.680 25.290 44.860 ;
        RECT 25.600 44.680 25.770 44.860 ;
        RECT 26.080 44.680 26.250 44.860 ;
        RECT 26.560 44.680 26.730 44.860 ;
        RECT 27.040 44.680 27.210 44.860 ;
        RECT 27.520 44.680 27.690 44.860 ;
        RECT 28.000 44.680 28.170 44.860 ;
        RECT 28.480 44.680 28.650 44.860 ;
        RECT 28.960 44.680 29.130 44.860 ;
        RECT 29.440 44.680 29.610 44.860 ;
        RECT 29.920 44.680 30.090 44.860 ;
        RECT 30.400 44.680 30.570 44.860 ;
        RECT 30.880 44.680 31.050 44.860 ;
        RECT 31.360 44.680 31.530 44.860 ;
        RECT 31.840 44.680 32.010 44.860 ;
        RECT 32.320 44.680 32.490 44.860 ;
        RECT 32.800 44.680 32.970 44.860 ;
        RECT 33.280 44.680 33.450 44.860 ;
        RECT 33.760 44.680 33.930 44.860 ;
        RECT 34.240 44.680 34.410 44.860 ;
        RECT 34.720 44.680 34.890 44.860 ;
        RECT 35.200 44.680 35.370 44.860 ;
        RECT 35.680 44.680 35.850 44.860 ;
        RECT 36.160 44.680 36.330 44.860 ;
        RECT 36.640 44.680 36.810 44.860 ;
        RECT 37.120 44.680 37.290 44.860 ;
        RECT 37.600 44.680 37.770 44.860 ;
        RECT 38.080 44.680 38.250 44.860 ;
        RECT 38.560 44.680 38.730 44.860 ;
        RECT 39.040 44.680 39.210 44.860 ;
        RECT 39.520 44.680 39.690 44.860 ;
        RECT 40.000 44.680 40.170 44.860 ;
        RECT 40.480 44.680 40.650 44.860 ;
        RECT 40.960 44.680 41.130 44.860 ;
        RECT 41.440 44.680 41.610 44.860 ;
        RECT 41.920 44.680 42.090 44.860 ;
        RECT 42.400 44.680 42.570 44.860 ;
        RECT 42.880 44.680 43.050 44.860 ;
        RECT 43.360 44.680 43.530 44.860 ;
        RECT 43.840 44.680 44.010 44.860 ;
        RECT 44.320 44.680 44.490 44.860 ;
        RECT 44.800 44.680 44.970 44.860 ;
        RECT 45.280 44.680 45.450 44.860 ;
        RECT 45.760 44.680 45.930 44.860 ;
        RECT 46.240 44.680 46.410 44.860 ;
        RECT 46.720 44.680 46.890 44.860 ;
        RECT 47.200 44.680 47.370 44.860 ;
        RECT 47.680 44.680 47.850 44.860 ;
        RECT 48.160 44.680 48.330 44.860 ;
        RECT 48.640 44.680 48.810 44.860 ;
        RECT 49.120 44.680 49.290 44.860 ;
        RECT 49.600 44.680 49.770 44.860 ;
        RECT 50.080 44.680 50.250 44.860 ;
      LAYER li1 ;
        RECT 50.400 44.680 50.880 44.860 ;
      LAYER li1 ;
        RECT 51.040 44.680 51.210 44.860 ;
        RECT 51.520 44.680 51.690 44.860 ;
        RECT 52.000 44.680 52.170 44.860 ;
        RECT 52.480 44.680 52.650 44.860 ;
        RECT 52.960 44.680 53.130 44.860 ;
        RECT 53.440 44.680 53.610 44.860 ;
        RECT 53.920 44.680 54.090 44.860 ;
        RECT 54.400 44.680 54.570 44.860 ;
        RECT 54.880 44.680 55.050 44.860 ;
        RECT 55.360 44.680 55.530 44.860 ;
        RECT 55.840 44.680 56.010 44.860 ;
        RECT 56.320 44.680 56.490 44.860 ;
        RECT 56.800 44.680 56.970 44.860 ;
        RECT 57.280 44.680 57.450 44.860 ;
        RECT 57.760 44.680 57.930 44.860 ;
        RECT 58.240 44.680 58.410 44.860 ;
        RECT 58.720 44.680 58.890 44.860 ;
        RECT 59.200 44.680 59.370 44.860 ;
        RECT 59.680 44.680 59.850 44.860 ;
        RECT 60.160 44.680 60.330 44.860 ;
        RECT 60.640 44.680 60.810 44.860 ;
        RECT 61.120 44.680 61.290 44.860 ;
        RECT 61.600 44.680 61.770 44.860 ;
        RECT 62.080 44.680 62.250 44.860 ;
        RECT 62.560 44.680 62.730 44.860 ;
        RECT 63.040 44.680 63.210 44.860 ;
        RECT 63.520 44.680 63.690 44.860 ;
        RECT 64.000 44.680 64.170 44.860 ;
        RECT 64.480 44.680 64.650 44.860 ;
        RECT 64.960 44.680 65.130 44.860 ;
        RECT 65.440 44.680 65.610 44.860 ;
        RECT 65.920 44.680 66.090 44.860 ;
        RECT 66.400 44.680 66.570 44.860 ;
        RECT 66.880 44.680 67.050 44.860 ;
        RECT 67.360 44.680 67.530 44.860 ;
        RECT 67.840 44.680 68.010 44.860 ;
        RECT 68.320 44.680 68.490 44.860 ;
        RECT 68.800 44.680 68.970 44.860 ;
        RECT 69.280 44.680 69.450 44.860 ;
        RECT 69.760 44.680 69.930 44.860 ;
        RECT 70.240 44.680 70.410 44.860 ;
        RECT 70.720 44.680 70.890 44.860 ;
        RECT 71.200 44.680 71.370 44.860 ;
        RECT 71.680 44.680 71.850 44.860 ;
        RECT 72.160 44.680 72.330 44.860 ;
        RECT 72.640 44.680 72.810 44.860 ;
        RECT 73.120 44.680 73.290 44.860 ;
        RECT 73.600 44.680 73.770 44.860 ;
        RECT 74.080 44.680 74.250 44.860 ;
        RECT 74.560 44.680 74.730 44.860 ;
        RECT 75.040 44.680 75.210 44.860 ;
        RECT 75.520 44.680 75.690 44.860 ;
        RECT 76.000 44.680 76.170 44.860 ;
        RECT 76.480 44.680 76.650 44.860 ;
        RECT 76.960 44.680 77.130 44.860 ;
        RECT 77.440 44.680 77.610 44.860 ;
        RECT 77.920 44.680 78.090 44.860 ;
        RECT 78.400 44.680 78.570 44.860 ;
        RECT 78.880 44.680 79.050 44.860 ;
        RECT 79.360 44.680 79.530 44.860 ;
        RECT 79.840 44.680 80.010 44.860 ;
        RECT 80.320 44.680 80.490 44.860 ;
        RECT 80.800 44.680 80.970 44.860 ;
        RECT 81.280 44.680 81.450 44.860 ;
        RECT 81.760 44.680 81.930 44.860 ;
        RECT 82.240 44.680 82.410 44.860 ;
        RECT 82.720 44.680 82.890 44.860 ;
        RECT 83.200 44.680 83.370 44.860 ;
        RECT 83.680 44.680 83.850 44.860 ;
        RECT 84.160 44.680 84.330 44.860 ;
        RECT 84.640 44.680 84.810 44.860 ;
        RECT 85.120 44.680 85.290 44.860 ;
        RECT 85.600 44.680 85.770 44.860 ;
        RECT 86.080 44.680 86.250 44.860 ;
        RECT 86.560 44.680 86.730 44.860 ;
        RECT 87.040 44.680 87.210 44.860 ;
        RECT 87.520 44.680 87.690 44.860 ;
        RECT 88.000 44.680 88.170 44.860 ;
        RECT 88.480 44.680 88.650 44.860 ;
        RECT 88.960 44.680 89.130 44.860 ;
        RECT 89.440 44.680 89.610 44.860 ;
        RECT 89.920 44.680 90.090 44.860 ;
        RECT 90.400 44.680 90.570 44.860 ;
        RECT 90.880 44.680 91.050 44.860 ;
        RECT 91.360 44.680 91.530 44.860 ;
        RECT 91.840 44.680 92.010 44.860 ;
        RECT 92.320 44.680 92.490 44.860 ;
        RECT 92.800 44.680 92.970 44.860 ;
        RECT 93.280 44.680 93.450 44.860 ;
        RECT 93.760 44.680 93.930 44.860 ;
        RECT 94.240 44.680 94.410 44.860 ;
      LAYER li1 ;
        RECT 94.560 44.680 95.040 44.860 ;
      LAYER li1 ;
        RECT 95.200 44.680 95.370 44.860 ;
        RECT 95.680 44.680 95.850 44.860 ;
        RECT 96.160 44.680 96.330 44.860 ;
        RECT 96.640 44.680 96.810 44.860 ;
        RECT 97.120 44.680 97.290 44.860 ;
        RECT 97.600 44.680 97.770 44.860 ;
        RECT 98.080 44.680 98.250 44.860 ;
        RECT 98.560 44.680 98.730 44.860 ;
        RECT 99.040 44.680 99.210 44.860 ;
        RECT 99.520 44.680 99.690 44.860 ;
        RECT 100.000 44.680 100.170 44.860 ;
        RECT 100.480 44.680 100.650 44.860 ;
        RECT 100.960 44.680 101.130 44.860 ;
        RECT 101.440 44.680 101.610 44.860 ;
        RECT 101.920 44.680 102.090 44.860 ;
        RECT 102.400 44.680 102.570 44.860 ;
        RECT 102.880 44.680 103.050 44.860 ;
        RECT 103.360 44.680 103.530 44.860 ;
        RECT 103.840 44.680 104.010 44.860 ;
        RECT 104.320 44.680 104.490 44.860 ;
        RECT 104.800 44.680 104.970 44.860 ;
        RECT 105.280 44.680 105.450 44.860 ;
        RECT 105.760 44.680 105.930 44.860 ;
        RECT 106.240 44.680 106.410 44.860 ;
        RECT 106.720 44.680 106.890 44.860 ;
        RECT 107.200 44.680 107.370 44.860 ;
        RECT 107.680 44.680 107.850 44.860 ;
      LAYER li1 ;
        RECT 108.000 44.680 108.480 44.860 ;
      LAYER li1 ;
        RECT 108.640 44.680 108.810 44.860 ;
        RECT 109.120 44.680 109.290 44.860 ;
        RECT 109.600 44.680 109.770 44.860 ;
        RECT 110.080 44.680 110.250 44.860 ;
        RECT 110.560 44.680 110.730 44.860 ;
        RECT 111.040 44.680 111.210 44.860 ;
        RECT 111.520 44.680 111.690 44.860 ;
        RECT 112.000 44.680 112.170 44.860 ;
        RECT 112.480 44.680 112.650 44.860 ;
        RECT 112.960 44.680 113.130 44.860 ;
        RECT 113.440 44.680 113.610 44.860 ;
        RECT 113.920 44.680 114.090 44.860 ;
        RECT 114.400 44.680 114.570 44.860 ;
        RECT 114.880 44.680 115.050 44.860 ;
        RECT 115.360 44.680 115.530 44.860 ;
        RECT 115.840 44.680 116.010 44.860 ;
        RECT 116.320 44.680 116.490 44.860 ;
        RECT 116.800 44.680 116.970 44.860 ;
        RECT 117.280 44.680 117.450 44.860 ;
        RECT 117.760 44.680 117.930 44.860 ;
        RECT 118.240 44.680 118.410 44.860 ;
        RECT 118.720 44.680 118.890 44.860 ;
        RECT 119.200 44.680 119.370 44.860 ;
        RECT 119.680 44.680 119.850 44.860 ;
        RECT 120.160 44.680 120.330 44.860 ;
        RECT 120.640 44.680 120.810 44.860 ;
        RECT 121.120 44.680 121.290 44.860 ;
        RECT 121.600 44.680 121.770 44.860 ;
        RECT 122.080 44.680 122.250 44.860 ;
        RECT 122.560 44.680 122.730 44.860 ;
        RECT 123.040 44.680 123.210 44.860 ;
        RECT 123.520 44.680 123.690 44.860 ;
        RECT 124.000 44.680 124.170 44.860 ;
        RECT 124.480 44.680 124.650 44.860 ;
        RECT 124.960 44.680 125.130 44.860 ;
        RECT 125.440 44.680 125.610 44.860 ;
        RECT 125.920 44.680 126.090 44.860 ;
        RECT 126.400 44.680 126.570 44.860 ;
        RECT 126.880 44.680 127.050 44.860 ;
        RECT 127.360 44.680 127.530 44.860 ;
        RECT 127.840 44.680 128.010 44.860 ;
        RECT 128.320 44.680 128.490 44.860 ;
        RECT 128.800 44.680 128.970 44.860 ;
        RECT 129.280 44.680 129.450 44.860 ;
        RECT 129.760 44.680 129.930 44.860 ;
        RECT 130.240 44.680 130.410 44.860 ;
        RECT 130.720 44.680 130.890 44.860 ;
        RECT 131.200 44.680 131.370 44.860 ;
        RECT 131.680 44.680 131.850 44.860 ;
        RECT 132.160 44.680 132.330 44.860 ;
        RECT 132.640 44.680 132.810 44.860 ;
        RECT 133.120 44.680 133.290 44.860 ;
        RECT 133.600 44.680 133.770 44.860 ;
        RECT 134.080 44.680 134.250 44.860 ;
        RECT 134.560 44.680 134.730 44.860 ;
        RECT 135.040 44.680 135.210 44.860 ;
        RECT 135.520 44.680 135.690 44.860 ;
        RECT 136.000 44.680 136.170 44.860 ;
        RECT 136.480 44.680 136.650 44.860 ;
        RECT 136.960 44.680 137.130 44.860 ;
        RECT 137.440 44.680 137.610 44.860 ;
        RECT 137.920 44.680 138.090 44.860 ;
        RECT 138.400 44.680 138.570 44.860 ;
        RECT 138.880 44.680 139.050 44.860 ;
        RECT 139.360 44.680 139.530 44.860 ;
        RECT 139.840 44.680 140.010 44.860 ;
        RECT 140.320 44.680 140.490 44.860 ;
        RECT 140.800 44.680 140.970 44.860 ;
        RECT 141.280 44.680 141.450 44.860 ;
        RECT 141.760 44.680 141.930 44.860 ;
        RECT 6.510 44.210 6.680 44.380 ;
        RECT 6.950 44.210 7.120 44.380 ;
        RECT 7.360 44.210 7.530 44.380 ;
        RECT 7.790 44.210 7.960 44.380 ;
        RECT 8.230 44.210 8.400 44.380 ;
        RECT 8.640 44.210 8.810 44.380 ;
        RECT 9.820 44.200 9.990 44.370 ;
        RECT 10.260 44.200 10.430 44.370 ;
        RECT 10.700 44.200 10.870 44.370 ;
        RECT 11.110 44.200 11.280 44.370 ;
        RECT 12.600 44.200 12.770 44.370 ;
        RECT 12.960 44.200 13.130 44.370 ;
        RECT 14.140 44.200 14.310 44.370 ;
        RECT 14.580 44.200 14.750 44.370 ;
        RECT 15.020 44.200 15.190 44.370 ;
        RECT 15.430 44.200 15.600 44.370 ;
        RECT 16.390 44.200 16.560 44.370 ;
        RECT 16.750 44.200 16.920 44.370 ;
        RECT 17.110 44.200 17.280 44.370 ;
        RECT 17.470 44.200 17.640 44.370 ;
        RECT 18.460 44.200 18.630 44.370 ;
        RECT 18.900 44.200 19.070 44.370 ;
        RECT 19.340 44.200 19.510 44.370 ;
        RECT 19.750 44.200 19.920 44.370 ;
        RECT 20.800 44.200 20.970 44.370 ;
        RECT 21.160 44.200 21.330 44.370 ;
        RECT 21.520 44.200 21.690 44.370 ;
        RECT 23.740 44.200 23.910 44.370 ;
        RECT 24.180 44.200 24.350 44.370 ;
        RECT 24.620 44.200 24.790 44.370 ;
        RECT 25.030 44.200 25.200 44.370 ;
        RECT 26.080 44.200 26.250 44.370 ;
        RECT 26.440 44.200 26.610 44.370 ;
        RECT 26.800 44.200 26.970 44.370 ;
        RECT 29.020 44.200 29.190 44.370 ;
        RECT 29.460 44.200 29.630 44.370 ;
        RECT 29.900 44.200 30.070 44.370 ;
        RECT 30.310 44.200 30.480 44.370 ;
        RECT 30.840 44.200 31.010 44.370 ;
        RECT 31.200 44.200 31.370 44.370 ;
        RECT 31.560 44.200 31.730 44.370 ;
        RECT 32.400 44.200 32.570 44.370 ;
        RECT 32.760 44.200 32.930 44.370 ;
        RECT 33.120 44.200 33.290 44.370 ;
        RECT 33.960 44.200 34.130 44.370 ;
        RECT 34.320 44.200 34.490 44.370 ;
        RECT 34.680 44.200 34.850 44.370 ;
        RECT 35.740 44.200 35.910 44.370 ;
        RECT 36.180 44.200 36.350 44.370 ;
        RECT 36.620 44.200 36.790 44.370 ;
        RECT 37.030 44.200 37.200 44.370 ;
        RECT 37.560 44.200 37.730 44.370 ;
        RECT 37.920 44.200 38.090 44.370 ;
        RECT 39.100 44.200 39.270 44.370 ;
        RECT 39.540 44.200 39.710 44.370 ;
        RECT 39.980 44.200 40.150 44.370 ;
        RECT 40.390 44.200 40.560 44.370 ;
        RECT 40.920 44.200 41.090 44.370 ;
        RECT 41.280 44.200 41.450 44.370 ;
        RECT 41.640 44.200 41.810 44.370 ;
        RECT 42.480 44.200 42.650 44.370 ;
        RECT 42.840 44.200 43.010 44.370 ;
        RECT 43.200 44.200 43.370 44.370 ;
        RECT 44.040 44.200 44.210 44.370 ;
        RECT 44.400 44.200 44.570 44.370 ;
        RECT 44.760 44.200 44.930 44.370 ;
        RECT 45.820 44.200 45.990 44.370 ;
        RECT 46.260 44.200 46.430 44.370 ;
        RECT 46.700 44.200 46.870 44.370 ;
        RECT 47.110 44.200 47.280 44.370 ;
        RECT 47.640 44.200 47.810 44.370 ;
        RECT 48.000 44.200 48.170 44.370 ;
        RECT 48.360 44.200 48.530 44.370 ;
        RECT 49.200 44.200 49.370 44.370 ;
        RECT 49.560 44.200 49.730 44.370 ;
        RECT 49.920 44.200 50.090 44.370 ;
        RECT 50.760 44.200 50.930 44.370 ;
        RECT 51.120 44.200 51.290 44.370 ;
        RECT 51.480 44.200 51.650 44.370 ;
        RECT 52.540 44.200 52.710 44.370 ;
        RECT 52.980 44.200 53.150 44.370 ;
        RECT 53.420 44.200 53.590 44.370 ;
        RECT 53.830 44.200 54.000 44.370 ;
        RECT 54.360 44.200 54.530 44.370 ;
        RECT 54.720 44.200 54.890 44.370 ;
        RECT 55.080 44.200 55.250 44.370 ;
        RECT 55.920 44.200 56.090 44.370 ;
        RECT 56.280 44.200 56.450 44.370 ;
        RECT 56.640 44.200 56.810 44.370 ;
        RECT 57.480 44.200 57.650 44.370 ;
        RECT 57.840 44.200 58.010 44.370 ;
        RECT 58.200 44.200 58.370 44.370 ;
        RECT 59.260 44.200 59.430 44.370 ;
        RECT 59.700 44.200 59.870 44.370 ;
        RECT 60.140 44.200 60.310 44.370 ;
        RECT 60.550 44.200 60.720 44.370 ;
        RECT 61.080 44.200 61.250 44.370 ;
        RECT 61.440 44.200 61.610 44.370 ;
        RECT 61.800 44.200 61.970 44.370 ;
        RECT 62.640 44.200 62.810 44.370 ;
        RECT 63.000 44.200 63.170 44.370 ;
        RECT 63.360 44.200 63.530 44.370 ;
        RECT 64.200 44.200 64.370 44.370 ;
        RECT 64.560 44.200 64.730 44.370 ;
        RECT 64.920 44.200 65.090 44.370 ;
        RECT 65.980 44.200 66.150 44.370 ;
        RECT 66.420 44.200 66.590 44.370 ;
        RECT 66.860 44.200 67.030 44.370 ;
        RECT 67.270 44.200 67.440 44.370 ;
        RECT 67.800 44.200 67.970 44.370 ;
        RECT 68.160 44.200 68.330 44.370 ;
        RECT 68.520 44.200 68.690 44.370 ;
        RECT 69.360 44.200 69.530 44.370 ;
        RECT 69.720 44.200 69.890 44.370 ;
        RECT 70.080 44.200 70.250 44.370 ;
        RECT 70.920 44.200 71.090 44.370 ;
        RECT 71.280 44.200 71.450 44.370 ;
        RECT 71.640 44.200 71.810 44.370 ;
        RECT 72.700 44.200 72.870 44.370 ;
        RECT 73.140 44.200 73.310 44.370 ;
        RECT 73.580 44.200 73.750 44.370 ;
        RECT 73.990 44.200 74.160 44.370 ;
        RECT 74.520 44.200 74.690 44.370 ;
        RECT 74.880 44.200 75.050 44.370 ;
        RECT 75.240 44.200 75.410 44.370 ;
        RECT 76.080 44.200 76.250 44.370 ;
        RECT 76.440 44.200 76.610 44.370 ;
        RECT 76.800 44.200 76.970 44.370 ;
        RECT 77.640 44.200 77.810 44.370 ;
        RECT 78.000 44.200 78.170 44.370 ;
        RECT 78.360 44.200 78.530 44.370 ;
        RECT 79.420 44.200 79.590 44.370 ;
        RECT 79.860 44.200 80.030 44.370 ;
        RECT 80.300 44.200 80.470 44.370 ;
        RECT 80.710 44.200 80.880 44.370 ;
        RECT 81.240 44.200 81.410 44.370 ;
        RECT 81.600 44.200 81.770 44.370 ;
        RECT 81.960 44.200 82.130 44.370 ;
        RECT 82.800 44.200 82.970 44.370 ;
        RECT 83.160 44.200 83.330 44.370 ;
        RECT 83.520 44.200 83.690 44.370 ;
        RECT 84.360 44.200 84.530 44.370 ;
        RECT 84.720 44.200 84.890 44.370 ;
        RECT 85.080 44.200 85.250 44.370 ;
        RECT 86.140 44.200 86.310 44.370 ;
        RECT 86.580 44.200 86.750 44.370 ;
        RECT 87.020 44.200 87.190 44.370 ;
        RECT 87.430 44.200 87.600 44.370 ;
        RECT 87.960 44.200 88.130 44.370 ;
        RECT 88.320 44.200 88.490 44.370 ;
        RECT 88.680 44.200 88.850 44.370 ;
        RECT 89.520 44.200 89.690 44.370 ;
        RECT 89.880 44.200 90.050 44.370 ;
        RECT 90.240 44.200 90.410 44.370 ;
        RECT 91.080 44.200 91.250 44.370 ;
        RECT 91.440 44.200 91.610 44.370 ;
        RECT 91.800 44.200 91.970 44.370 ;
        RECT 92.860 44.200 93.030 44.370 ;
        RECT 93.300 44.200 93.470 44.370 ;
        RECT 93.740 44.200 93.910 44.370 ;
        RECT 94.150 44.200 94.320 44.370 ;
        RECT 96.760 44.200 96.930 44.370 ;
        RECT 97.120 44.200 97.290 44.370 ;
        RECT 97.480 44.200 97.650 44.370 ;
        RECT 98.620 44.200 98.790 44.370 ;
        RECT 99.060 44.200 99.230 44.370 ;
        RECT 99.500 44.200 99.670 44.370 ;
        RECT 99.910 44.200 100.080 44.370 ;
        RECT 101.400 44.200 101.570 44.370 ;
        RECT 101.760 44.200 101.930 44.370 ;
        RECT 102.120 44.200 102.290 44.370 ;
        RECT 102.960 44.200 103.130 44.370 ;
        RECT 103.320 44.200 103.490 44.370 ;
        RECT 103.680 44.200 103.850 44.370 ;
        RECT 104.520 44.200 104.690 44.370 ;
        RECT 104.880 44.200 105.050 44.370 ;
        RECT 105.240 44.200 105.410 44.370 ;
        RECT 106.300 44.200 106.470 44.370 ;
        RECT 106.740 44.200 106.910 44.370 ;
        RECT 107.180 44.200 107.350 44.370 ;
        RECT 107.590 44.200 107.760 44.370 ;
        RECT 108.120 44.200 108.290 44.370 ;
        RECT 108.480 44.200 108.650 44.370 ;
        RECT 108.840 44.200 109.010 44.370 ;
        RECT 109.680 44.200 109.850 44.370 ;
        RECT 110.040 44.200 110.210 44.370 ;
        RECT 110.400 44.200 110.570 44.370 ;
        RECT 111.240 44.200 111.410 44.370 ;
        RECT 111.600 44.200 111.770 44.370 ;
        RECT 111.960 44.200 112.130 44.370 ;
        RECT 113.020 44.200 113.190 44.370 ;
        RECT 113.460 44.200 113.630 44.370 ;
        RECT 113.900 44.200 114.070 44.370 ;
        RECT 114.310 44.200 114.480 44.370 ;
        RECT 116.280 44.200 116.450 44.370 ;
        RECT 116.640 44.200 116.810 44.370 ;
        RECT 117.000 44.200 117.170 44.370 ;
        RECT 117.840 44.200 118.010 44.370 ;
        RECT 118.200 44.200 118.370 44.370 ;
        RECT 118.560 44.200 118.730 44.370 ;
        RECT 119.400 44.200 119.570 44.370 ;
        RECT 119.760 44.200 119.930 44.370 ;
        RECT 120.120 44.200 120.290 44.370 ;
        RECT 121.180 44.200 121.350 44.370 ;
        RECT 121.620 44.200 121.790 44.370 ;
        RECT 122.060 44.200 122.230 44.370 ;
        RECT 122.470 44.200 122.640 44.370 ;
        RECT 123.000 44.200 123.170 44.370 ;
        RECT 123.360 44.200 123.530 44.370 ;
        RECT 123.720 44.200 123.890 44.370 ;
        RECT 124.560 44.200 124.730 44.370 ;
        RECT 124.920 44.200 125.090 44.370 ;
        RECT 125.280 44.200 125.450 44.370 ;
        RECT 126.120 44.200 126.290 44.370 ;
        RECT 126.480 44.200 126.650 44.370 ;
        RECT 126.840 44.200 127.010 44.370 ;
        RECT 127.900 44.200 128.070 44.370 ;
        RECT 128.340 44.200 128.510 44.370 ;
        RECT 128.780 44.200 128.950 44.370 ;
        RECT 129.190 44.200 129.360 44.370 ;
        RECT 129.720 44.200 129.890 44.370 ;
        RECT 130.080 44.200 130.250 44.370 ;
        RECT 130.440 44.200 130.610 44.370 ;
        RECT 131.280 44.200 131.450 44.370 ;
        RECT 131.640 44.200 131.810 44.370 ;
        RECT 132.000 44.200 132.170 44.370 ;
        RECT 132.840 44.200 133.010 44.370 ;
        RECT 133.200 44.200 133.370 44.370 ;
        RECT 133.560 44.200 133.730 44.370 ;
        RECT 134.620 44.200 134.790 44.370 ;
        RECT 135.060 44.200 135.230 44.370 ;
        RECT 135.500 44.200 135.670 44.370 ;
        RECT 135.910 44.200 136.080 44.370 ;
        RECT 136.700 44.200 136.870 44.370 ;
        RECT 137.060 44.200 137.230 44.370 ;
        RECT 137.420 44.200 137.590 44.370 ;
        RECT 137.780 44.200 137.950 44.370 ;
        RECT 138.140 44.200 138.310 44.370 ;
        RECT 139.030 44.200 139.200 44.370 ;
        RECT 139.390 44.200 139.560 44.370 ;
        RECT 139.900 44.200 140.070 44.370 ;
        RECT 140.340 44.200 140.510 44.370 ;
        RECT 140.780 44.200 140.950 44.370 ;
        RECT 141.190 44.200 141.360 44.370 ;
        RECT 5.920 36.540 6.090 36.720 ;
        RECT 6.400 36.540 6.570 36.720 ;
        RECT 6.880 36.540 7.050 36.720 ;
        RECT 7.360 36.540 7.530 36.720 ;
        RECT 7.840 36.540 8.010 36.720 ;
        RECT 8.320 36.540 8.490 36.720 ;
        RECT 8.800 36.540 8.970 36.720 ;
        RECT 9.280 36.540 9.450 36.720 ;
        RECT 9.760 36.540 9.930 36.720 ;
        RECT 10.240 36.540 10.410 36.720 ;
        RECT 10.720 36.540 10.890 36.720 ;
        RECT 11.200 36.540 11.370 36.720 ;
        RECT 11.680 36.540 11.850 36.720 ;
        RECT 12.160 36.540 12.330 36.720 ;
        RECT 12.640 36.540 12.810 36.720 ;
        RECT 13.120 36.540 13.290 36.720 ;
        RECT 13.600 36.540 13.770 36.720 ;
        RECT 14.080 36.540 14.250 36.720 ;
      LAYER li1 ;
        RECT 14.400 36.540 14.880 36.720 ;
      LAYER li1 ;
        RECT 15.040 36.540 15.210 36.720 ;
        RECT 15.520 36.540 15.690 36.720 ;
        RECT 16.000 36.540 16.170 36.720 ;
        RECT 16.480 36.540 16.650 36.720 ;
        RECT 16.960 36.540 17.130 36.720 ;
        RECT 17.440 36.540 17.610 36.720 ;
        RECT 17.920 36.540 18.090 36.720 ;
        RECT 18.400 36.540 18.570 36.720 ;
        RECT 18.880 36.540 19.050 36.720 ;
        RECT 19.360 36.540 19.530 36.720 ;
        RECT 19.840 36.540 20.010 36.720 ;
        RECT 20.320 36.540 20.490 36.720 ;
        RECT 20.800 36.540 20.970 36.720 ;
        RECT 21.280 36.540 21.450 36.720 ;
        RECT 21.760 36.540 21.930 36.720 ;
        RECT 22.240 36.540 22.410 36.720 ;
        RECT 22.720 36.540 22.890 36.720 ;
        RECT 23.200 36.540 23.370 36.720 ;
        RECT 23.680 36.540 23.850 36.720 ;
        RECT 24.160 36.540 24.330 36.720 ;
        RECT 24.640 36.540 24.810 36.720 ;
        RECT 25.120 36.540 25.290 36.720 ;
        RECT 25.600 36.540 25.770 36.720 ;
        RECT 26.080 36.540 26.250 36.720 ;
        RECT 26.560 36.540 26.730 36.720 ;
        RECT 27.040 36.540 27.210 36.720 ;
        RECT 27.520 36.540 27.690 36.720 ;
        RECT 28.000 36.540 28.170 36.720 ;
        RECT 28.480 36.540 28.650 36.720 ;
        RECT 28.960 36.540 29.130 36.720 ;
        RECT 29.440 36.540 29.610 36.720 ;
        RECT 29.920 36.540 30.090 36.720 ;
        RECT 30.400 36.540 30.570 36.720 ;
        RECT 30.880 36.540 31.050 36.720 ;
        RECT 31.360 36.540 31.530 36.720 ;
        RECT 31.840 36.540 32.010 36.720 ;
        RECT 32.320 36.540 32.490 36.720 ;
        RECT 32.800 36.540 32.970 36.720 ;
        RECT 33.280 36.540 33.450 36.720 ;
        RECT 33.760 36.540 33.930 36.720 ;
        RECT 34.240 36.540 34.410 36.720 ;
        RECT 34.720 36.540 34.890 36.720 ;
        RECT 35.200 36.540 35.370 36.720 ;
        RECT 35.680 36.540 35.850 36.720 ;
        RECT 36.160 36.540 36.330 36.720 ;
        RECT 36.640 36.540 36.810 36.720 ;
        RECT 37.120 36.540 37.290 36.720 ;
        RECT 37.600 36.540 37.770 36.720 ;
        RECT 38.080 36.540 38.250 36.720 ;
        RECT 38.560 36.540 38.730 36.720 ;
        RECT 39.040 36.540 39.210 36.720 ;
        RECT 39.520 36.540 39.690 36.720 ;
        RECT 40.000 36.540 40.170 36.720 ;
        RECT 40.480 36.540 40.650 36.720 ;
        RECT 40.960 36.540 41.130 36.720 ;
        RECT 41.440 36.540 41.610 36.720 ;
        RECT 41.920 36.540 42.090 36.720 ;
        RECT 42.400 36.540 42.570 36.720 ;
        RECT 42.880 36.540 43.050 36.720 ;
        RECT 43.360 36.540 43.530 36.720 ;
        RECT 43.840 36.540 44.010 36.720 ;
        RECT 44.320 36.540 44.490 36.720 ;
        RECT 44.800 36.540 44.970 36.720 ;
        RECT 45.280 36.540 45.450 36.720 ;
        RECT 45.760 36.540 45.930 36.720 ;
        RECT 46.240 36.540 46.410 36.720 ;
        RECT 46.720 36.540 46.890 36.720 ;
        RECT 47.200 36.540 47.370 36.720 ;
        RECT 47.680 36.540 47.850 36.720 ;
        RECT 48.160 36.540 48.330 36.720 ;
        RECT 48.640 36.540 48.810 36.720 ;
        RECT 49.120 36.540 49.290 36.720 ;
        RECT 49.600 36.540 49.770 36.720 ;
        RECT 50.080 36.540 50.250 36.720 ;
        RECT 50.560 36.540 50.730 36.720 ;
        RECT 51.040 36.540 51.210 36.720 ;
        RECT 51.520 36.540 51.690 36.720 ;
        RECT 52.000 36.540 52.170 36.720 ;
        RECT 52.480 36.540 52.650 36.720 ;
        RECT 52.960 36.540 53.130 36.720 ;
        RECT 53.440 36.540 53.610 36.720 ;
        RECT 53.920 36.540 54.090 36.720 ;
        RECT 54.400 36.540 54.570 36.720 ;
        RECT 54.880 36.540 55.050 36.720 ;
        RECT 55.360 36.540 55.530 36.720 ;
        RECT 55.840 36.540 56.010 36.720 ;
        RECT 56.320 36.540 56.490 36.720 ;
        RECT 56.800 36.540 56.970 36.720 ;
        RECT 57.280 36.540 57.450 36.720 ;
        RECT 57.760 36.540 57.930 36.720 ;
        RECT 58.240 36.540 58.410 36.720 ;
        RECT 58.720 36.540 58.890 36.720 ;
        RECT 59.200 36.540 59.370 36.720 ;
        RECT 59.680 36.540 59.850 36.720 ;
        RECT 60.160 36.540 60.330 36.720 ;
        RECT 60.640 36.540 60.810 36.720 ;
        RECT 61.120 36.540 61.290 36.720 ;
        RECT 61.600 36.540 61.770 36.720 ;
        RECT 62.080 36.540 62.250 36.720 ;
        RECT 62.560 36.540 62.730 36.720 ;
        RECT 63.040 36.540 63.210 36.720 ;
        RECT 63.520 36.540 63.690 36.720 ;
        RECT 64.000 36.540 64.170 36.720 ;
        RECT 64.480 36.540 64.650 36.720 ;
        RECT 64.960 36.540 65.130 36.720 ;
        RECT 65.440 36.540 65.610 36.720 ;
        RECT 65.920 36.540 66.090 36.720 ;
        RECT 66.400 36.540 66.570 36.720 ;
        RECT 66.880 36.540 67.050 36.720 ;
        RECT 67.360 36.540 67.530 36.720 ;
        RECT 67.840 36.540 68.010 36.720 ;
        RECT 68.320 36.540 68.490 36.720 ;
        RECT 68.800 36.540 68.970 36.720 ;
        RECT 69.280 36.540 69.450 36.720 ;
        RECT 69.760 36.540 69.930 36.720 ;
        RECT 70.240 36.540 70.410 36.720 ;
        RECT 70.720 36.540 70.890 36.720 ;
        RECT 71.200 36.540 71.370 36.720 ;
        RECT 71.680 36.540 71.850 36.720 ;
        RECT 72.160 36.540 72.330 36.720 ;
        RECT 72.640 36.540 72.810 36.720 ;
        RECT 73.120 36.540 73.290 36.720 ;
        RECT 73.600 36.540 73.770 36.720 ;
        RECT 74.080 36.540 74.250 36.720 ;
        RECT 74.560 36.540 74.730 36.720 ;
        RECT 75.040 36.540 75.210 36.720 ;
        RECT 75.520 36.540 75.690 36.720 ;
        RECT 76.000 36.540 76.170 36.720 ;
        RECT 76.480 36.540 76.650 36.720 ;
        RECT 76.960 36.540 77.130 36.720 ;
        RECT 77.440 36.540 77.610 36.720 ;
      LAYER li1 ;
        RECT 77.760 36.540 78.240 36.720 ;
      LAYER li1 ;
        RECT 78.400 36.540 78.570 36.720 ;
        RECT 78.880 36.540 79.050 36.720 ;
        RECT 79.360 36.540 79.530 36.720 ;
        RECT 79.840 36.540 80.010 36.720 ;
        RECT 80.320 36.540 80.490 36.720 ;
        RECT 80.800 36.540 80.970 36.720 ;
        RECT 81.280 36.540 81.450 36.720 ;
        RECT 81.760 36.540 81.930 36.720 ;
        RECT 82.240 36.540 82.410 36.720 ;
        RECT 82.720 36.540 82.890 36.720 ;
        RECT 83.200 36.540 83.370 36.720 ;
        RECT 83.680 36.540 83.850 36.720 ;
        RECT 84.160 36.540 84.330 36.720 ;
        RECT 84.640 36.540 84.810 36.720 ;
        RECT 85.120 36.540 85.290 36.720 ;
        RECT 85.600 36.540 85.770 36.720 ;
        RECT 86.080 36.540 86.250 36.720 ;
        RECT 86.560 36.540 86.730 36.720 ;
        RECT 87.040 36.540 87.210 36.720 ;
        RECT 87.520 36.540 87.690 36.720 ;
        RECT 88.000 36.540 88.170 36.720 ;
        RECT 88.480 36.540 88.650 36.720 ;
        RECT 88.960 36.540 89.130 36.720 ;
        RECT 89.440 36.540 89.610 36.720 ;
        RECT 89.920 36.540 90.090 36.720 ;
        RECT 90.400 36.540 90.570 36.720 ;
        RECT 90.880 36.540 91.050 36.720 ;
        RECT 91.360 36.540 91.530 36.720 ;
        RECT 91.840 36.540 92.010 36.720 ;
        RECT 92.320 36.540 92.490 36.720 ;
        RECT 92.800 36.540 92.970 36.720 ;
        RECT 93.280 36.540 93.450 36.720 ;
        RECT 93.760 36.540 93.930 36.720 ;
        RECT 94.240 36.540 94.410 36.720 ;
        RECT 94.720 36.540 94.890 36.720 ;
        RECT 95.200 36.540 95.370 36.720 ;
        RECT 95.680 36.540 95.850 36.720 ;
        RECT 96.160 36.540 96.330 36.720 ;
        RECT 96.640 36.540 96.810 36.720 ;
        RECT 97.120 36.540 97.290 36.720 ;
        RECT 97.600 36.540 97.770 36.720 ;
        RECT 98.080 36.540 98.250 36.720 ;
        RECT 98.560 36.540 98.730 36.720 ;
        RECT 99.040 36.540 99.210 36.720 ;
        RECT 99.520 36.540 99.690 36.720 ;
        RECT 100.000 36.540 100.170 36.720 ;
        RECT 100.480 36.540 100.650 36.720 ;
        RECT 100.960 36.540 101.130 36.720 ;
        RECT 101.440 36.540 101.610 36.720 ;
        RECT 101.920 36.540 102.090 36.720 ;
        RECT 102.400 36.540 102.570 36.720 ;
        RECT 102.880 36.540 103.050 36.720 ;
        RECT 103.360 36.540 103.530 36.720 ;
        RECT 103.840 36.540 104.010 36.720 ;
        RECT 104.320 36.540 104.490 36.720 ;
        RECT 104.800 36.540 104.970 36.720 ;
        RECT 105.280 36.540 105.450 36.720 ;
        RECT 105.760 36.540 105.930 36.720 ;
        RECT 106.240 36.540 106.410 36.720 ;
        RECT 106.720 36.540 106.890 36.720 ;
        RECT 107.200 36.540 107.370 36.720 ;
        RECT 107.680 36.540 107.850 36.720 ;
        RECT 108.160 36.540 108.330 36.720 ;
        RECT 108.640 36.540 108.810 36.720 ;
        RECT 109.120 36.540 109.290 36.720 ;
        RECT 109.600 36.540 109.770 36.720 ;
        RECT 110.080 36.540 110.250 36.720 ;
      LAYER li1 ;
        RECT 110.400 36.540 110.880 36.720 ;
      LAYER li1 ;
        RECT 111.040 36.540 111.210 36.720 ;
        RECT 111.520 36.540 111.690 36.720 ;
        RECT 112.000 36.540 112.170 36.720 ;
        RECT 112.480 36.540 112.650 36.720 ;
        RECT 112.960 36.540 113.130 36.720 ;
        RECT 113.440 36.540 113.610 36.720 ;
        RECT 113.920 36.540 114.090 36.720 ;
        RECT 114.400 36.540 114.570 36.720 ;
        RECT 114.880 36.540 115.050 36.720 ;
        RECT 115.360 36.540 115.530 36.720 ;
        RECT 115.840 36.540 116.010 36.720 ;
        RECT 116.320 36.540 116.490 36.720 ;
        RECT 116.800 36.540 116.970 36.720 ;
        RECT 117.280 36.540 117.450 36.720 ;
        RECT 117.760 36.540 117.930 36.720 ;
        RECT 118.240 36.540 118.410 36.720 ;
        RECT 118.720 36.540 118.890 36.720 ;
        RECT 119.200 36.540 119.370 36.720 ;
        RECT 119.680 36.540 119.850 36.720 ;
        RECT 120.160 36.540 120.330 36.720 ;
        RECT 120.640 36.540 120.810 36.720 ;
        RECT 121.120 36.540 121.290 36.720 ;
        RECT 121.600 36.540 121.770 36.720 ;
        RECT 122.080 36.540 122.250 36.720 ;
        RECT 122.560 36.540 122.730 36.720 ;
        RECT 123.040 36.540 123.210 36.720 ;
        RECT 123.520 36.540 123.690 36.720 ;
        RECT 124.000 36.540 124.170 36.720 ;
        RECT 124.480 36.540 124.650 36.720 ;
        RECT 124.960 36.540 125.130 36.720 ;
        RECT 125.440 36.540 125.610 36.720 ;
        RECT 125.920 36.540 126.090 36.720 ;
        RECT 126.400 36.540 126.570 36.720 ;
        RECT 126.880 36.540 127.050 36.720 ;
        RECT 127.360 36.540 127.530 36.720 ;
        RECT 127.840 36.540 128.010 36.720 ;
        RECT 128.320 36.540 128.490 36.720 ;
        RECT 128.800 36.540 128.970 36.720 ;
        RECT 129.280 36.540 129.450 36.720 ;
        RECT 129.760 36.540 129.930 36.720 ;
        RECT 130.240 36.540 130.410 36.720 ;
        RECT 130.720 36.540 130.890 36.720 ;
        RECT 131.200 36.540 131.370 36.720 ;
        RECT 131.680 36.540 131.850 36.720 ;
        RECT 132.160 36.540 132.330 36.720 ;
        RECT 132.640 36.540 132.810 36.720 ;
        RECT 133.120 36.540 133.290 36.720 ;
        RECT 133.600 36.540 133.770 36.720 ;
        RECT 134.080 36.540 134.250 36.720 ;
        RECT 134.560 36.540 134.730 36.720 ;
        RECT 135.040 36.540 135.210 36.720 ;
        RECT 135.520 36.540 135.690 36.720 ;
        RECT 136.000 36.540 136.170 36.720 ;
        RECT 136.480 36.540 136.650 36.720 ;
        RECT 136.960 36.540 137.130 36.720 ;
        RECT 137.440 36.540 137.610 36.720 ;
        RECT 137.920 36.540 138.090 36.720 ;
        RECT 138.400 36.540 138.570 36.720 ;
        RECT 138.880 36.540 139.050 36.720 ;
        RECT 139.360 36.540 139.530 36.720 ;
        RECT 139.840 36.540 140.010 36.720 ;
        RECT 140.320 36.540 140.490 36.720 ;
        RECT 140.800 36.540 140.970 36.720 ;
        RECT 141.280 36.540 141.450 36.720 ;
        RECT 141.760 36.540 141.930 36.720 ;
        RECT 6.510 36.070 6.680 36.240 ;
        RECT 6.950 36.070 7.120 36.240 ;
        RECT 7.360 36.070 7.530 36.240 ;
        RECT 7.790 36.070 7.960 36.240 ;
        RECT 8.230 36.070 8.400 36.240 ;
        RECT 8.640 36.070 8.810 36.240 ;
        RECT 10.680 36.060 10.850 36.230 ;
        RECT 11.040 36.060 11.210 36.230 ;
        RECT 12.220 36.060 12.390 36.230 ;
        RECT 12.660 36.060 12.830 36.230 ;
        RECT 13.100 36.060 13.270 36.230 ;
        RECT 13.510 36.060 13.680 36.230 ;
        RECT 14.470 36.060 14.640 36.230 ;
        RECT 14.830 36.060 15.000 36.230 ;
        RECT 15.190 36.060 15.360 36.230 ;
        RECT 15.550 36.060 15.720 36.230 ;
        RECT 17.070 36.070 17.240 36.240 ;
        RECT 17.510 36.070 17.680 36.240 ;
        RECT 17.920 36.070 18.090 36.240 ;
        RECT 18.350 36.070 18.520 36.240 ;
        RECT 18.790 36.070 18.960 36.240 ;
        RECT 19.200 36.070 19.370 36.240 ;
        RECT 21.240 36.060 21.410 36.230 ;
        RECT 21.600 36.060 21.770 36.230 ;
        RECT 21.960 36.060 22.130 36.230 ;
        RECT 22.320 36.060 22.490 36.230 ;
        RECT 23.740 36.060 23.910 36.230 ;
        RECT 24.180 36.060 24.350 36.230 ;
        RECT 24.620 36.060 24.790 36.230 ;
        RECT 25.030 36.060 25.200 36.230 ;
        RECT 27.640 36.060 27.810 36.230 ;
        RECT 28.000 36.060 28.170 36.230 ;
        RECT 28.360 36.060 28.530 36.230 ;
        RECT 29.500 36.060 29.670 36.230 ;
        RECT 29.940 36.060 30.110 36.230 ;
        RECT 30.380 36.060 30.550 36.230 ;
        RECT 30.790 36.060 30.960 36.230 ;
        RECT 31.760 36.060 31.930 36.230 ;
        RECT 32.120 36.060 32.290 36.230 ;
        RECT 32.480 36.060 32.650 36.230 ;
        RECT 35.120 36.060 35.290 36.230 ;
        RECT 35.480 36.060 35.650 36.230 ;
        RECT 35.840 36.060 36.010 36.230 ;
        RECT 36.200 36.060 36.370 36.230 ;
        RECT 37.230 36.070 37.400 36.240 ;
        RECT 37.670 36.070 37.840 36.240 ;
        RECT 38.080 36.070 38.250 36.240 ;
        RECT 38.510 36.070 38.680 36.240 ;
        RECT 38.950 36.070 39.120 36.240 ;
        RECT 39.360 36.070 39.530 36.240 ;
        RECT 40.920 36.060 41.090 36.230 ;
        RECT 41.280 36.060 41.450 36.230 ;
        RECT 41.640 36.060 41.810 36.230 ;
        RECT 42.480 36.060 42.650 36.230 ;
        RECT 42.840 36.060 43.010 36.230 ;
        RECT 43.200 36.060 43.370 36.230 ;
        RECT 44.040 36.060 44.210 36.230 ;
        RECT 44.400 36.060 44.570 36.230 ;
        RECT 44.760 36.060 44.930 36.230 ;
        RECT 45.820 36.060 45.990 36.230 ;
        RECT 46.260 36.060 46.430 36.230 ;
        RECT 46.700 36.060 46.870 36.230 ;
        RECT 47.110 36.060 47.280 36.230 ;
        RECT 47.640 36.060 47.810 36.230 ;
        RECT 48.000 36.060 48.170 36.230 ;
        RECT 48.360 36.060 48.530 36.230 ;
        RECT 49.200 36.060 49.370 36.230 ;
        RECT 49.560 36.060 49.730 36.230 ;
        RECT 49.920 36.060 50.090 36.230 ;
        RECT 50.760 36.060 50.930 36.230 ;
        RECT 51.120 36.060 51.290 36.230 ;
        RECT 51.480 36.060 51.650 36.230 ;
        RECT 52.540 36.060 52.710 36.230 ;
        RECT 52.980 36.060 53.150 36.230 ;
        RECT 53.420 36.060 53.590 36.230 ;
        RECT 53.830 36.060 54.000 36.230 ;
        RECT 54.360 36.060 54.530 36.230 ;
        RECT 54.720 36.060 54.890 36.230 ;
        RECT 55.080 36.060 55.250 36.230 ;
        RECT 55.920 36.060 56.090 36.230 ;
        RECT 56.280 36.060 56.450 36.230 ;
        RECT 56.640 36.060 56.810 36.230 ;
        RECT 57.480 36.060 57.650 36.230 ;
        RECT 57.840 36.060 58.010 36.230 ;
        RECT 58.200 36.060 58.370 36.230 ;
        RECT 59.260 36.060 59.430 36.230 ;
        RECT 59.700 36.060 59.870 36.230 ;
        RECT 60.140 36.060 60.310 36.230 ;
        RECT 60.550 36.060 60.720 36.230 ;
        RECT 61.550 36.060 61.720 36.230 ;
        RECT 61.910 36.060 62.080 36.230 ;
        RECT 62.270 36.060 62.440 36.230 ;
        RECT 63.190 36.060 63.360 36.230 ;
        RECT 63.550 36.060 63.720 36.230 ;
        RECT 68.150 36.060 68.320 36.230 ;
        RECT 68.510 36.060 68.680 36.230 ;
        RECT 68.870 36.060 69.040 36.230 ;
        RECT 72.120 36.060 72.290 36.230 ;
        RECT 72.480 36.060 72.650 36.230 ;
        RECT 72.840 36.060 73.010 36.230 ;
        RECT 74.730 36.060 74.900 36.230 ;
        RECT 75.090 36.060 75.260 36.230 ;
        RECT 75.450 36.060 75.620 36.230 ;
        RECT 76.540 36.060 76.710 36.230 ;
        RECT 76.980 36.060 77.150 36.230 ;
        RECT 77.420 36.060 77.590 36.230 ;
        RECT 77.830 36.060 78.000 36.230 ;
        RECT 78.360 36.060 78.530 36.230 ;
        RECT 78.720 36.060 78.890 36.230 ;
        RECT 79.900 36.060 80.070 36.230 ;
        RECT 80.340 36.060 80.510 36.230 ;
        RECT 80.780 36.060 80.950 36.230 ;
        RECT 81.190 36.060 81.360 36.230 ;
        RECT 81.720 36.060 81.890 36.230 ;
        RECT 82.080 36.060 82.250 36.230 ;
        RECT 82.440 36.060 82.610 36.230 ;
        RECT 83.280 36.060 83.450 36.230 ;
        RECT 83.640 36.060 83.810 36.230 ;
        RECT 84.000 36.060 84.170 36.230 ;
        RECT 84.840 36.060 85.010 36.230 ;
        RECT 85.200 36.060 85.370 36.230 ;
        RECT 85.560 36.060 85.730 36.230 ;
        RECT 86.620 36.060 86.790 36.230 ;
        RECT 87.060 36.060 87.230 36.230 ;
        RECT 87.500 36.060 87.670 36.230 ;
        RECT 87.910 36.060 88.080 36.230 ;
        RECT 89.400 36.060 89.570 36.230 ;
        RECT 89.760 36.060 89.930 36.230 ;
        RECT 90.120 36.060 90.290 36.230 ;
        RECT 90.960 36.060 91.130 36.230 ;
        RECT 91.320 36.060 91.490 36.230 ;
        RECT 91.680 36.060 91.850 36.230 ;
        RECT 92.520 36.060 92.690 36.230 ;
        RECT 92.880 36.060 93.050 36.230 ;
        RECT 93.240 36.060 93.410 36.230 ;
        RECT 94.300 36.060 94.470 36.230 ;
        RECT 94.740 36.060 94.910 36.230 ;
        RECT 95.180 36.060 95.350 36.230 ;
        RECT 95.590 36.060 95.760 36.230 ;
        RECT 98.200 36.060 98.370 36.230 ;
        RECT 98.560 36.060 98.730 36.230 ;
        RECT 98.920 36.060 99.090 36.230 ;
        RECT 100.590 36.070 100.760 36.240 ;
        RECT 101.030 36.070 101.200 36.240 ;
        RECT 101.440 36.070 101.610 36.240 ;
        RECT 101.870 36.070 102.040 36.240 ;
        RECT 102.310 36.070 102.480 36.240 ;
        RECT 102.720 36.070 102.890 36.240 ;
        RECT 104.740 36.060 104.910 36.230 ;
        RECT 105.100 36.060 105.270 36.230 ;
        RECT 105.460 36.060 105.630 36.230 ;
        RECT 106.710 36.060 106.880 36.230 ;
        RECT 107.070 36.060 107.240 36.230 ;
        RECT 108.220 36.060 108.390 36.230 ;
        RECT 108.660 36.060 108.830 36.230 ;
        RECT 109.100 36.060 109.270 36.230 ;
        RECT 109.510 36.060 109.680 36.230 ;
        RECT 110.040 36.060 110.210 36.230 ;
        RECT 110.400 36.060 110.570 36.230 ;
        RECT 111.310 36.060 111.480 36.230 ;
        RECT 111.670 36.060 111.840 36.230 ;
        RECT 112.030 36.060 112.200 36.230 ;
        RECT 113.500 36.060 113.670 36.230 ;
        RECT 113.940 36.060 114.110 36.230 ;
        RECT 114.380 36.060 114.550 36.230 ;
        RECT 114.790 36.060 114.960 36.230 ;
        RECT 116.280 36.060 116.450 36.230 ;
        RECT 116.640 36.060 116.810 36.230 ;
        RECT 117.000 36.060 117.170 36.230 ;
        RECT 117.840 36.060 118.010 36.230 ;
        RECT 118.200 36.060 118.370 36.230 ;
        RECT 118.560 36.060 118.730 36.230 ;
        RECT 119.400 36.060 119.570 36.230 ;
        RECT 119.760 36.060 119.930 36.230 ;
        RECT 120.120 36.060 120.290 36.230 ;
        RECT 121.180 36.060 121.350 36.230 ;
        RECT 121.620 36.060 121.790 36.230 ;
        RECT 122.060 36.060 122.230 36.230 ;
        RECT 122.470 36.060 122.640 36.230 ;
        RECT 123.460 36.060 123.630 36.230 ;
        RECT 124.050 36.060 124.220 36.230 ;
        RECT 125.570 36.060 125.740 36.230 ;
        RECT 125.930 36.060 126.100 36.230 ;
        RECT 126.940 36.060 127.110 36.230 ;
        RECT 127.380 36.060 127.550 36.230 ;
        RECT 127.820 36.060 127.990 36.230 ;
        RECT 128.230 36.060 128.400 36.230 ;
        RECT 128.750 36.060 128.920 36.230 ;
        RECT 129.110 36.060 129.280 36.230 ;
        RECT 129.470 36.060 129.640 36.230 ;
        RECT 130.390 36.060 130.560 36.230 ;
        RECT 130.750 36.060 130.920 36.230 ;
        RECT 131.790 36.070 131.960 36.240 ;
        RECT 132.230 36.070 132.400 36.240 ;
        RECT 132.640 36.070 132.810 36.240 ;
        RECT 133.070 36.070 133.240 36.240 ;
        RECT 133.510 36.070 133.680 36.240 ;
        RECT 133.920 36.070 134.090 36.240 ;
        RECT 135.000 36.060 135.170 36.230 ;
        RECT 135.360 36.060 135.530 36.230 ;
        RECT 136.540 36.060 136.710 36.230 ;
        RECT 136.980 36.060 137.150 36.230 ;
        RECT 137.420 36.060 137.590 36.230 ;
        RECT 137.830 36.060 138.000 36.230 ;
        RECT 138.360 36.060 138.530 36.230 ;
        RECT 138.720 36.060 138.890 36.230 ;
        RECT 139.900 36.060 140.070 36.230 ;
        RECT 140.340 36.060 140.510 36.230 ;
        RECT 140.780 36.060 140.950 36.230 ;
        RECT 141.190 36.060 141.360 36.230 ;
        RECT 5.920 28.400 6.090 28.580 ;
        RECT 6.400 28.400 6.570 28.580 ;
        RECT 6.880 28.400 7.050 28.580 ;
        RECT 7.360 28.400 7.530 28.580 ;
        RECT 7.840 28.400 8.010 28.580 ;
        RECT 8.320 28.400 8.490 28.580 ;
        RECT 8.800 28.400 8.970 28.580 ;
        RECT 9.280 28.400 9.450 28.580 ;
        RECT 9.760 28.400 9.930 28.580 ;
        RECT 10.240 28.400 10.410 28.580 ;
        RECT 10.720 28.400 10.890 28.580 ;
        RECT 11.200 28.400 11.370 28.580 ;
        RECT 11.680 28.400 11.850 28.580 ;
        RECT 12.160 28.400 12.330 28.580 ;
        RECT 12.640 28.400 12.810 28.580 ;
        RECT 13.120 28.400 13.290 28.580 ;
        RECT 13.600 28.400 13.770 28.580 ;
        RECT 14.080 28.400 14.250 28.580 ;
        RECT 14.560 28.400 14.730 28.580 ;
        RECT 15.040 28.400 15.210 28.580 ;
        RECT 15.520 28.400 15.690 28.580 ;
        RECT 16.000 28.400 16.170 28.580 ;
        RECT 16.480 28.400 16.650 28.580 ;
        RECT 16.960 28.400 17.130 28.580 ;
        RECT 17.440 28.400 17.610 28.580 ;
        RECT 17.920 28.400 18.090 28.580 ;
        RECT 18.400 28.400 18.570 28.580 ;
        RECT 18.880 28.400 19.050 28.580 ;
        RECT 19.360 28.400 19.530 28.580 ;
        RECT 19.840 28.400 20.010 28.580 ;
        RECT 20.320 28.400 20.490 28.580 ;
        RECT 20.800 28.400 20.970 28.580 ;
        RECT 21.280 28.400 21.450 28.580 ;
        RECT 21.760 28.400 21.930 28.580 ;
        RECT 22.240 28.400 22.410 28.580 ;
        RECT 22.720 28.400 22.890 28.580 ;
        RECT 23.200 28.400 23.370 28.580 ;
        RECT 23.680 28.400 23.850 28.580 ;
        RECT 24.160 28.400 24.330 28.580 ;
        RECT 24.640 28.400 24.810 28.580 ;
        RECT 25.120 28.400 25.290 28.580 ;
        RECT 25.600 28.400 25.770 28.580 ;
        RECT 26.080 28.400 26.250 28.580 ;
        RECT 26.560 28.400 26.730 28.580 ;
        RECT 27.040 28.400 27.210 28.580 ;
        RECT 27.520 28.400 27.690 28.580 ;
        RECT 28.000 28.400 28.170 28.580 ;
        RECT 28.480 28.400 28.650 28.580 ;
        RECT 28.960 28.400 29.130 28.580 ;
        RECT 29.440 28.400 29.610 28.580 ;
        RECT 29.920 28.400 30.090 28.580 ;
        RECT 30.400 28.400 30.570 28.580 ;
        RECT 30.880 28.400 31.050 28.580 ;
        RECT 31.360 28.400 31.530 28.580 ;
        RECT 31.840 28.400 32.010 28.580 ;
        RECT 32.320 28.400 32.490 28.580 ;
        RECT 32.800 28.400 32.970 28.580 ;
        RECT 33.280 28.400 33.450 28.580 ;
        RECT 33.760 28.400 33.930 28.580 ;
        RECT 34.240 28.400 34.410 28.580 ;
        RECT 34.720 28.400 34.890 28.580 ;
        RECT 35.200 28.400 35.370 28.580 ;
        RECT 35.680 28.400 35.850 28.580 ;
        RECT 36.160 28.400 36.330 28.580 ;
        RECT 36.640 28.400 36.810 28.580 ;
        RECT 37.120 28.400 37.290 28.580 ;
        RECT 37.600 28.400 37.770 28.580 ;
        RECT 38.080 28.400 38.250 28.580 ;
        RECT 38.560 28.400 38.730 28.580 ;
        RECT 39.040 28.400 39.210 28.580 ;
        RECT 39.520 28.400 39.690 28.580 ;
        RECT 40.000 28.400 40.170 28.580 ;
        RECT 40.480 28.400 40.650 28.580 ;
        RECT 40.960 28.400 41.130 28.580 ;
        RECT 41.440 28.400 41.610 28.580 ;
        RECT 41.920 28.400 42.090 28.580 ;
        RECT 42.400 28.400 42.570 28.580 ;
        RECT 42.880 28.400 43.050 28.580 ;
        RECT 43.360 28.400 43.530 28.580 ;
        RECT 43.840 28.400 44.010 28.580 ;
        RECT 44.320 28.400 44.490 28.580 ;
        RECT 44.800 28.400 44.970 28.580 ;
        RECT 45.280 28.400 45.450 28.580 ;
        RECT 45.760 28.400 45.930 28.580 ;
        RECT 46.240 28.400 46.410 28.580 ;
        RECT 46.720 28.400 46.890 28.580 ;
        RECT 47.200 28.400 47.370 28.580 ;
        RECT 47.680 28.400 47.850 28.580 ;
        RECT 48.160 28.400 48.330 28.580 ;
        RECT 48.640 28.400 48.810 28.580 ;
        RECT 49.120 28.400 49.290 28.580 ;
        RECT 49.600 28.400 49.770 28.580 ;
        RECT 50.080 28.400 50.250 28.580 ;
        RECT 50.560 28.400 50.730 28.580 ;
        RECT 51.040 28.400 51.210 28.580 ;
        RECT 51.520 28.400 51.690 28.580 ;
        RECT 52.000 28.400 52.170 28.580 ;
        RECT 52.480 28.400 52.650 28.580 ;
        RECT 52.960 28.400 53.130 28.580 ;
        RECT 53.440 28.400 53.610 28.580 ;
        RECT 53.920 28.400 54.090 28.580 ;
        RECT 54.400 28.400 54.570 28.580 ;
        RECT 54.880 28.400 55.050 28.580 ;
        RECT 55.360 28.400 55.530 28.580 ;
        RECT 55.840 28.400 56.010 28.580 ;
        RECT 56.320 28.400 56.490 28.580 ;
        RECT 56.800 28.400 56.970 28.580 ;
        RECT 57.280 28.400 57.450 28.580 ;
        RECT 57.760 28.400 57.930 28.580 ;
        RECT 58.240 28.400 58.410 28.580 ;
        RECT 58.720 28.400 58.890 28.580 ;
        RECT 59.200 28.400 59.370 28.580 ;
        RECT 59.680 28.400 59.850 28.580 ;
        RECT 60.160 28.400 60.330 28.580 ;
        RECT 60.640 28.400 60.810 28.580 ;
        RECT 61.120 28.400 61.290 28.580 ;
        RECT 61.600 28.400 61.770 28.580 ;
        RECT 62.080 28.400 62.250 28.580 ;
        RECT 62.560 28.400 62.730 28.580 ;
        RECT 63.040 28.400 63.210 28.580 ;
        RECT 63.520 28.400 63.690 28.580 ;
        RECT 64.000 28.400 64.170 28.580 ;
        RECT 64.480 28.400 64.650 28.580 ;
        RECT 64.960 28.400 65.130 28.580 ;
        RECT 65.440 28.400 65.610 28.580 ;
        RECT 65.920 28.400 66.090 28.580 ;
        RECT 66.400 28.400 66.570 28.580 ;
        RECT 66.880 28.400 67.050 28.580 ;
        RECT 67.360 28.400 67.530 28.580 ;
        RECT 67.840 28.400 68.010 28.580 ;
        RECT 68.320 28.400 68.490 28.580 ;
        RECT 68.800 28.400 68.970 28.580 ;
        RECT 69.280 28.400 69.450 28.580 ;
        RECT 69.760 28.400 69.930 28.580 ;
        RECT 70.240 28.400 70.410 28.580 ;
        RECT 70.720 28.400 70.890 28.580 ;
        RECT 71.200 28.400 71.370 28.580 ;
        RECT 71.680 28.400 71.850 28.580 ;
        RECT 72.160 28.400 72.330 28.580 ;
        RECT 72.640 28.400 72.810 28.580 ;
        RECT 73.120 28.400 73.290 28.580 ;
        RECT 73.600 28.400 73.770 28.580 ;
        RECT 74.080 28.400 74.250 28.580 ;
        RECT 74.560 28.400 74.730 28.580 ;
        RECT 75.040 28.400 75.210 28.580 ;
        RECT 75.520 28.400 75.690 28.580 ;
        RECT 76.000 28.400 76.170 28.580 ;
        RECT 76.480 28.400 76.650 28.580 ;
        RECT 76.960 28.400 77.130 28.580 ;
        RECT 77.440 28.400 77.610 28.580 ;
        RECT 77.920 28.400 78.090 28.580 ;
        RECT 78.400 28.400 78.570 28.580 ;
        RECT 78.880 28.400 79.050 28.580 ;
        RECT 79.360 28.400 79.530 28.580 ;
        RECT 79.840 28.400 80.010 28.580 ;
        RECT 80.320 28.400 80.490 28.580 ;
        RECT 80.800 28.400 80.970 28.580 ;
        RECT 81.280 28.400 81.450 28.580 ;
        RECT 81.760 28.400 81.930 28.580 ;
        RECT 82.240 28.400 82.410 28.580 ;
        RECT 82.720 28.400 82.890 28.580 ;
        RECT 83.200 28.400 83.370 28.580 ;
        RECT 83.680 28.400 83.850 28.580 ;
        RECT 84.160 28.400 84.330 28.580 ;
        RECT 84.640 28.400 84.810 28.580 ;
        RECT 85.120 28.400 85.290 28.580 ;
        RECT 85.600 28.400 85.770 28.580 ;
        RECT 86.080 28.400 86.250 28.580 ;
        RECT 86.560 28.400 86.730 28.580 ;
        RECT 87.040 28.400 87.210 28.580 ;
        RECT 87.520 28.400 87.690 28.580 ;
        RECT 88.000 28.400 88.170 28.580 ;
        RECT 88.480 28.400 88.650 28.580 ;
        RECT 88.960 28.400 89.130 28.580 ;
        RECT 89.440 28.400 89.610 28.580 ;
        RECT 89.920 28.400 90.090 28.580 ;
        RECT 90.400 28.400 90.570 28.580 ;
        RECT 90.880 28.400 91.050 28.580 ;
        RECT 91.360 28.400 91.530 28.580 ;
        RECT 91.840 28.400 92.010 28.580 ;
        RECT 92.320 28.400 92.490 28.580 ;
        RECT 92.800 28.400 92.970 28.580 ;
        RECT 93.280 28.400 93.450 28.580 ;
        RECT 93.760 28.400 93.930 28.580 ;
        RECT 94.240 28.400 94.410 28.580 ;
        RECT 94.720 28.400 94.890 28.580 ;
        RECT 95.200 28.400 95.370 28.580 ;
        RECT 95.680 28.400 95.850 28.580 ;
        RECT 96.160 28.400 96.330 28.580 ;
        RECT 96.640 28.400 96.810 28.580 ;
        RECT 97.120 28.400 97.290 28.580 ;
        RECT 97.600 28.400 97.770 28.580 ;
        RECT 98.080 28.400 98.250 28.580 ;
        RECT 98.560 28.400 98.730 28.580 ;
        RECT 99.040 28.400 99.210 28.580 ;
        RECT 99.520 28.400 99.690 28.580 ;
        RECT 100.000 28.400 100.170 28.580 ;
        RECT 100.480 28.400 100.650 28.580 ;
        RECT 100.960 28.400 101.130 28.580 ;
        RECT 101.440 28.400 101.610 28.580 ;
        RECT 101.920 28.400 102.090 28.580 ;
        RECT 102.400 28.400 102.570 28.580 ;
        RECT 102.880 28.400 103.050 28.580 ;
        RECT 103.360 28.400 103.530 28.580 ;
        RECT 103.840 28.400 104.010 28.580 ;
      LAYER li1 ;
        RECT 104.160 28.400 104.640 28.580 ;
      LAYER li1 ;
        RECT 104.800 28.400 104.970 28.580 ;
        RECT 105.280 28.400 105.450 28.580 ;
        RECT 105.760 28.400 105.930 28.580 ;
        RECT 106.240 28.400 106.410 28.580 ;
        RECT 106.720 28.400 106.890 28.580 ;
        RECT 107.200 28.400 107.370 28.580 ;
        RECT 107.680 28.400 107.850 28.580 ;
        RECT 108.160 28.400 108.330 28.580 ;
        RECT 108.640 28.400 108.810 28.580 ;
        RECT 109.120 28.400 109.290 28.580 ;
        RECT 109.600 28.400 109.770 28.580 ;
        RECT 110.080 28.400 110.250 28.580 ;
        RECT 110.560 28.400 110.730 28.580 ;
        RECT 111.040 28.400 111.210 28.580 ;
        RECT 111.520 28.400 111.690 28.580 ;
        RECT 112.000 28.400 112.170 28.580 ;
        RECT 112.480 28.400 112.650 28.580 ;
        RECT 112.960 28.400 113.130 28.580 ;
        RECT 113.440 28.400 113.610 28.580 ;
        RECT 113.920 28.400 114.090 28.580 ;
        RECT 114.400 28.400 114.570 28.580 ;
        RECT 114.880 28.400 115.050 28.580 ;
        RECT 115.360 28.400 115.530 28.580 ;
        RECT 115.840 28.400 116.010 28.580 ;
        RECT 116.320 28.400 116.490 28.580 ;
        RECT 116.800 28.400 116.970 28.580 ;
        RECT 117.280 28.400 117.450 28.580 ;
        RECT 117.760 28.400 117.930 28.580 ;
        RECT 118.240 28.400 118.410 28.580 ;
        RECT 118.720 28.400 118.890 28.580 ;
        RECT 119.200 28.400 119.370 28.580 ;
      LAYER li1 ;
        RECT 119.520 28.400 120.000 28.580 ;
      LAYER li1 ;
        RECT 120.160 28.400 120.330 28.580 ;
        RECT 120.640 28.400 120.810 28.580 ;
        RECT 121.120 28.400 121.290 28.580 ;
        RECT 121.600 28.400 121.770 28.580 ;
        RECT 122.080 28.400 122.250 28.580 ;
        RECT 122.560 28.400 122.730 28.580 ;
        RECT 123.040 28.400 123.210 28.580 ;
        RECT 123.520 28.400 123.690 28.580 ;
        RECT 124.000 28.400 124.170 28.580 ;
        RECT 124.480 28.400 124.650 28.580 ;
        RECT 124.960 28.400 125.130 28.580 ;
        RECT 125.440 28.400 125.610 28.580 ;
        RECT 125.920 28.400 126.090 28.580 ;
        RECT 126.400 28.400 126.570 28.580 ;
        RECT 126.880 28.400 127.050 28.580 ;
        RECT 127.360 28.400 127.530 28.580 ;
        RECT 127.840 28.400 128.010 28.580 ;
        RECT 128.320 28.400 128.490 28.580 ;
        RECT 128.800 28.400 128.970 28.580 ;
        RECT 129.280 28.400 129.450 28.580 ;
        RECT 129.760 28.400 129.930 28.580 ;
        RECT 130.240 28.400 130.410 28.580 ;
        RECT 130.720 28.400 130.890 28.580 ;
        RECT 131.200 28.400 131.370 28.580 ;
        RECT 131.680 28.400 131.850 28.580 ;
      LAYER li1 ;
        RECT 132.000 28.400 132.480 28.580 ;
      LAYER li1 ;
        RECT 132.640 28.400 132.810 28.580 ;
        RECT 133.120 28.400 133.290 28.580 ;
        RECT 133.600 28.400 133.770 28.580 ;
        RECT 134.080 28.400 134.250 28.580 ;
        RECT 134.560 28.400 134.730 28.580 ;
        RECT 135.040 28.400 135.210 28.580 ;
        RECT 135.520 28.400 135.690 28.580 ;
        RECT 136.000 28.400 136.170 28.580 ;
        RECT 136.480 28.400 136.650 28.580 ;
        RECT 136.960 28.400 137.130 28.580 ;
        RECT 137.440 28.400 137.610 28.580 ;
        RECT 137.920 28.400 138.090 28.580 ;
        RECT 138.400 28.400 138.570 28.580 ;
        RECT 138.880 28.400 139.050 28.580 ;
        RECT 139.360 28.400 139.530 28.580 ;
        RECT 139.840 28.400 140.010 28.580 ;
        RECT 140.320 28.400 140.490 28.580 ;
        RECT 140.800 28.400 140.970 28.580 ;
        RECT 141.280 28.400 141.450 28.580 ;
      LAYER li1 ;
        RECT 141.600 28.400 142.080 28.580 ;
      LAYER li1 ;
        RECT 6.510 27.930 6.680 28.100 ;
        RECT 6.950 27.930 7.120 28.100 ;
        RECT 7.360 27.930 7.530 28.100 ;
        RECT 7.790 27.930 7.960 28.100 ;
        RECT 8.230 27.930 8.400 28.100 ;
        RECT 8.640 27.930 8.810 28.100 ;
        RECT 10.350 27.930 10.520 28.100 ;
        RECT 10.790 27.930 10.960 28.100 ;
        RECT 11.200 27.930 11.370 28.100 ;
        RECT 11.630 27.930 11.800 28.100 ;
        RECT 12.070 27.930 12.240 28.100 ;
        RECT 12.480 27.930 12.650 28.100 ;
        RECT 15.000 27.920 15.170 28.090 ;
        RECT 15.360 27.920 15.530 28.090 ;
        RECT 16.540 27.920 16.710 28.090 ;
        RECT 16.980 27.920 17.150 28.090 ;
        RECT 17.420 27.920 17.590 28.090 ;
        RECT 17.830 27.920 18.000 28.090 ;
        RECT 18.350 27.920 18.520 28.090 ;
        RECT 18.710 27.920 18.880 28.090 ;
        RECT 19.070 27.920 19.240 28.090 ;
        RECT 19.990 27.920 20.160 28.090 ;
        RECT 20.350 27.920 20.520 28.090 ;
        RECT 20.860 27.920 21.030 28.090 ;
        RECT 21.300 27.920 21.470 28.090 ;
        RECT 21.740 27.920 21.910 28.090 ;
        RECT 22.150 27.920 22.320 28.090 ;
        RECT 23.110 27.920 23.280 28.090 ;
        RECT 23.470 27.920 23.640 28.090 ;
        RECT 23.830 27.920 24.000 28.090 ;
        RECT 24.190 27.920 24.360 28.090 ;
        RECT 25.180 27.920 25.350 28.090 ;
        RECT 25.620 27.920 25.790 28.090 ;
        RECT 26.060 27.920 26.230 28.090 ;
        RECT 26.470 27.920 26.640 28.090 ;
        RECT 26.990 27.920 27.160 28.090 ;
        RECT 27.350 27.920 27.520 28.090 ;
        RECT 27.710 27.920 27.880 28.090 ;
        RECT 28.630 27.920 28.800 28.090 ;
        RECT 28.990 27.920 29.160 28.090 ;
        RECT 29.500 27.920 29.670 28.090 ;
        RECT 29.940 27.920 30.110 28.090 ;
        RECT 30.380 27.920 30.550 28.090 ;
        RECT 30.790 27.920 30.960 28.090 ;
        RECT 31.300 27.920 31.470 28.090 ;
        RECT 31.660 27.920 31.830 28.090 ;
        RECT 32.020 27.920 32.190 28.090 ;
        RECT 32.380 27.920 32.550 28.090 ;
        RECT 32.740 27.920 32.910 28.090 ;
        RECT 35.310 27.930 35.480 28.100 ;
        RECT 35.750 27.930 35.920 28.100 ;
        RECT 36.160 27.930 36.330 28.100 ;
        RECT 36.590 27.930 36.760 28.100 ;
        RECT 37.030 27.930 37.200 28.100 ;
        RECT 37.440 27.930 37.610 28.100 ;
        RECT 39.480 27.920 39.650 28.090 ;
        RECT 39.840 27.920 40.010 28.090 ;
        RECT 40.750 27.920 40.920 28.090 ;
        RECT 41.110 27.920 41.280 28.090 ;
        RECT 41.470 27.920 41.640 28.090 ;
        RECT 42.940 27.920 43.110 28.090 ;
        RECT 43.380 27.920 43.550 28.090 ;
        RECT 43.820 27.920 43.990 28.090 ;
        RECT 44.230 27.920 44.400 28.090 ;
        RECT 45.220 27.920 45.390 28.090 ;
        RECT 45.810 27.920 45.980 28.090 ;
        RECT 47.330 27.920 47.500 28.090 ;
        RECT 47.690 27.920 47.860 28.090 ;
        RECT 49.230 27.930 49.400 28.100 ;
        RECT 49.670 27.930 49.840 28.100 ;
        RECT 50.080 27.930 50.250 28.100 ;
        RECT 50.510 27.930 50.680 28.100 ;
        RECT 50.950 27.930 51.120 28.100 ;
        RECT 51.360 27.930 51.530 28.100 ;
        RECT 52.920 27.920 53.090 28.090 ;
        RECT 53.280 27.920 53.450 28.090 ;
        RECT 53.640 27.920 53.810 28.090 ;
        RECT 54.480 27.920 54.650 28.090 ;
        RECT 54.840 27.920 55.010 28.090 ;
        RECT 55.200 27.920 55.370 28.090 ;
        RECT 56.040 27.920 56.210 28.090 ;
        RECT 56.400 27.920 56.570 28.090 ;
        RECT 56.760 27.920 56.930 28.090 ;
        RECT 57.820 27.920 57.990 28.090 ;
        RECT 58.260 27.920 58.430 28.090 ;
        RECT 58.700 27.920 58.870 28.090 ;
        RECT 59.110 27.920 59.280 28.090 ;
        RECT 59.640 27.920 59.810 28.090 ;
        RECT 60.000 27.920 60.170 28.090 ;
        RECT 60.360 27.920 60.530 28.090 ;
        RECT 61.200 27.920 61.370 28.090 ;
        RECT 61.560 27.920 61.730 28.090 ;
        RECT 61.920 27.920 62.090 28.090 ;
        RECT 62.760 27.920 62.930 28.090 ;
        RECT 63.120 27.920 63.290 28.090 ;
        RECT 63.480 27.920 63.650 28.090 ;
        RECT 64.540 27.920 64.710 28.090 ;
        RECT 64.980 27.920 65.150 28.090 ;
        RECT 65.420 27.920 65.590 28.090 ;
        RECT 65.830 27.920 66.000 28.090 ;
        RECT 66.360 27.920 66.530 28.090 ;
        RECT 66.720 27.920 66.890 28.090 ;
        RECT 67.080 27.920 67.250 28.090 ;
        RECT 67.920 27.920 68.090 28.090 ;
        RECT 68.280 27.920 68.450 28.090 ;
        RECT 68.640 27.920 68.810 28.090 ;
        RECT 69.480 27.920 69.650 28.090 ;
        RECT 69.840 27.920 70.010 28.090 ;
        RECT 70.200 27.920 70.370 28.090 ;
        RECT 71.260 27.920 71.430 28.090 ;
        RECT 71.700 27.920 71.870 28.090 ;
        RECT 72.140 27.920 72.310 28.090 ;
        RECT 72.550 27.920 72.720 28.090 ;
        RECT 73.080 27.920 73.250 28.090 ;
        RECT 73.440 27.920 73.610 28.090 ;
        RECT 73.800 27.920 73.970 28.090 ;
        RECT 74.640 27.920 74.810 28.090 ;
        RECT 75.000 27.920 75.170 28.090 ;
        RECT 75.360 27.920 75.530 28.090 ;
        RECT 76.200 27.920 76.370 28.090 ;
        RECT 76.560 27.920 76.730 28.090 ;
        RECT 76.920 27.920 77.090 28.090 ;
        RECT 78.510 27.930 78.680 28.100 ;
        RECT 78.950 27.930 79.120 28.100 ;
        RECT 79.360 27.930 79.530 28.100 ;
        RECT 79.790 27.930 79.960 28.100 ;
        RECT 80.230 27.930 80.400 28.100 ;
        RECT 80.640 27.930 80.810 28.100 ;
        RECT 82.630 27.920 82.800 28.090 ;
        RECT 82.990 27.920 83.160 28.090 ;
        RECT 83.350 27.920 83.520 28.090 ;
        RECT 83.710 27.920 83.880 28.090 ;
        RECT 85.230 27.930 85.400 28.100 ;
        RECT 85.670 27.930 85.840 28.100 ;
        RECT 86.080 27.930 86.250 28.100 ;
        RECT 86.510 27.930 86.680 28.100 ;
        RECT 86.950 27.930 87.120 28.100 ;
        RECT 87.360 27.930 87.530 28.100 ;
        RECT 88.910 27.920 89.080 28.090 ;
        RECT 89.270 27.920 89.440 28.090 ;
        RECT 89.630 27.920 89.800 28.090 ;
        RECT 90.550 27.920 90.720 28.090 ;
        RECT 90.910 27.920 91.080 28.090 ;
        RECT 91.420 27.920 91.590 28.090 ;
        RECT 91.860 27.920 92.030 28.090 ;
        RECT 92.300 27.920 92.470 28.090 ;
        RECT 92.710 27.920 92.880 28.090 ;
        RECT 94.680 27.920 94.850 28.090 ;
        RECT 95.040 27.920 95.210 28.090 ;
        RECT 95.400 27.920 95.570 28.090 ;
        RECT 95.760 27.920 95.930 28.090 ;
        RECT 97.180 27.920 97.350 28.090 ;
        RECT 97.620 27.920 97.790 28.090 ;
        RECT 98.060 27.920 98.230 28.090 ;
        RECT 98.470 27.920 98.640 28.090 ;
        RECT 99.000 27.920 99.170 28.090 ;
        RECT 99.360 27.920 99.530 28.090 ;
        RECT 100.540 27.920 100.710 28.090 ;
        RECT 100.980 27.920 101.150 28.090 ;
        RECT 101.420 27.920 101.590 28.090 ;
        RECT 101.830 27.920 102.000 28.090 ;
        RECT 102.790 27.920 102.960 28.090 ;
        RECT 103.150 27.920 103.320 28.090 ;
        RECT 103.510 27.920 103.680 28.090 ;
        RECT 103.870 27.920 104.040 28.090 ;
        RECT 104.860 27.920 105.030 28.090 ;
        RECT 105.300 27.920 105.470 28.090 ;
        RECT 105.740 27.920 105.910 28.090 ;
        RECT 106.150 27.920 106.320 28.090 ;
        RECT 107.110 27.920 107.280 28.090 ;
        RECT 107.470 27.920 107.640 28.090 ;
        RECT 107.830 27.920 108.000 28.090 ;
        RECT 108.190 27.920 108.360 28.090 ;
        RECT 109.180 27.920 109.350 28.090 ;
        RECT 109.620 27.920 109.790 28.090 ;
        RECT 110.060 27.920 110.230 28.090 ;
        RECT 110.470 27.920 110.640 28.090 ;
        RECT 111.000 27.920 111.170 28.090 ;
        RECT 111.360 27.920 111.530 28.090 ;
        RECT 111.720 27.920 111.890 28.090 ;
        RECT 112.080 27.920 112.250 28.090 ;
        RECT 113.500 27.920 113.670 28.090 ;
        RECT 113.940 27.920 114.110 28.090 ;
        RECT 114.380 27.920 114.550 28.090 ;
        RECT 114.790 27.920 114.960 28.090 ;
        RECT 115.320 27.920 115.490 28.090 ;
        RECT 115.680 27.920 115.850 28.090 ;
        RECT 116.590 27.920 116.760 28.090 ;
        RECT 116.950 27.920 117.120 28.090 ;
        RECT 117.310 27.920 117.480 28.090 ;
        RECT 118.780 27.920 118.950 28.090 ;
        RECT 119.220 27.920 119.390 28.090 ;
        RECT 119.660 27.920 119.830 28.090 ;
        RECT 120.070 27.920 120.240 28.090 ;
        RECT 120.860 27.920 121.030 28.090 ;
        RECT 121.220 27.920 121.390 28.090 ;
        RECT 121.580 27.920 121.750 28.090 ;
        RECT 121.940 27.920 122.110 28.090 ;
        RECT 122.300 27.920 122.470 28.090 ;
        RECT 123.190 27.920 123.360 28.090 ;
        RECT 123.550 27.920 123.720 28.090 ;
        RECT 124.060 27.920 124.230 28.090 ;
        RECT 124.500 27.920 124.670 28.090 ;
        RECT 124.940 27.920 125.110 28.090 ;
        RECT 125.350 27.920 125.520 28.090 ;
        RECT 125.880 27.920 126.050 28.090 ;
        RECT 126.240 27.920 126.410 28.090 ;
        RECT 127.420 27.920 127.590 28.090 ;
        RECT 127.860 27.920 128.030 28.090 ;
        RECT 128.300 27.920 128.470 28.090 ;
        RECT 128.710 27.920 128.880 28.090 ;
        RECT 129.670 27.920 129.840 28.090 ;
        RECT 130.030 27.920 130.200 28.090 ;
        RECT 130.390 27.920 130.560 28.090 ;
        RECT 130.750 27.920 130.920 28.090 ;
        RECT 131.740 27.920 131.910 28.090 ;
        RECT 132.180 27.920 132.350 28.090 ;
        RECT 132.620 27.920 132.790 28.090 ;
        RECT 133.030 27.920 133.200 28.090 ;
        RECT 136.000 27.920 136.170 28.090 ;
        RECT 136.360 27.920 136.530 28.090 ;
        RECT 137.550 27.930 137.720 28.100 ;
        RECT 137.990 27.930 138.160 28.100 ;
        RECT 138.400 27.930 138.570 28.100 ;
        RECT 138.830 27.930 139.000 28.100 ;
        RECT 139.270 27.930 139.440 28.100 ;
        RECT 139.680 27.930 139.850 28.100 ;
        RECT 5.920 20.260 6.090 20.440 ;
        RECT 6.400 20.260 6.570 20.440 ;
        RECT 6.880 20.260 7.050 20.440 ;
        RECT 7.360 20.260 7.530 20.440 ;
        RECT 7.840 20.260 8.010 20.440 ;
        RECT 8.320 20.260 8.490 20.440 ;
        RECT 8.800 20.260 8.970 20.440 ;
        RECT 9.280 20.260 9.450 20.440 ;
        RECT 9.760 20.260 9.930 20.440 ;
        RECT 10.240 20.260 10.410 20.440 ;
        RECT 10.720 20.260 10.890 20.440 ;
        RECT 11.200 20.260 11.370 20.440 ;
        RECT 11.680 20.260 11.850 20.440 ;
        RECT 12.160 20.260 12.330 20.440 ;
        RECT 12.640 20.260 12.810 20.440 ;
        RECT 13.120 20.260 13.290 20.440 ;
        RECT 13.600 20.260 13.770 20.440 ;
        RECT 14.080 20.260 14.250 20.440 ;
        RECT 14.560 20.260 14.730 20.440 ;
        RECT 15.040 20.260 15.210 20.440 ;
        RECT 15.520 20.260 15.690 20.440 ;
        RECT 16.000 20.260 16.170 20.440 ;
        RECT 16.480 20.260 16.650 20.440 ;
        RECT 16.960 20.260 17.130 20.440 ;
        RECT 17.440 20.260 17.610 20.440 ;
        RECT 17.920 20.260 18.090 20.440 ;
        RECT 18.400 20.260 18.570 20.440 ;
        RECT 18.880 20.260 19.050 20.440 ;
        RECT 19.360 20.260 19.530 20.440 ;
        RECT 19.840 20.260 20.010 20.440 ;
        RECT 20.320 20.260 20.490 20.440 ;
        RECT 20.800 20.260 20.970 20.440 ;
        RECT 21.280 20.260 21.450 20.440 ;
        RECT 21.760 20.260 21.930 20.440 ;
        RECT 22.240 20.260 22.410 20.440 ;
        RECT 22.720 20.260 22.890 20.440 ;
        RECT 23.200 20.260 23.370 20.440 ;
        RECT 23.680 20.260 23.850 20.440 ;
        RECT 24.160 20.260 24.330 20.440 ;
        RECT 24.640 20.260 24.810 20.440 ;
        RECT 25.120 20.260 25.290 20.440 ;
        RECT 25.600 20.260 25.770 20.440 ;
        RECT 26.080 20.260 26.250 20.440 ;
        RECT 26.560 20.260 26.730 20.440 ;
        RECT 27.040 20.260 27.210 20.440 ;
        RECT 27.520 20.260 27.690 20.440 ;
        RECT 28.000 20.260 28.170 20.440 ;
        RECT 28.480 20.260 28.650 20.440 ;
        RECT 28.960 20.260 29.130 20.440 ;
        RECT 29.440 20.260 29.610 20.440 ;
        RECT 29.920 20.260 30.090 20.440 ;
        RECT 30.400 20.260 30.570 20.440 ;
        RECT 30.880 20.260 31.050 20.440 ;
        RECT 31.360 20.260 31.530 20.440 ;
        RECT 31.840 20.260 32.010 20.440 ;
        RECT 32.320 20.260 32.490 20.440 ;
        RECT 32.800 20.260 32.970 20.440 ;
        RECT 33.280 20.260 33.450 20.440 ;
        RECT 33.760 20.260 33.930 20.440 ;
        RECT 34.240 20.260 34.410 20.440 ;
        RECT 34.720 20.260 34.890 20.440 ;
        RECT 35.200 20.260 35.370 20.440 ;
        RECT 35.680 20.260 35.850 20.440 ;
        RECT 36.160 20.260 36.330 20.440 ;
        RECT 36.640 20.260 36.810 20.440 ;
        RECT 37.120 20.260 37.290 20.440 ;
        RECT 37.600 20.260 37.770 20.440 ;
        RECT 38.080 20.260 38.250 20.440 ;
        RECT 38.560 20.260 38.730 20.440 ;
        RECT 39.040 20.260 39.210 20.440 ;
        RECT 39.520 20.260 39.690 20.440 ;
        RECT 40.000 20.260 40.170 20.440 ;
        RECT 40.480 20.260 40.650 20.440 ;
        RECT 40.960 20.260 41.130 20.440 ;
        RECT 41.440 20.260 41.610 20.440 ;
        RECT 41.920 20.260 42.090 20.440 ;
        RECT 42.400 20.260 42.570 20.440 ;
        RECT 42.880 20.260 43.050 20.440 ;
        RECT 43.360 20.260 43.530 20.440 ;
        RECT 43.840 20.260 44.010 20.440 ;
        RECT 44.320 20.260 44.490 20.440 ;
        RECT 44.800 20.260 44.970 20.440 ;
        RECT 45.280 20.260 45.450 20.440 ;
        RECT 45.760 20.260 45.930 20.440 ;
        RECT 46.240 20.260 46.410 20.440 ;
        RECT 46.720 20.260 46.890 20.440 ;
        RECT 47.200 20.260 47.370 20.440 ;
        RECT 47.680 20.260 47.850 20.440 ;
        RECT 48.160 20.260 48.330 20.440 ;
        RECT 48.640 20.260 48.810 20.440 ;
        RECT 49.120 20.260 49.290 20.440 ;
        RECT 49.600 20.260 49.770 20.440 ;
        RECT 50.080 20.260 50.250 20.440 ;
        RECT 50.560 20.260 50.730 20.440 ;
        RECT 51.040 20.260 51.210 20.440 ;
        RECT 51.520 20.260 51.690 20.440 ;
        RECT 52.000 20.260 52.170 20.440 ;
        RECT 52.480 20.260 52.650 20.440 ;
        RECT 52.960 20.260 53.130 20.440 ;
        RECT 53.440 20.260 53.610 20.440 ;
        RECT 53.920 20.260 54.090 20.440 ;
        RECT 54.400 20.260 54.570 20.440 ;
        RECT 54.880 20.260 55.050 20.440 ;
        RECT 55.360 20.260 55.530 20.440 ;
        RECT 55.840 20.260 56.010 20.440 ;
        RECT 56.320 20.260 56.490 20.440 ;
        RECT 56.800 20.260 56.970 20.440 ;
        RECT 57.280 20.260 57.450 20.440 ;
        RECT 57.760 20.260 57.930 20.440 ;
        RECT 58.240 20.260 58.410 20.440 ;
        RECT 58.720 20.260 58.890 20.440 ;
        RECT 59.200 20.260 59.370 20.440 ;
        RECT 59.680 20.260 59.850 20.440 ;
        RECT 60.160 20.260 60.330 20.440 ;
        RECT 60.640 20.260 60.810 20.440 ;
        RECT 61.120 20.260 61.290 20.440 ;
        RECT 61.600 20.260 61.770 20.440 ;
        RECT 62.080 20.260 62.250 20.440 ;
        RECT 62.560 20.260 62.730 20.440 ;
        RECT 63.040 20.260 63.210 20.440 ;
        RECT 63.520 20.260 63.690 20.440 ;
        RECT 64.000 20.260 64.170 20.440 ;
        RECT 64.480 20.260 64.650 20.440 ;
        RECT 64.960 20.260 65.130 20.440 ;
        RECT 65.440 20.260 65.610 20.440 ;
        RECT 65.920 20.260 66.090 20.440 ;
        RECT 66.400 20.260 66.570 20.440 ;
        RECT 66.880 20.260 67.050 20.440 ;
        RECT 67.360 20.260 67.530 20.440 ;
        RECT 67.840 20.260 68.010 20.440 ;
        RECT 68.320 20.260 68.490 20.440 ;
        RECT 68.800 20.260 68.970 20.440 ;
        RECT 69.280 20.260 69.450 20.440 ;
        RECT 69.760 20.260 69.930 20.440 ;
        RECT 70.240 20.260 70.410 20.440 ;
        RECT 70.720 20.260 70.890 20.440 ;
        RECT 71.200 20.260 71.370 20.440 ;
        RECT 71.680 20.260 71.850 20.440 ;
        RECT 72.160 20.260 72.330 20.440 ;
        RECT 72.640 20.260 72.810 20.440 ;
        RECT 73.120 20.260 73.290 20.440 ;
        RECT 73.600 20.260 73.770 20.440 ;
        RECT 74.080 20.260 74.250 20.440 ;
        RECT 74.560 20.260 74.730 20.440 ;
        RECT 75.040 20.260 75.210 20.440 ;
        RECT 75.520 20.260 75.690 20.440 ;
        RECT 76.000 20.260 76.170 20.440 ;
        RECT 76.480 20.260 76.650 20.440 ;
        RECT 76.960 20.260 77.130 20.440 ;
        RECT 77.440 20.260 77.610 20.440 ;
        RECT 77.920 20.260 78.090 20.440 ;
        RECT 78.400 20.260 78.570 20.440 ;
        RECT 78.880 20.260 79.050 20.440 ;
        RECT 79.360 20.260 79.530 20.440 ;
        RECT 79.840 20.260 80.010 20.440 ;
        RECT 80.320 20.260 80.490 20.440 ;
        RECT 80.800 20.260 80.970 20.440 ;
        RECT 81.280 20.260 81.450 20.440 ;
        RECT 81.760 20.260 81.930 20.440 ;
        RECT 82.240 20.260 82.410 20.440 ;
        RECT 82.720 20.260 82.890 20.440 ;
        RECT 83.200 20.260 83.370 20.440 ;
        RECT 83.680 20.260 83.850 20.440 ;
        RECT 84.160 20.260 84.330 20.440 ;
        RECT 84.640 20.260 84.810 20.440 ;
        RECT 85.120 20.260 85.290 20.440 ;
        RECT 85.600 20.260 85.770 20.440 ;
        RECT 86.080 20.260 86.250 20.440 ;
        RECT 86.560 20.260 86.730 20.440 ;
        RECT 87.040 20.260 87.210 20.440 ;
        RECT 87.520 20.260 87.690 20.440 ;
        RECT 88.000 20.260 88.170 20.440 ;
        RECT 88.480 20.260 88.650 20.440 ;
        RECT 88.960 20.260 89.130 20.440 ;
        RECT 89.440 20.260 89.610 20.440 ;
        RECT 89.920 20.260 90.090 20.440 ;
        RECT 90.400 20.260 90.570 20.440 ;
        RECT 90.880 20.260 91.050 20.440 ;
        RECT 91.360 20.260 91.530 20.440 ;
        RECT 91.840 20.260 92.010 20.440 ;
        RECT 92.320 20.260 92.490 20.440 ;
        RECT 92.800 20.260 92.970 20.440 ;
        RECT 93.280 20.260 93.450 20.440 ;
        RECT 93.760 20.260 93.930 20.440 ;
        RECT 94.240 20.260 94.410 20.440 ;
        RECT 94.720 20.260 94.890 20.440 ;
        RECT 95.200 20.260 95.370 20.440 ;
        RECT 95.680 20.260 95.850 20.440 ;
        RECT 96.160 20.260 96.330 20.440 ;
        RECT 96.640 20.260 96.810 20.440 ;
        RECT 97.120 20.260 97.290 20.440 ;
        RECT 97.600 20.260 97.770 20.440 ;
        RECT 98.080 20.260 98.250 20.440 ;
        RECT 98.560 20.260 98.730 20.440 ;
        RECT 99.040 20.260 99.210 20.440 ;
        RECT 99.520 20.260 99.690 20.440 ;
        RECT 100.000 20.260 100.170 20.440 ;
        RECT 100.480 20.260 100.650 20.440 ;
        RECT 100.960 20.260 101.130 20.440 ;
        RECT 101.440 20.260 101.610 20.440 ;
        RECT 101.920 20.260 102.090 20.440 ;
        RECT 102.400 20.260 102.570 20.440 ;
        RECT 102.880 20.260 103.050 20.440 ;
        RECT 103.360 20.260 103.530 20.440 ;
        RECT 103.840 20.260 104.010 20.440 ;
        RECT 104.320 20.260 104.490 20.440 ;
        RECT 104.800 20.260 104.970 20.440 ;
        RECT 105.280 20.260 105.450 20.440 ;
        RECT 105.760 20.260 105.930 20.440 ;
        RECT 106.240 20.260 106.410 20.440 ;
        RECT 106.720 20.260 106.890 20.440 ;
        RECT 107.200 20.260 107.370 20.440 ;
        RECT 107.680 20.260 107.850 20.440 ;
        RECT 108.160 20.260 108.330 20.440 ;
        RECT 108.640 20.260 108.810 20.440 ;
        RECT 109.120 20.260 109.290 20.440 ;
        RECT 109.600 20.260 109.770 20.440 ;
        RECT 110.080 20.260 110.250 20.440 ;
        RECT 110.560 20.260 110.730 20.440 ;
        RECT 111.040 20.260 111.210 20.440 ;
        RECT 111.520 20.260 111.690 20.440 ;
        RECT 112.000 20.260 112.170 20.440 ;
        RECT 112.480 20.260 112.650 20.440 ;
        RECT 112.960 20.260 113.130 20.440 ;
        RECT 113.440 20.260 113.610 20.440 ;
        RECT 113.920 20.260 114.090 20.440 ;
        RECT 114.400 20.260 114.570 20.440 ;
        RECT 114.880 20.260 115.050 20.440 ;
        RECT 115.360 20.260 115.530 20.440 ;
        RECT 115.840 20.260 116.010 20.440 ;
        RECT 116.320 20.260 116.490 20.440 ;
        RECT 116.800 20.260 116.970 20.440 ;
        RECT 117.280 20.260 117.450 20.440 ;
        RECT 117.760 20.260 117.930 20.440 ;
        RECT 118.240 20.260 118.410 20.440 ;
        RECT 118.720 20.260 118.890 20.440 ;
        RECT 119.200 20.260 119.370 20.440 ;
        RECT 119.680 20.260 119.850 20.440 ;
        RECT 120.160 20.260 120.330 20.440 ;
        RECT 120.640 20.260 120.810 20.440 ;
        RECT 121.120 20.260 121.290 20.440 ;
        RECT 121.600 20.260 121.770 20.440 ;
        RECT 122.080 20.260 122.250 20.440 ;
        RECT 122.560 20.260 122.730 20.440 ;
        RECT 123.040 20.260 123.210 20.440 ;
        RECT 123.520 20.260 123.690 20.440 ;
        RECT 124.000 20.260 124.170 20.440 ;
        RECT 124.480 20.260 124.650 20.440 ;
        RECT 124.960 20.260 125.130 20.440 ;
        RECT 125.440 20.260 125.610 20.440 ;
        RECT 125.920 20.260 126.090 20.440 ;
        RECT 126.400 20.260 126.570 20.440 ;
        RECT 126.880 20.260 127.050 20.440 ;
        RECT 127.360 20.260 127.530 20.440 ;
        RECT 127.840 20.260 128.010 20.440 ;
        RECT 128.320 20.260 128.490 20.440 ;
        RECT 128.800 20.260 128.970 20.440 ;
        RECT 129.280 20.260 129.450 20.440 ;
        RECT 129.760 20.260 129.930 20.440 ;
        RECT 130.240 20.260 130.410 20.440 ;
        RECT 130.720 20.260 130.890 20.440 ;
        RECT 131.200 20.260 131.370 20.440 ;
        RECT 131.680 20.260 131.850 20.440 ;
        RECT 132.160 20.260 132.330 20.440 ;
        RECT 132.640 20.260 132.810 20.440 ;
        RECT 133.120 20.260 133.290 20.440 ;
        RECT 133.600 20.260 133.770 20.440 ;
        RECT 134.080 20.260 134.250 20.440 ;
        RECT 134.560 20.260 134.730 20.440 ;
        RECT 135.040 20.260 135.210 20.440 ;
        RECT 135.520 20.260 135.690 20.440 ;
        RECT 136.000 20.260 136.170 20.440 ;
        RECT 136.480 20.260 136.650 20.440 ;
        RECT 136.960 20.260 137.130 20.440 ;
        RECT 137.440 20.260 137.610 20.440 ;
        RECT 137.920 20.260 138.090 20.440 ;
        RECT 138.400 20.260 138.570 20.440 ;
        RECT 138.880 20.260 139.050 20.440 ;
        RECT 139.360 20.260 139.530 20.440 ;
        RECT 139.840 20.260 140.010 20.440 ;
        RECT 140.320 20.260 140.490 20.440 ;
        RECT 140.800 20.260 140.970 20.440 ;
        RECT 141.280 20.260 141.450 20.440 ;
        RECT 141.760 20.260 141.930 20.440 ;
        RECT 6.510 19.790 6.680 19.960 ;
        RECT 6.950 19.790 7.120 19.960 ;
        RECT 7.360 19.790 7.530 19.960 ;
        RECT 7.790 19.790 7.960 19.960 ;
        RECT 8.230 19.790 8.400 19.960 ;
        RECT 8.640 19.790 8.810 19.960 ;
        RECT 9.820 19.780 9.990 19.950 ;
        RECT 10.260 19.780 10.430 19.950 ;
        RECT 10.700 19.780 10.870 19.950 ;
        RECT 11.110 19.780 11.280 19.950 ;
        RECT 13.120 19.780 13.290 19.950 ;
        RECT 13.480 19.780 13.650 19.950 ;
        RECT 14.140 19.780 14.310 19.950 ;
        RECT 14.580 19.780 14.750 19.950 ;
        RECT 15.020 19.780 15.190 19.950 ;
        RECT 15.430 19.780 15.600 19.950 ;
        RECT 17.440 19.780 17.610 19.950 ;
        RECT 17.800 19.780 17.970 19.950 ;
        RECT 18.460 19.780 18.630 19.950 ;
        RECT 18.900 19.780 19.070 19.950 ;
        RECT 19.340 19.780 19.510 19.950 ;
        RECT 19.750 19.780 19.920 19.950 ;
        RECT 21.760 19.780 21.930 19.950 ;
        RECT 22.120 19.780 22.290 19.950 ;
        RECT 22.780 19.780 22.950 19.950 ;
        RECT 23.220 19.780 23.390 19.950 ;
        RECT 23.660 19.780 23.830 19.950 ;
        RECT 24.070 19.780 24.240 19.950 ;
        RECT 25.030 19.780 25.200 19.950 ;
        RECT 25.390 19.780 25.560 19.950 ;
        RECT 25.750 19.780 25.920 19.950 ;
        RECT 26.110 19.780 26.280 19.950 ;
        RECT 27.100 19.780 27.270 19.950 ;
        RECT 27.540 19.780 27.710 19.950 ;
        RECT 27.980 19.780 28.150 19.950 ;
        RECT 28.390 19.780 28.560 19.950 ;
        RECT 29.350 19.780 29.520 19.950 ;
        RECT 29.710 19.780 29.880 19.950 ;
        RECT 30.070 19.780 30.240 19.950 ;
        RECT 30.430 19.780 30.600 19.950 ;
        RECT 31.420 19.780 31.590 19.950 ;
        RECT 31.860 19.780 32.030 19.950 ;
        RECT 32.300 19.780 32.470 19.950 ;
        RECT 32.710 19.780 32.880 19.950 ;
        RECT 33.670 19.780 33.840 19.950 ;
        RECT 34.030 19.780 34.200 19.950 ;
        RECT 34.390 19.780 34.560 19.950 ;
        RECT 34.750 19.780 34.920 19.950 ;
        RECT 35.740 19.780 35.910 19.950 ;
        RECT 36.180 19.780 36.350 19.950 ;
        RECT 36.620 19.780 36.790 19.950 ;
        RECT 37.030 19.780 37.200 19.950 ;
        RECT 38.040 19.780 38.210 19.950 ;
        RECT 38.400 19.780 38.570 19.950 ;
        RECT 39.580 19.780 39.750 19.950 ;
        RECT 40.020 19.780 40.190 19.950 ;
        RECT 40.460 19.780 40.630 19.950 ;
        RECT 40.870 19.780 41.040 19.950 ;
        RECT 41.830 19.780 42.000 19.950 ;
        RECT 42.190 19.780 42.360 19.950 ;
        RECT 42.550 19.780 42.720 19.950 ;
        RECT 42.910 19.780 43.080 19.950 ;
        RECT 43.900 19.780 44.070 19.950 ;
        RECT 44.340 19.780 44.510 19.950 ;
        RECT 44.780 19.780 44.950 19.950 ;
        RECT 45.190 19.780 45.360 19.950 ;
        RECT 45.720 19.780 45.890 19.950 ;
        RECT 46.080 19.780 46.250 19.950 ;
        RECT 46.990 19.780 47.160 19.950 ;
        RECT 47.350 19.780 47.520 19.950 ;
        RECT 47.710 19.780 47.880 19.950 ;
        RECT 49.180 19.780 49.350 19.950 ;
        RECT 49.620 19.780 49.790 19.950 ;
        RECT 50.060 19.780 50.230 19.950 ;
        RECT 50.470 19.780 50.640 19.950 ;
        RECT 51.000 19.780 51.170 19.950 ;
        RECT 51.360 19.780 51.530 19.950 ;
        RECT 52.270 19.780 52.440 19.950 ;
        RECT 52.630 19.780 52.800 19.950 ;
        RECT 52.990 19.780 53.160 19.950 ;
        RECT 54.460 19.780 54.630 19.950 ;
        RECT 54.900 19.780 55.070 19.950 ;
        RECT 55.340 19.780 55.510 19.950 ;
        RECT 55.750 19.780 55.920 19.950 ;
        RECT 56.280 19.780 56.450 19.950 ;
        RECT 56.640 19.780 56.810 19.950 ;
        RECT 57.820 19.780 57.990 19.950 ;
        RECT 58.260 19.780 58.430 19.950 ;
        RECT 58.700 19.780 58.870 19.950 ;
        RECT 59.110 19.780 59.280 19.950 ;
        RECT 59.640 19.780 59.810 19.950 ;
        RECT 60.000 19.780 60.170 19.950 ;
        RECT 60.360 19.780 60.530 19.950 ;
        RECT 61.200 19.780 61.370 19.950 ;
        RECT 61.560 19.780 61.730 19.950 ;
        RECT 61.920 19.780 62.090 19.950 ;
        RECT 62.760 19.780 62.930 19.950 ;
        RECT 63.120 19.780 63.290 19.950 ;
        RECT 63.480 19.780 63.650 19.950 ;
        RECT 64.540 19.780 64.710 19.950 ;
        RECT 64.980 19.780 65.150 19.950 ;
        RECT 65.420 19.780 65.590 19.950 ;
        RECT 65.830 19.780 66.000 19.950 ;
        RECT 68.440 19.780 68.610 19.950 ;
        RECT 68.800 19.780 68.970 19.950 ;
        RECT 69.160 19.780 69.330 19.950 ;
        RECT 70.300 19.780 70.470 19.950 ;
        RECT 70.740 19.780 70.910 19.950 ;
        RECT 71.180 19.780 71.350 19.950 ;
        RECT 71.590 19.780 71.760 19.950 ;
        RECT 72.550 19.780 72.720 19.950 ;
        RECT 72.910 19.780 73.080 19.950 ;
        RECT 73.270 19.780 73.440 19.950 ;
        RECT 73.630 19.780 73.800 19.950 ;
        RECT 74.620 19.780 74.790 19.950 ;
        RECT 75.060 19.780 75.230 19.950 ;
        RECT 75.500 19.780 75.670 19.950 ;
        RECT 75.910 19.780 76.080 19.950 ;
        RECT 76.870 19.780 77.040 19.950 ;
        RECT 77.230 19.780 77.400 19.950 ;
        RECT 77.590 19.780 77.760 19.950 ;
        RECT 77.950 19.780 78.120 19.950 ;
        RECT 79.470 19.790 79.640 19.960 ;
        RECT 79.910 19.790 80.080 19.960 ;
        RECT 80.320 19.790 80.490 19.960 ;
        RECT 80.750 19.790 80.920 19.960 ;
        RECT 81.190 19.790 81.360 19.960 ;
        RECT 81.600 19.790 81.770 19.960 ;
        RECT 83.150 19.780 83.320 19.950 ;
        RECT 83.510 19.780 83.680 19.950 ;
        RECT 83.870 19.780 84.040 19.950 ;
        RECT 84.790 19.780 84.960 19.950 ;
        RECT 85.150 19.780 85.320 19.950 ;
        RECT 89.750 19.780 89.920 19.950 ;
        RECT 90.110 19.780 90.280 19.950 ;
        RECT 90.470 19.780 90.640 19.950 ;
        RECT 93.720 19.780 93.890 19.950 ;
        RECT 94.080 19.780 94.250 19.950 ;
        RECT 94.440 19.780 94.610 19.950 ;
        RECT 96.330 19.780 96.500 19.950 ;
        RECT 96.690 19.780 96.860 19.950 ;
        RECT 97.050 19.780 97.220 19.950 ;
        RECT 98.670 19.790 98.840 19.960 ;
        RECT 99.110 19.790 99.280 19.960 ;
        RECT 99.520 19.790 99.690 19.960 ;
        RECT 99.950 19.790 100.120 19.960 ;
        RECT 100.390 19.790 100.560 19.960 ;
        RECT 100.800 19.790 100.970 19.960 ;
        RECT 103.310 19.780 103.480 19.950 ;
        RECT 103.670 19.780 103.840 19.950 ;
        RECT 104.030 19.780 104.200 19.950 ;
        RECT 104.950 19.780 105.120 19.950 ;
        RECT 105.310 19.780 105.480 19.950 ;
        RECT 109.910 19.780 110.080 19.950 ;
        RECT 110.270 19.780 110.440 19.950 ;
        RECT 110.630 19.780 110.800 19.950 ;
        RECT 113.880 19.780 114.050 19.950 ;
        RECT 114.240 19.780 114.410 19.950 ;
        RECT 114.600 19.780 114.770 19.950 ;
        RECT 116.490 19.780 116.660 19.950 ;
        RECT 116.850 19.780 117.020 19.950 ;
        RECT 117.210 19.780 117.380 19.950 ;
        RECT 118.300 19.780 118.470 19.950 ;
        RECT 118.740 19.780 118.910 19.950 ;
        RECT 119.180 19.780 119.350 19.950 ;
        RECT 119.590 19.780 119.760 19.950 ;
        RECT 121.600 19.780 121.770 19.950 ;
        RECT 121.960 19.780 122.130 19.950 ;
        RECT 122.620 19.780 122.790 19.950 ;
        RECT 123.060 19.780 123.230 19.950 ;
        RECT 123.500 19.780 123.670 19.950 ;
        RECT 123.910 19.780 124.080 19.950 ;
        RECT 125.920 19.780 126.090 19.950 ;
        RECT 126.280 19.780 126.450 19.950 ;
        RECT 127.470 19.790 127.640 19.960 ;
        RECT 127.910 19.790 128.080 19.960 ;
        RECT 128.320 19.790 128.490 19.960 ;
        RECT 128.750 19.790 128.920 19.960 ;
        RECT 129.190 19.790 129.360 19.960 ;
        RECT 129.600 19.790 129.770 19.960 ;
        RECT 131.310 19.790 131.480 19.960 ;
        RECT 131.750 19.790 131.920 19.960 ;
        RECT 132.160 19.790 132.330 19.960 ;
        RECT 132.590 19.790 132.760 19.960 ;
        RECT 133.030 19.790 133.200 19.960 ;
        RECT 133.440 19.790 133.610 19.960 ;
        RECT 136.000 19.780 136.170 19.950 ;
        RECT 136.360 19.780 136.530 19.950 ;
        RECT 137.550 19.790 137.720 19.960 ;
        RECT 137.990 19.790 138.160 19.960 ;
        RECT 138.400 19.790 138.570 19.960 ;
        RECT 138.830 19.790 139.000 19.960 ;
        RECT 139.270 19.790 139.440 19.960 ;
        RECT 139.680 19.790 139.850 19.960 ;
      LAYER L1M1_PR_C ;
        RECT 141.760 150.500 141.930 150.680 ;
        RECT 17.920 142.360 18.090 142.540 ;
        RECT 36.160 142.360 36.330 142.540 ;
        RECT 43.840 142.360 44.010 142.540 ;
        RECT 85.600 142.360 85.770 142.540 ;
        RECT 141.760 142.360 141.930 142.540 ;
        RECT 30.400 134.220 30.570 134.400 ;
        RECT 62.560 134.220 62.730 134.400 ;
        RECT 75.040 134.220 75.210 134.400 ;
        RECT 98.080 134.220 98.250 134.400 ;
        RECT 109.600 134.220 109.770 134.400 ;
        RECT 141.760 134.220 141.930 134.400 ;
        RECT 34.240 126.080 34.410 126.260 ;
        RECT 43.840 126.080 44.010 126.260 ;
        RECT 74.080 126.080 74.250 126.260 ;
        RECT 110.560 126.080 110.730 126.260 ;
        RECT 118.240 126.080 118.410 126.260 ;
        RECT 10.720 117.940 10.890 118.120 ;
        RECT 28.480 117.940 28.650 118.120 ;
        RECT 43.360 117.940 43.530 118.120 ;
        RECT 50.080 117.940 50.250 118.120 ;
        RECT 67.360 117.940 67.530 118.120 ;
        RECT 100.480 117.940 100.650 118.120 ;
        RECT 141.760 117.940 141.930 118.120 ;
        RECT 24.160 109.800 24.330 109.980 ;
        RECT 37.120 109.800 37.290 109.980 ;
        RECT 71.680 109.800 71.850 109.980 ;
        RECT 40.480 101.660 40.650 101.840 ;
        RECT 61.120 101.660 61.290 101.840 ;
        RECT 121.120 101.660 121.290 101.840 ;
        RECT 32.800 93.520 32.970 93.700 ;
        RECT 74.080 93.520 74.250 93.700 ;
        RECT 98.560 93.520 98.730 93.700 ;
        RECT 121.120 93.520 121.290 93.700 ;
        RECT 20.320 85.380 20.490 85.560 ;
        RECT 68.320 85.380 68.490 85.560 ;
        RECT 101.440 85.380 101.610 85.560 ;
        RECT 117.760 85.380 117.930 85.560 ;
        RECT 134.080 85.380 134.250 85.560 ;
        RECT 141.760 85.380 141.930 85.560 ;
        RECT 14.560 77.240 14.730 77.420 ;
        RECT 71.200 77.240 71.370 77.420 ;
        RECT 80.800 77.240 80.970 77.420 ;
        RECT 47.680 69.100 47.850 69.280 ;
        RECT 59.200 69.100 59.370 69.280 ;
        RECT 76.480 69.100 76.650 69.280 ;
        RECT 91.360 60.960 91.530 61.140 ;
        RECT 105.760 60.960 105.930 61.140 ;
        RECT 141.760 60.960 141.930 61.140 ;
        RECT 7.840 52.820 8.010 53.000 ;
        RECT 47.680 52.820 47.850 53.000 ;
        RECT 81.280 52.820 81.450 53.000 ;
        RECT 107.200 52.820 107.370 53.000 ;
        RECT 123.040 52.820 123.210 53.000 ;
        RECT 50.560 44.680 50.730 44.860 ;
        RECT 94.720 44.680 94.890 44.860 ;
        RECT 108.160 44.680 108.330 44.860 ;
        RECT 14.560 36.540 14.730 36.720 ;
        RECT 77.920 36.540 78.090 36.720 ;
        RECT 110.560 36.540 110.730 36.720 ;
        RECT 104.320 28.400 104.490 28.580 ;
        RECT 119.680 28.400 119.850 28.580 ;
        RECT 132.160 28.400 132.330 28.580 ;
        RECT 141.760 28.400 141.930 28.580 ;
      LAYER met1 ;
        RECT 5.760 149.960 142.080 150.840 ;
        RECT 5.760 141.820 142.080 142.700 ;
        RECT 5.760 133.680 142.080 134.560 ;
        RECT 5.760 125.540 142.080 126.420 ;
        RECT 5.760 117.400 142.080 118.280 ;
        RECT 5.760 109.260 142.080 110.140 ;
        RECT 5.760 101.120 142.080 102.000 ;
        RECT 5.760 92.980 142.080 93.860 ;
        RECT 5.760 84.840 142.080 85.720 ;
        RECT 5.760 76.700 142.080 77.580 ;
        RECT 5.760 68.560 142.080 69.440 ;
        RECT 5.760 60.420 142.080 61.300 ;
        RECT 5.760 52.280 142.080 53.160 ;
        RECT 5.760 44.140 142.080 45.020 ;
        RECT 5.760 36.000 142.080 36.880 ;
        RECT 5.760 27.860 142.080 28.740 ;
        RECT 5.760 19.720 142.080 20.600 ;
      LAYER via ;
        RECT 50.590 150.460 50.850 150.720 ;
        RECT 50.910 150.460 51.170 150.720 ;
        RECT 51.230 150.460 51.490 150.720 ;
        RECT 51.550 150.460 51.810 150.720 ;
        RECT 96.030 150.460 96.290 150.720 ;
        RECT 96.350 150.460 96.610 150.720 ;
        RECT 96.670 150.460 96.930 150.720 ;
        RECT 96.990 150.460 97.250 150.720 ;
        RECT 50.590 142.320 50.850 142.580 ;
        RECT 50.910 142.320 51.170 142.580 ;
        RECT 51.230 142.320 51.490 142.580 ;
        RECT 51.550 142.320 51.810 142.580 ;
        RECT 96.030 142.320 96.290 142.580 ;
        RECT 96.350 142.320 96.610 142.580 ;
        RECT 96.670 142.320 96.930 142.580 ;
        RECT 96.990 142.320 97.250 142.580 ;
        RECT 50.590 134.180 50.850 134.440 ;
        RECT 50.910 134.180 51.170 134.440 ;
        RECT 51.230 134.180 51.490 134.440 ;
        RECT 51.550 134.180 51.810 134.440 ;
        RECT 96.030 134.180 96.290 134.440 ;
        RECT 96.350 134.180 96.610 134.440 ;
        RECT 96.670 134.180 96.930 134.440 ;
        RECT 96.990 134.180 97.250 134.440 ;
        RECT 50.590 126.040 50.850 126.300 ;
        RECT 50.910 126.040 51.170 126.300 ;
        RECT 51.230 126.040 51.490 126.300 ;
        RECT 51.550 126.040 51.810 126.300 ;
        RECT 96.030 126.040 96.290 126.300 ;
        RECT 96.350 126.040 96.610 126.300 ;
        RECT 96.670 126.040 96.930 126.300 ;
        RECT 96.990 126.040 97.250 126.300 ;
        RECT 50.590 117.900 50.850 118.160 ;
        RECT 50.910 117.900 51.170 118.160 ;
        RECT 51.230 117.900 51.490 118.160 ;
        RECT 51.550 117.900 51.810 118.160 ;
        RECT 96.030 117.900 96.290 118.160 ;
        RECT 96.350 117.900 96.610 118.160 ;
        RECT 96.670 117.900 96.930 118.160 ;
        RECT 96.990 117.900 97.250 118.160 ;
        RECT 50.590 109.760 50.850 110.020 ;
        RECT 50.910 109.760 51.170 110.020 ;
        RECT 51.230 109.760 51.490 110.020 ;
        RECT 51.550 109.760 51.810 110.020 ;
        RECT 96.030 109.760 96.290 110.020 ;
        RECT 96.350 109.760 96.610 110.020 ;
        RECT 96.670 109.760 96.930 110.020 ;
        RECT 96.990 109.760 97.250 110.020 ;
        RECT 50.590 101.620 50.850 101.880 ;
        RECT 50.910 101.620 51.170 101.880 ;
        RECT 51.230 101.620 51.490 101.880 ;
        RECT 51.550 101.620 51.810 101.880 ;
        RECT 96.030 101.620 96.290 101.880 ;
        RECT 96.350 101.620 96.610 101.880 ;
        RECT 96.670 101.620 96.930 101.880 ;
        RECT 96.990 101.620 97.250 101.880 ;
        RECT 50.590 93.480 50.850 93.740 ;
        RECT 50.910 93.480 51.170 93.740 ;
        RECT 51.230 93.480 51.490 93.740 ;
        RECT 51.550 93.480 51.810 93.740 ;
        RECT 96.030 93.480 96.290 93.740 ;
        RECT 96.350 93.480 96.610 93.740 ;
        RECT 96.670 93.480 96.930 93.740 ;
        RECT 96.990 93.480 97.250 93.740 ;
        RECT 50.590 85.340 50.850 85.600 ;
        RECT 50.910 85.340 51.170 85.600 ;
        RECT 51.230 85.340 51.490 85.600 ;
        RECT 51.550 85.340 51.810 85.600 ;
        RECT 96.030 85.340 96.290 85.600 ;
        RECT 96.350 85.340 96.610 85.600 ;
        RECT 96.670 85.340 96.930 85.600 ;
        RECT 96.990 85.340 97.250 85.600 ;
        RECT 50.590 77.200 50.850 77.460 ;
        RECT 50.910 77.200 51.170 77.460 ;
        RECT 51.230 77.200 51.490 77.460 ;
        RECT 51.550 77.200 51.810 77.460 ;
        RECT 96.030 77.200 96.290 77.460 ;
        RECT 96.350 77.200 96.610 77.460 ;
        RECT 96.670 77.200 96.930 77.460 ;
        RECT 96.990 77.200 97.250 77.460 ;
        RECT 50.590 69.060 50.850 69.320 ;
        RECT 50.910 69.060 51.170 69.320 ;
        RECT 51.230 69.060 51.490 69.320 ;
        RECT 51.550 69.060 51.810 69.320 ;
        RECT 96.030 69.060 96.290 69.320 ;
        RECT 96.350 69.060 96.610 69.320 ;
        RECT 96.670 69.060 96.930 69.320 ;
        RECT 96.990 69.060 97.250 69.320 ;
        RECT 50.590 60.920 50.850 61.180 ;
        RECT 50.910 60.920 51.170 61.180 ;
        RECT 51.230 60.920 51.490 61.180 ;
        RECT 51.550 60.920 51.810 61.180 ;
        RECT 96.030 60.920 96.290 61.180 ;
        RECT 96.350 60.920 96.610 61.180 ;
        RECT 96.670 60.920 96.930 61.180 ;
        RECT 96.990 60.920 97.250 61.180 ;
        RECT 50.590 52.780 50.850 53.040 ;
        RECT 50.910 52.780 51.170 53.040 ;
        RECT 51.230 52.780 51.490 53.040 ;
        RECT 51.550 52.780 51.810 53.040 ;
        RECT 96.030 52.780 96.290 53.040 ;
        RECT 96.350 52.780 96.610 53.040 ;
        RECT 96.670 52.780 96.930 53.040 ;
        RECT 96.990 52.780 97.250 53.040 ;
        RECT 50.590 44.640 50.850 44.900 ;
        RECT 50.910 44.640 51.170 44.900 ;
        RECT 51.230 44.640 51.490 44.900 ;
        RECT 51.550 44.640 51.810 44.900 ;
        RECT 96.030 44.640 96.290 44.900 ;
        RECT 96.350 44.640 96.610 44.900 ;
        RECT 96.670 44.640 96.930 44.900 ;
        RECT 96.990 44.640 97.250 44.900 ;
        RECT 50.590 36.500 50.850 36.760 ;
        RECT 50.910 36.500 51.170 36.760 ;
        RECT 51.230 36.500 51.490 36.760 ;
        RECT 51.550 36.500 51.810 36.760 ;
        RECT 96.030 36.500 96.290 36.760 ;
        RECT 96.350 36.500 96.610 36.760 ;
        RECT 96.670 36.500 96.930 36.760 ;
        RECT 96.990 36.500 97.250 36.760 ;
        RECT 50.590 28.360 50.850 28.620 ;
        RECT 50.910 28.360 51.170 28.620 ;
        RECT 51.230 28.360 51.490 28.620 ;
        RECT 51.550 28.360 51.810 28.620 ;
        RECT 96.030 28.360 96.290 28.620 ;
        RECT 96.350 28.360 96.610 28.620 ;
        RECT 96.670 28.360 96.930 28.620 ;
        RECT 96.990 28.360 97.250 28.620 ;
        RECT 50.590 20.220 50.850 20.480 ;
        RECT 50.910 20.220 51.170 20.480 ;
        RECT 51.230 20.220 51.490 20.480 ;
        RECT 51.550 20.220 51.810 20.480 ;
        RECT 96.030 20.220 96.290 20.480 ;
        RECT 96.350 20.220 96.610 20.480 ;
        RECT 96.670 20.220 96.930 20.480 ;
        RECT 96.990 20.220 97.250 20.480 ;
      LAYER met2 ;
        RECT 50.460 150.330 51.940 150.840 ;
        RECT 95.900 150.330 97.380 150.840 ;
        RECT 50.460 142.190 51.940 142.700 ;
        RECT 95.900 142.190 97.380 142.700 ;
        RECT 50.460 134.050 51.940 134.560 ;
        RECT 95.900 134.050 97.380 134.560 ;
        RECT 50.460 125.910 51.940 126.420 ;
        RECT 95.900 125.910 97.380 126.420 ;
        RECT 50.460 117.770 51.940 118.280 ;
        RECT 95.900 117.770 97.380 118.280 ;
        RECT 50.460 109.630 51.940 110.140 ;
        RECT 95.900 109.630 97.380 110.140 ;
        RECT 50.460 101.490 51.940 102.000 ;
        RECT 95.900 101.490 97.380 102.000 ;
        RECT 50.460 93.350 51.940 93.860 ;
        RECT 95.900 93.350 97.380 93.860 ;
        RECT 50.460 85.210 51.940 85.720 ;
        RECT 95.900 85.210 97.380 85.720 ;
        RECT 50.460 77.070 51.940 77.580 ;
        RECT 95.900 77.070 97.380 77.580 ;
        RECT 50.460 68.930 51.940 69.440 ;
        RECT 95.900 68.930 97.380 69.440 ;
        RECT 50.460 60.790 51.940 61.300 ;
        RECT 95.900 60.790 97.380 61.300 ;
        RECT 50.460 52.650 51.940 53.160 ;
        RECT 95.900 52.650 97.380 53.160 ;
        RECT 50.460 44.510 51.940 45.020 ;
        RECT 95.900 44.510 97.380 45.020 ;
        RECT 50.460 36.370 51.940 36.880 ;
        RECT 95.900 36.370 97.380 36.880 ;
        RECT 50.460 28.230 51.940 28.740 ;
        RECT 95.900 28.230 97.380 28.740 ;
        RECT 50.460 20.090 51.940 20.600 ;
        RECT 95.900 20.090 97.380 20.600 ;
      LAYER via2 ;
        RECT 50.460 150.450 50.740 150.730 ;
        RECT 50.860 150.450 51.140 150.730 ;
        RECT 51.260 150.450 51.540 150.730 ;
        RECT 51.660 150.450 51.940 150.730 ;
        RECT 95.900 150.450 96.180 150.730 ;
        RECT 96.300 150.450 96.580 150.730 ;
        RECT 96.700 150.450 96.980 150.730 ;
        RECT 97.100 150.450 97.380 150.730 ;
        RECT 50.460 142.310 50.740 142.590 ;
        RECT 50.860 142.310 51.140 142.590 ;
        RECT 51.260 142.310 51.540 142.590 ;
        RECT 51.660 142.310 51.940 142.590 ;
        RECT 95.900 142.310 96.180 142.590 ;
        RECT 96.300 142.310 96.580 142.590 ;
        RECT 96.700 142.310 96.980 142.590 ;
        RECT 97.100 142.310 97.380 142.590 ;
        RECT 50.460 134.170 50.740 134.450 ;
        RECT 50.860 134.170 51.140 134.450 ;
        RECT 51.260 134.170 51.540 134.450 ;
        RECT 51.660 134.170 51.940 134.450 ;
        RECT 95.900 134.170 96.180 134.450 ;
        RECT 96.300 134.170 96.580 134.450 ;
        RECT 96.700 134.170 96.980 134.450 ;
        RECT 97.100 134.170 97.380 134.450 ;
        RECT 50.460 126.030 50.740 126.310 ;
        RECT 50.860 126.030 51.140 126.310 ;
        RECT 51.260 126.030 51.540 126.310 ;
        RECT 51.660 126.030 51.940 126.310 ;
        RECT 95.900 126.030 96.180 126.310 ;
        RECT 96.300 126.030 96.580 126.310 ;
        RECT 96.700 126.030 96.980 126.310 ;
        RECT 97.100 126.030 97.380 126.310 ;
        RECT 50.460 117.890 50.740 118.170 ;
        RECT 50.860 117.890 51.140 118.170 ;
        RECT 51.260 117.890 51.540 118.170 ;
        RECT 51.660 117.890 51.940 118.170 ;
        RECT 95.900 117.890 96.180 118.170 ;
        RECT 96.300 117.890 96.580 118.170 ;
        RECT 96.700 117.890 96.980 118.170 ;
        RECT 97.100 117.890 97.380 118.170 ;
        RECT 50.460 109.750 50.740 110.030 ;
        RECT 50.860 109.750 51.140 110.030 ;
        RECT 51.260 109.750 51.540 110.030 ;
        RECT 51.660 109.750 51.940 110.030 ;
        RECT 95.900 109.750 96.180 110.030 ;
        RECT 96.300 109.750 96.580 110.030 ;
        RECT 96.700 109.750 96.980 110.030 ;
        RECT 97.100 109.750 97.380 110.030 ;
        RECT 50.460 101.610 50.740 101.890 ;
        RECT 50.860 101.610 51.140 101.890 ;
        RECT 51.260 101.610 51.540 101.890 ;
        RECT 51.660 101.610 51.940 101.890 ;
        RECT 95.900 101.610 96.180 101.890 ;
        RECT 96.300 101.610 96.580 101.890 ;
        RECT 96.700 101.610 96.980 101.890 ;
        RECT 97.100 101.610 97.380 101.890 ;
        RECT 50.460 93.470 50.740 93.750 ;
        RECT 50.860 93.470 51.140 93.750 ;
        RECT 51.260 93.470 51.540 93.750 ;
        RECT 51.660 93.470 51.940 93.750 ;
        RECT 95.900 93.470 96.180 93.750 ;
        RECT 96.300 93.470 96.580 93.750 ;
        RECT 96.700 93.470 96.980 93.750 ;
        RECT 97.100 93.470 97.380 93.750 ;
        RECT 50.460 85.330 50.740 85.610 ;
        RECT 50.860 85.330 51.140 85.610 ;
        RECT 51.260 85.330 51.540 85.610 ;
        RECT 51.660 85.330 51.940 85.610 ;
        RECT 95.900 85.330 96.180 85.610 ;
        RECT 96.300 85.330 96.580 85.610 ;
        RECT 96.700 85.330 96.980 85.610 ;
        RECT 97.100 85.330 97.380 85.610 ;
        RECT 50.460 77.190 50.740 77.470 ;
        RECT 50.860 77.190 51.140 77.470 ;
        RECT 51.260 77.190 51.540 77.470 ;
        RECT 51.660 77.190 51.940 77.470 ;
        RECT 95.900 77.190 96.180 77.470 ;
        RECT 96.300 77.190 96.580 77.470 ;
        RECT 96.700 77.190 96.980 77.470 ;
        RECT 97.100 77.190 97.380 77.470 ;
        RECT 50.460 69.050 50.740 69.330 ;
        RECT 50.860 69.050 51.140 69.330 ;
        RECT 51.260 69.050 51.540 69.330 ;
        RECT 51.660 69.050 51.940 69.330 ;
        RECT 95.900 69.050 96.180 69.330 ;
        RECT 96.300 69.050 96.580 69.330 ;
        RECT 96.700 69.050 96.980 69.330 ;
        RECT 97.100 69.050 97.380 69.330 ;
        RECT 50.460 60.910 50.740 61.190 ;
        RECT 50.860 60.910 51.140 61.190 ;
        RECT 51.260 60.910 51.540 61.190 ;
        RECT 51.660 60.910 51.940 61.190 ;
        RECT 95.900 60.910 96.180 61.190 ;
        RECT 96.300 60.910 96.580 61.190 ;
        RECT 96.700 60.910 96.980 61.190 ;
        RECT 97.100 60.910 97.380 61.190 ;
        RECT 50.460 52.770 50.740 53.050 ;
        RECT 50.860 52.770 51.140 53.050 ;
        RECT 51.260 52.770 51.540 53.050 ;
        RECT 51.660 52.770 51.940 53.050 ;
        RECT 95.900 52.770 96.180 53.050 ;
        RECT 96.300 52.770 96.580 53.050 ;
        RECT 96.700 52.770 96.980 53.050 ;
        RECT 97.100 52.770 97.380 53.050 ;
        RECT 50.460 44.630 50.740 44.910 ;
        RECT 50.860 44.630 51.140 44.910 ;
        RECT 51.260 44.630 51.540 44.910 ;
        RECT 51.660 44.630 51.940 44.910 ;
        RECT 95.900 44.630 96.180 44.910 ;
        RECT 96.300 44.630 96.580 44.910 ;
        RECT 96.700 44.630 96.980 44.910 ;
        RECT 97.100 44.630 97.380 44.910 ;
        RECT 50.460 36.490 50.740 36.770 ;
        RECT 50.860 36.490 51.140 36.770 ;
        RECT 51.260 36.490 51.540 36.770 ;
        RECT 51.660 36.490 51.940 36.770 ;
        RECT 95.900 36.490 96.180 36.770 ;
        RECT 96.300 36.490 96.580 36.770 ;
        RECT 96.700 36.490 96.980 36.770 ;
        RECT 97.100 36.490 97.380 36.770 ;
        RECT 50.460 28.350 50.740 28.630 ;
        RECT 50.860 28.350 51.140 28.630 ;
        RECT 51.260 28.350 51.540 28.630 ;
        RECT 51.660 28.350 51.940 28.630 ;
        RECT 95.900 28.350 96.180 28.630 ;
        RECT 96.300 28.350 96.580 28.630 ;
        RECT 96.700 28.350 96.980 28.630 ;
        RECT 97.100 28.350 97.380 28.630 ;
        RECT 50.460 20.210 50.740 20.490 ;
        RECT 50.860 20.210 51.140 20.490 ;
        RECT 51.260 20.210 51.540 20.490 ;
        RECT 51.660 20.210 51.940 20.490 ;
        RECT 95.900 20.210 96.180 20.490 ;
        RECT 96.300 20.210 96.580 20.490 ;
        RECT 96.700 20.210 96.980 20.490 ;
        RECT 97.100 20.210 97.380 20.490 ;
      LAYER met3 ;
        RECT 50.400 150.420 52.000 150.750 ;
        RECT 95.840 150.420 97.440 150.750 ;
        RECT 50.400 142.280 52.000 142.610 ;
        RECT 95.840 142.280 97.440 142.610 ;
        RECT 50.400 134.140 52.000 134.470 ;
        RECT 95.840 134.140 97.440 134.470 ;
        RECT 50.400 126.000 52.000 126.330 ;
        RECT 95.840 126.000 97.440 126.330 ;
        RECT 50.400 117.860 52.000 118.190 ;
        RECT 95.840 117.860 97.440 118.190 ;
        RECT 50.400 109.720 52.000 110.050 ;
        RECT 95.840 109.720 97.440 110.050 ;
        RECT 50.400 101.580 52.000 101.910 ;
        RECT 95.840 101.580 97.440 101.910 ;
        RECT 50.400 93.440 52.000 93.770 ;
        RECT 95.840 93.440 97.440 93.770 ;
        RECT 50.400 85.300 52.000 85.630 ;
        RECT 95.840 85.300 97.440 85.630 ;
        RECT 50.400 77.160 52.000 77.490 ;
        RECT 95.840 77.160 97.440 77.490 ;
        RECT 50.400 69.020 52.000 69.350 ;
        RECT 95.840 69.020 97.440 69.350 ;
        RECT 50.400 60.880 52.000 61.210 ;
        RECT 95.840 60.880 97.440 61.210 ;
        RECT 50.400 52.740 52.000 53.070 ;
        RECT 95.840 52.740 97.440 53.070 ;
        RECT 50.400 44.600 52.000 44.930 ;
        RECT 95.840 44.600 97.440 44.930 ;
        RECT 50.400 36.460 52.000 36.790 ;
        RECT 95.840 36.460 97.440 36.790 ;
        RECT 50.400 28.320 52.000 28.650 ;
        RECT 95.840 28.320 97.440 28.650 ;
        RECT 50.400 20.180 52.000 20.510 ;
        RECT 95.840 20.180 97.440 20.510 ;
      LAYER via3 ;
        RECT 50.440 150.430 50.760 150.750 ;
        RECT 50.840 150.430 51.160 150.750 ;
        RECT 51.240 150.430 51.560 150.750 ;
        RECT 51.640 150.430 51.960 150.750 ;
        RECT 95.880 150.430 96.200 150.750 ;
        RECT 96.280 150.430 96.600 150.750 ;
        RECT 96.680 150.430 97.000 150.750 ;
        RECT 97.080 150.430 97.400 150.750 ;
        RECT 50.440 142.290 50.760 142.610 ;
        RECT 50.840 142.290 51.160 142.610 ;
        RECT 51.240 142.290 51.560 142.610 ;
        RECT 51.640 142.290 51.960 142.610 ;
        RECT 95.880 142.290 96.200 142.610 ;
        RECT 96.280 142.290 96.600 142.610 ;
        RECT 96.680 142.290 97.000 142.610 ;
        RECT 97.080 142.290 97.400 142.610 ;
        RECT 50.440 134.150 50.760 134.470 ;
        RECT 50.840 134.150 51.160 134.470 ;
        RECT 51.240 134.150 51.560 134.470 ;
        RECT 51.640 134.150 51.960 134.470 ;
        RECT 95.880 134.150 96.200 134.470 ;
        RECT 96.280 134.150 96.600 134.470 ;
        RECT 96.680 134.150 97.000 134.470 ;
        RECT 97.080 134.150 97.400 134.470 ;
        RECT 50.440 126.010 50.760 126.330 ;
        RECT 50.840 126.010 51.160 126.330 ;
        RECT 51.240 126.010 51.560 126.330 ;
        RECT 51.640 126.010 51.960 126.330 ;
        RECT 95.880 126.010 96.200 126.330 ;
        RECT 96.280 126.010 96.600 126.330 ;
        RECT 96.680 126.010 97.000 126.330 ;
        RECT 97.080 126.010 97.400 126.330 ;
        RECT 50.440 117.870 50.760 118.190 ;
        RECT 50.840 117.870 51.160 118.190 ;
        RECT 51.240 117.870 51.560 118.190 ;
        RECT 51.640 117.870 51.960 118.190 ;
        RECT 95.880 117.870 96.200 118.190 ;
        RECT 96.280 117.870 96.600 118.190 ;
        RECT 96.680 117.870 97.000 118.190 ;
        RECT 97.080 117.870 97.400 118.190 ;
        RECT 50.440 109.730 50.760 110.050 ;
        RECT 50.840 109.730 51.160 110.050 ;
        RECT 51.240 109.730 51.560 110.050 ;
        RECT 51.640 109.730 51.960 110.050 ;
        RECT 95.880 109.730 96.200 110.050 ;
        RECT 96.280 109.730 96.600 110.050 ;
        RECT 96.680 109.730 97.000 110.050 ;
        RECT 97.080 109.730 97.400 110.050 ;
        RECT 50.440 101.590 50.760 101.910 ;
        RECT 50.840 101.590 51.160 101.910 ;
        RECT 51.240 101.590 51.560 101.910 ;
        RECT 51.640 101.590 51.960 101.910 ;
        RECT 95.880 101.590 96.200 101.910 ;
        RECT 96.280 101.590 96.600 101.910 ;
        RECT 96.680 101.590 97.000 101.910 ;
        RECT 97.080 101.590 97.400 101.910 ;
        RECT 50.440 93.450 50.760 93.770 ;
        RECT 50.840 93.450 51.160 93.770 ;
        RECT 51.240 93.450 51.560 93.770 ;
        RECT 51.640 93.450 51.960 93.770 ;
        RECT 95.880 93.450 96.200 93.770 ;
        RECT 96.280 93.450 96.600 93.770 ;
        RECT 96.680 93.450 97.000 93.770 ;
        RECT 97.080 93.450 97.400 93.770 ;
        RECT 50.440 85.310 50.760 85.630 ;
        RECT 50.840 85.310 51.160 85.630 ;
        RECT 51.240 85.310 51.560 85.630 ;
        RECT 51.640 85.310 51.960 85.630 ;
        RECT 95.880 85.310 96.200 85.630 ;
        RECT 96.280 85.310 96.600 85.630 ;
        RECT 96.680 85.310 97.000 85.630 ;
        RECT 97.080 85.310 97.400 85.630 ;
        RECT 50.440 77.170 50.760 77.490 ;
        RECT 50.840 77.170 51.160 77.490 ;
        RECT 51.240 77.170 51.560 77.490 ;
        RECT 51.640 77.170 51.960 77.490 ;
        RECT 95.880 77.170 96.200 77.490 ;
        RECT 96.280 77.170 96.600 77.490 ;
        RECT 96.680 77.170 97.000 77.490 ;
        RECT 97.080 77.170 97.400 77.490 ;
        RECT 50.440 69.030 50.760 69.350 ;
        RECT 50.840 69.030 51.160 69.350 ;
        RECT 51.240 69.030 51.560 69.350 ;
        RECT 51.640 69.030 51.960 69.350 ;
        RECT 95.880 69.030 96.200 69.350 ;
        RECT 96.280 69.030 96.600 69.350 ;
        RECT 96.680 69.030 97.000 69.350 ;
        RECT 97.080 69.030 97.400 69.350 ;
        RECT 50.440 60.890 50.760 61.210 ;
        RECT 50.840 60.890 51.160 61.210 ;
        RECT 51.240 60.890 51.560 61.210 ;
        RECT 51.640 60.890 51.960 61.210 ;
        RECT 95.880 60.890 96.200 61.210 ;
        RECT 96.280 60.890 96.600 61.210 ;
        RECT 96.680 60.890 97.000 61.210 ;
        RECT 97.080 60.890 97.400 61.210 ;
        RECT 50.440 52.750 50.760 53.070 ;
        RECT 50.840 52.750 51.160 53.070 ;
        RECT 51.240 52.750 51.560 53.070 ;
        RECT 51.640 52.750 51.960 53.070 ;
        RECT 95.880 52.750 96.200 53.070 ;
        RECT 96.280 52.750 96.600 53.070 ;
        RECT 96.680 52.750 97.000 53.070 ;
        RECT 97.080 52.750 97.400 53.070 ;
        RECT 50.440 44.610 50.760 44.930 ;
        RECT 50.840 44.610 51.160 44.930 ;
        RECT 51.240 44.610 51.560 44.930 ;
        RECT 51.640 44.610 51.960 44.930 ;
        RECT 95.880 44.610 96.200 44.930 ;
        RECT 96.280 44.610 96.600 44.930 ;
        RECT 96.680 44.610 97.000 44.930 ;
        RECT 97.080 44.610 97.400 44.930 ;
        RECT 50.440 36.470 50.760 36.790 ;
        RECT 50.840 36.470 51.160 36.790 ;
        RECT 51.240 36.470 51.560 36.790 ;
        RECT 51.640 36.470 51.960 36.790 ;
        RECT 95.880 36.470 96.200 36.790 ;
        RECT 96.280 36.470 96.600 36.790 ;
        RECT 96.680 36.470 97.000 36.790 ;
        RECT 97.080 36.470 97.400 36.790 ;
        RECT 50.440 28.330 50.760 28.650 ;
        RECT 50.840 28.330 51.160 28.650 ;
        RECT 51.240 28.330 51.560 28.650 ;
        RECT 51.640 28.330 51.960 28.650 ;
        RECT 95.880 28.330 96.200 28.650 ;
        RECT 96.280 28.330 96.600 28.650 ;
        RECT 96.680 28.330 97.000 28.650 ;
        RECT 97.080 28.330 97.400 28.650 ;
        RECT 50.440 20.190 50.760 20.510 ;
        RECT 50.840 20.190 51.160 20.510 ;
        RECT 51.240 20.190 51.560 20.510 ;
        RECT 51.640 20.190 51.960 20.510 ;
        RECT 95.880 20.190 96.200 20.510 ;
        RECT 96.280 20.190 96.600 20.510 ;
        RECT 96.680 20.190 97.000 20.510 ;
        RECT 97.080 20.190 97.400 20.510 ;
      LAYER met4 ;
        RECT 50.400 16.020 52.000 150.850 ;
        RECT 95.840 16.020 97.440 150.850 ;
      LAYER M4M5_PR_C ;
        RECT 50.610 104.970 51.790 106.150 ;
        RECT 50.610 60.200 51.790 61.380 ;
        RECT 96.050 104.970 97.230 106.150 ;
        RECT 96.050 60.200 97.230 61.380 ;
      LAYER met5 ;
        RECT 5.760 104.760 142.080 106.370 ;
        RECT 5.760 59.990 142.080 61.600 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.760 150.500 5.920 150.680 ;
        RECT 6.090 150.500 6.400 150.680 ;
        RECT 6.570 150.500 6.880 150.680 ;
        RECT 7.050 150.500 7.360 150.680 ;
        RECT 7.530 150.500 7.840 150.680 ;
        RECT 8.010 150.500 8.320 150.680 ;
        RECT 8.490 150.500 8.800 150.680 ;
        RECT 8.970 150.500 9.280 150.680 ;
        RECT 9.450 150.500 9.760 150.680 ;
        RECT 9.930 150.500 10.240 150.680 ;
        RECT 10.410 150.500 10.720 150.680 ;
        RECT 10.890 150.500 11.200 150.680 ;
        RECT 11.370 150.500 11.680 150.680 ;
        RECT 11.850 150.500 12.160 150.680 ;
        RECT 12.330 150.500 12.640 150.680 ;
        RECT 12.810 150.500 13.120 150.680 ;
        RECT 13.290 150.500 13.600 150.680 ;
        RECT 13.770 150.500 14.080 150.680 ;
        RECT 14.250 150.500 14.560 150.680 ;
        RECT 14.730 150.500 15.040 150.680 ;
        RECT 15.210 150.500 15.520 150.680 ;
        RECT 15.690 150.500 16.000 150.680 ;
        RECT 16.170 150.500 16.480 150.680 ;
        RECT 16.650 150.500 16.960 150.680 ;
        RECT 17.130 150.500 17.440 150.680 ;
        RECT 17.610 150.500 17.920 150.680 ;
        RECT 18.090 150.500 18.400 150.680 ;
        RECT 18.570 150.500 18.880 150.680 ;
        RECT 19.050 150.500 19.360 150.680 ;
        RECT 19.530 150.500 19.840 150.680 ;
        RECT 20.010 150.500 20.320 150.680 ;
        RECT 20.490 150.500 20.800 150.680 ;
        RECT 20.970 150.500 21.280 150.680 ;
        RECT 21.450 150.500 21.760 150.680 ;
        RECT 21.930 150.500 22.240 150.680 ;
        RECT 22.410 150.500 22.720 150.680 ;
        RECT 22.890 150.500 23.200 150.680 ;
        RECT 23.370 150.500 23.680 150.680 ;
        RECT 23.850 150.500 24.160 150.680 ;
        RECT 24.330 150.500 24.640 150.680 ;
        RECT 24.810 150.500 25.120 150.680 ;
        RECT 25.290 150.500 25.600 150.680 ;
        RECT 25.770 150.500 26.080 150.680 ;
        RECT 26.250 150.500 26.560 150.680 ;
        RECT 26.730 150.500 27.040 150.680 ;
        RECT 27.210 150.500 27.520 150.680 ;
        RECT 27.690 150.500 28.000 150.680 ;
        RECT 28.170 150.500 28.480 150.680 ;
        RECT 28.650 150.500 28.960 150.680 ;
        RECT 29.130 150.500 29.440 150.680 ;
        RECT 29.610 150.500 29.920 150.680 ;
        RECT 30.090 150.500 30.400 150.680 ;
        RECT 30.570 150.500 30.880 150.680 ;
        RECT 31.050 150.500 31.360 150.680 ;
        RECT 31.530 150.500 31.840 150.680 ;
        RECT 32.010 150.500 32.320 150.680 ;
        RECT 32.490 150.500 32.800 150.680 ;
        RECT 32.970 150.500 33.280 150.680 ;
        RECT 33.450 150.500 33.760 150.680 ;
        RECT 33.930 150.500 34.240 150.680 ;
        RECT 34.410 150.500 34.720 150.680 ;
        RECT 34.890 150.500 35.200 150.680 ;
        RECT 35.370 150.500 35.680 150.680 ;
        RECT 35.850 150.500 36.160 150.680 ;
        RECT 36.330 150.500 36.640 150.680 ;
        RECT 36.810 150.500 37.120 150.680 ;
        RECT 37.290 150.500 37.600 150.680 ;
        RECT 37.770 150.500 38.080 150.680 ;
        RECT 38.250 150.500 38.560 150.680 ;
        RECT 38.730 150.500 39.040 150.680 ;
        RECT 39.210 150.500 39.520 150.680 ;
        RECT 39.690 150.500 40.000 150.680 ;
        RECT 40.170 150.500 40.480 150.680 ;
        RECT 40.650 150.500 40.960 150.680 ;
        RECT 41.130 150.500 41.440 150.680 ;
        RECT 41.610 150.500 41.920 150.680 ;
        RECT 42.090 150.500 42.400 150.680 ;
        RECT 42.570 150.500 42.880 150.680 ;
        RECT 43.050 150.500 43.360 150.680 ;
        RECT 43.530 150.500 43.840 150.680 ;
        RECT 44.010 150.500 44.320 150.680 ;
        RECT 44.490 150.500 44.800 150.680 ;
        RECT 44.970 150.500 45.280 150.680 ;
        RECT 45.450 150.500 45.760 150.680 ;
        RECT 45.930 150.500 46.240 150.680 ;
        RECT 46.410 150.500 46.720 150.680 ;
        RECT 46.890 150.500 47.200 150.680 ;
        RECT 47.370 150.500 47.680 150.680 ;
        RECT 47.850 150.500 48.160 150.680 ;
        RECT 48.330 150.500 48.640 150.680 ;
        RECT 48.810 150.500 49.120 150.680 ;
        RECT 49.290 150.500 49.600 150.680 ;
        RECT 49.770 150.500 50.080 150.680 ;
        RECT 50.250 150.500 50.560 150.680 ;
        RECT 50.730 150.500 51.040 150.680 ;
        RECT 51.210 150.500 51.520 150.680 ;
        RECT 51.690 150.500 52.000 150.680 ;
        RECT 52.170 150.500 52.480 150.680 ;
        RECT 52.650 150.500 52.960 150.680 ;
        RECT 53.130 150.500 53.440 150.680 ;
        RECT 53.610 150.500 53.920 150.680 ;
        RECT 54.090 150.500 54.400 150.680 ;
        RECT 54.570 150.500 54.880 150.680 ;
        RECT 55.050 150.500 55.360 150.680 ;
        RECT 55.530 150.500 55.840 150.680 ;
        RECT 56.010 150.500 56.320 150.680 ;
        RECT 56.490 150.500 56.800 150.680 ;
        RECT 56.970 150.500 57.280 150.680 ;
        RECT 57.450 150.500 57.760 150.680 ;
        RECT 57.930 150.500 58.240 150.680 ;
        RECT 58.410 150.500 58.720 150.680 ;
        RECT 58.890 150.500 59.200 150.680 ;
        RECT 59.370 150.500 59.680 150.680 ;
        RECT 59.850 150.500 60.160 150.680 ;
        RECT 60.330 150.500 60.640 150.680 ;
        RECT 60.810 150.500 61.120 150.680 ;
        RECT 61.290 150.500 61.600 150.680 ;
        RECT 61.770 150.500 62.080 150.680 ;
        RECT 62.250 150.500 62.560 150.680 ;
        RECT 62.730 150.500 63.040 150.680 ;
        RECT 63.210 150.500 63.520 150.680 ;
        RECT 63.690 150.500 64.000 150.680 ;
        RECT 64.170 150.500 64.480 150.680 ;
        RECT 64.650 150.500 64.960 150.680 ;
        RECT 65.130 150.500 65.440 150.680 ;
        RECT 65.610 150.500 65.920 150.680 ;
        RECT 66.090 150.500 66.400 150.680 ;
        RECT 66.570 150.500 66.880 150.680 ;
        RECT 67.050 150.500 67.360 150.680 ;
        RECT 67.530 150.500 67.840 150.680 ;
        RECT 68.010 150.500 68.320 150.680 ;
        RECT 68.490 150.500 68.800 150.680 ;
        RECT 68.970 150.500 69.280 150.680 ;
        RECT 69.450 150.500 69.760 150.680 ;
        RECT 69.930 150.500 70.240 150.680 ;
        RECT 70.410 150.500 70.720 150.680 ;
        RECT 70.890 150.500 71.200 150.680 ;
        RECT 71.370 150.500 71.680 150.680 ;
        RECT 71.850 150.500 72.160 150.680 ;
        RECT 72.330 150.500 72.640 150.680 ;
        RECT 72.810 150.500 73.120 150.680 ;
        RECT 73.290 150.500 73.600 150.680 ;
        RECT 73.770 150.500 74.080 150.680 ;
        RECT 74.250 150.500 74.560 150.680 ;
        RECT 74.730 150.500 75.040 150.680 ;
        RECT 75.210 150.500 75.520 150.680 ;
        RECT 75.690 150.500 76.000 150.680 ;
        RECT 76.170 150.500 76.480 150.680 ;
        RECT 76.650 150.500 76.960 150.680 ;
        RECT 77.130 150.500 77.440 150.680 ;
        RECT 77.610 150.500 77.920 150.680 ;
        RECT 78.090 150.500 78.400 150.680 ;
        RECT 78.570 150.500 78.880 150.680 ;
        RECT 79.050 150.500 79.360 150.680 ;
        RECT 79.530 150.500 79.840 150.680 ;
        RECT 80.010 150.500 80.320 150.680 ;
        RECT 80.490 150.500 80.800 150.680 ;
        RECT 80.970 150.500 81.280 150.680 ;
        RECT 81.450 150.500 81.760 150.680 ;
        RECT 81.930 150.500 82.240 150.680 ;
        RECT 82.410 150.500 82.720 150.680 ;
        RECT 82.890 150.500 83.200 150.680 ;
        RECT 83.370 150.500 83.680 150.680 ;
        RECT 83.850 150.500 84.160 150.680 ;
        RECT 84.330 150.500 84.640 150.680 ;
        RECT 84.810 150.500 85.120 150.680 ;
        RECT 85.290 150.500 85.600 150.680 ;
        RECT 85.770 150.500 86.080 150.680 ;
        RECT 86.250 150.500 86.560 150.680 ;
        RECT 86.730 150.500 87.040 150.680 ;
        RECT 87.210 150.500 87.520 150.680 ;
        RECT 87.690 150.500 88.000 150.680 ;
        RECT 88.170 150.500 88.480 150.680 ;
        RECT 88.650 150.500 88.960 150.680 ;
        RECT 89.130 150.500 89.440 150.680 ;
        RECT 89.610 150.500 89.920 150.680 ;
        RECT 90.090 150.500 90.400 150.680 ;
        RECT 90.570 150.500 90.880 150.680 ;
        RECT 91.050 150.500 91.360 150.680 ;
        RECT 91.530 150.500 91.840 150.680 ;
        RECT 92.010 150.500 92.320 150.680 ;
        RECT 92.490 150.500 92.800 150.680 ;
        RECT 92.970 150.500 93.280 150.680 ;
        RECT 93.450 150.500 93.760 150.680 ;
        RECT 93.930 150.500 94.240 150.680 ;
        RECT 94.410 150.500 94.720 150.680 ;
        RECT 94.890 150.500 95.200 150.680 ;
        RECT 95.370 150.500 95.680 150.680 ;
        RECT 95.850 150.500 96.160 150.680 ;
        RECT 96.330 150.500 96.640 150.680 ;
        RECT 96.810 150.500 97.120 150.680 ;
        RECT 97.290 150.500 97.600 150.680 ;
        RECT 97.770 150.500 98.080 150.680 ;
        RECT 98.250 150.500 98.560 150.680 ;
        RECT 98.730 150.500 99.040 150.680 ;
        RECT 99.210 150.500 99.520 150.680 ;
        RECT 99.690 150.500 100.000 150.680 ;
        RECT 100.170 150.500 100.480 150.680 ;
        RECT 100.650 150.500 100.960 150.680 ;
        RECT 101.130 150.500 101.440 150.680 ;
        RECT 101.610 150.500 101.920 150.680 ;
        RECT 102.090 150.500 102.400 150.680 ;
        RECT 102.570 150.500 102.880 150.680 ;
        RECT 103.050 150.500 103.360 150.680 ;
        RECT 103.530 150.500 103.840 150.680 ;
        RECT 104.010 150.500 104.320 150.680 ;
        RECT 104.490 150.500 104.800 150.680 ;
        RECT 104.970 150.500 105.280 150.680 ;
        RECT 105.450 150.500 105.760 150.680 ;
        RECT 105.930 150.500 106.240 150.680 ;
        RECT 106.410 150.500 106.720 150.680 ;
        RECT 106.890 150.500 107.200 150.680 ;
        RECT 107.370 150.500 107.680 150.680 ;
        RECT 107.850 150.500 108.160 150.680 ;
        RECT 108.330 150.500 108.640 150.680 ;
        RECT 108.810 150.500 109.120 150.680 ;
        RECT 109.290 150.500 109.600 150.680 ;
        RECT 109.770 150.500 110.080 150.680 ;
        RECT 110.250 150.500 110.560 150.680 ;
        RECT 110.730 150.500 111.040 150.680 ;
        RECT 111.210 150.500 111.520 150.680 ;
        RECT 111.690 150.500 112.000 150.680 ;
        RECT 112.170 150.500 112.480 150.680 ;
        RECT 112.650 150.500 112.960 150.680 ;
        RECT 113.130 150.500 113.440 150.680 ;
        RECT 113.610 150.500 113.920 150.680 ;
        RECT 114.090 150.500 114.400 150.680 ;
        RECT 114.570 150.500 114.880 150.680 ;
        RECT 115.050 150.500 115.360 150.680 ;
        RECT 115.530 150.500 115.840 150.680 ;
        RECT 116.010 150.500 116.320 150.680 ;
        RECT 116.490 150.500 116.800 150.680 ;
        RECT 116.970 150.500 117.280 150.680 ;
        RECT 117.450 150.500 117.760 150.680 ;
        RECT 117.930 150.500 118.240 150.680 ;
        RECT 118.410 150.500 118.720 150.680 ;
        RECT 118.890 150.500 119.200 150.680 ;
        RECT 119.370 150.500 119.680 150.680 ;
        RECT 119.850 150.500 120.160 150.680 ;
        RECT 120.330 150.500 120.640 150.680 ;
        RECT 120.810 150.500 121.120 150.680 ;
        RECT 121.290 150.500 121.600 150.680 ;
        RECT 121.770 150.500 122.080 150.680 ;
        RECT 122.250 150.500 122.560 150.680 ;
        RECT 122.730 150.500 123.040 150.680 ;
        RECT 123.210 150.500 123.520 150.680 ;
        RECT 123.690 150.500 124.000 150.680 ;
        RECT 124.170 150.500 124.480 150.680 ;
        RECT 124.650 150.500 124.960 150.680 ;
        RECT 125.130 150.500 125.440 150.680 ;
        RECT 125.610 150.500 125.920 150.680 ;
        RECT 126.090 150.500 126.400 150.680 ;
        RECT 126.570 150.500 126.880 150.680 ;
        RECT 127.050 150.500 127.360 150.680 ;
        RECT 127.530 150.500 127.840 150.680 ;
        RECT 128.010 150.500 128.320 150.680 ;
        RECT 128.490 150.500 128.800 150.680 ;
        RECT 128.970 150.500 129.280 150.680 ;
        RECT 129.450 150.500 129.760 150.680 ;
        RECT 129.930 150.500 130.240 150.680 ;
        RECT 130.410 150.500 130.720 150.680 ;
        RECT 130.890 150.500 131.200 150.680 ;
        RECT 131.370 150.500 131.680 150.680 ;
        RECT 131.850 150.500 132.160 150.680 ;
        RECT 132.330 150.500 132.640 150.680 ;
        RECT 132.810 150.500 133.120 150.680 ;
        RECT 133.290 150.500 133.600 150.680 ;
        RECT 133.770 150.500 134.080 150.680 ;
        RECT 134.250 150.500 134.560 150.680 ;
        RECT 134.730 150.500 135.040 150.680 ;
        RECT 135.210 150.500 135.520 150.680 ;
        RECT 135.690 150.500 136.000 150.680 ;
        RECT 136.170 150.500 136.480 150.680 ;
        RECT 136.650 150.500 136.960 150.680 ;
        RECT 137.130 150.500 137.440 150.680 ;
        RECT 137.610 150.500 137.920 150.680 ;
        RECT 138.090 150.500 138.400 150.680 ;
        RECT 138.570 150.500 138.880 150.680 ;
        RECT 139.050 150.500 139.360 150.680 ;
        RECT 139.530 150.500 139.840 150.680 ;
        RECT 140.010 150.500 140.320 150.680 ;
        RECT 140.490 150.500 140.800 150.680 ;
        RECT 140.970 150.500 141.280 150.680 ;
        RECT 141.450 150.500 141.600 150.680 ;
        RECT 6.340 150.200 9.070 150.230 ;
        RECT 6.340 150.030 6.510 150.200 ;
        RECT 6.680 150.030 6.950 150.200 ;
        RECT 7.120 150.030 7.360 150.200 ;
        RECT 7.530 150.030 7.790 150.200 ;
        RECT 7.960 150.030 8.230 150.200 ;
        RECT 8.400 150.030 8.640 150.200 ;
        RECT 8.810 150.030 9.070 150.200 ;
        RECT 6.340 149.230 9.070 150.030 ;
        RECT 10.180 150.200 12.910 150.230 ;
        RECT 10.180 150.030 10.350 150.200 ;
        RECT 10.520 150.030 10.790 150.200 ;
        RECT 10.960 150.030 11.200 150.200 ;
        RECT 11.370 150.030 11.630 150.200 ;
        RECT 11.800 150.030 12.070 150.200 ;
        RECT 12.240 150.030 12.480 150.200 ;
        RECT 12.650 150.030 12.910 150.200 ;
        RECT 10.180 149.230 12.910 150.030 ;
        RECT 14.020 150.200 16.750 150.230 ;
        RECT 14.020 150.030 14.190 150.200 ;
        RECT 14.360 150.030 14.630 150.200 ;
        RECT 14.800 150.030 15.040 150.200 ;
        RECT 15.210 150.030 15.470 150.200 ;
        RECT 15.640 150.030 15.910 150.200 ;
        RECT 16.080 150.030 16.320 150.200 ;
        RECT 16.490 150.030 16.750 150.200 ;
        RECT 14.020 149.230 16.750 150.030 ;
        RECT 17.860 150.200 20.590 150.230 ;
        RECT 17.860 150.030 18.030 150.200 ;
        RECT 18.200 150.030 18.470 150.200 ;
        RECT 18.640 150.030 18.880 150.200 ;
        RECT 19.050 150.030 19.310 150.200 ;
        RECT 19.480 150.030 19.750 150.200 ;
        RECT 19.920 150.030 20.160 150.200 ;
        RECT 20.330 150.030 20.590 150.200 ;
        RECT 23.620 150.190 24.270 150.300 ;
        RECT 17.860 149.230 20.590 150.030 ;
      LAYER li1 ;
        RECT 22.370 149.520 22.950 150.160 ;
      LAYER li1 ;
        RECT 23.620 150.020 23.680 150.190 ;
        RECT 23.850 150.020 24.040 150.190 ;
        RECT 24.210 150.020 24.270 150.190 ;
        RECT 23.620 149.960 24.270 150.020 ;
        RECT 23.860 149.520 24.270 149.960 ;
        RECT 25.060 150.200 27.790 150.230 ;
        RECT 25.060 150.030 25.230 150.200 ;
        RECT 25.400 150.030 25.670 150.200 ;
        RECT 25.840 150.030 26.080 150.200 ;
        RECT 26.250 150.030 26.510 150.200 ;
        RECT 26.680 150.030 26.950 150.200 ;
        RECT 27.120 150.030 27.360 150.200 ;
        RECT 27.530 150.030 27.790 150.200 ;
        RECT 6.500 148.560 6.830 149.230 ;
        RECT 7.230 147.910 7.560 148.890 ;
        RECT 7.780 148.560 8.110 149.230 ;
        RECT 8.510 147.910 8.840 148.890 ;
        RECT 10.340 148.560 10.670 149.230 ;
        RECT 11.070 147.910 11.400 148.890 ;
        RECT 11.620 148.560 11.950 149.230 ;
        RECT 12.350 147.910 12.680 148.890 ;
        RECT 14.180 148.560 14.510 149.230 ;
        RECT 14.910 147.910 15.240 148.890 ;
        RECT 15.460 148.560 15.790 149.230 ;
        RECT 16.190 147.910 16.520 148.890 ;
        RECT 18.020 148.560 18.350 149.230 ;
        RECT 18.750 147.910 19.080 148.890 ;
        RECT 19.300 148.560 19.630 149.230 ;
        RECT 20.030 147.910 20.360 148.890 ;
      LAYER li1 ;
        RECT 22.700 148.650 22.950 149.520 ;
      LAYER li1 ;
        RECT 25.060 149.230 27.790 150.030 ;
        RECT 28.900 150.200 31.630 150.230 ;
        RECT 28.900 150.030 29.070 150.200 ;
        RECT 29.240 150.030 29.510 150.200 ;
        RECT 29.680 150.030 29.920 150.200 ;
        RECT 30.090 150.030 30.350 150.200 ;
        RECT 30.520 150.030 30.790 150.200 ;
        RECT 30.960 150.030 31.200 150.200 ;
        RECT 31.370 150.030 31.630 150.200 ;
        RECT 28.900 149.230 31.630 150.030 ;
        RECT 32.740 150.200 35.470 150.230 ;
        RECT 32.740 150.030 32.910 150.200 ;
        RECT 33.080 150.030 33.350 150.200 ;
        RECT 33.520 150.030 33.760 150.200 ;
        RECT 33.930 150.030 34.190 150.200 ;
        RECT 34.360 150.030 34.630 150.200 ;
        RECT 34.800 150.030 35.040 150.200 ;
        RECT 35.210 150.030 35.470 150.200 ;
        RECT 32.740 149.230 35.470 150.030 ;
        RECT 36.580 150.200 39.310 150.230 ;
        RECT 36.580 150.030 36.750 150.200 ;
        RECT 36.920 150.030 37.190 150.200 ;
        RECT 37.360 150.030 37.600 150.200 ;
        RECT 37.770 150.030 38.030 150.200 ;
        RECT 38.200 150.030 38.470 150.200 ;
        RECT 38.640 150.030 38.880 150.200 ;
        RECT 39.050 150.030 39.310 150.200 ;
        RECT 36.580 149.230 39.310 150.030 ;
        RECT 40.420 150.200 43.150 150.230 ;
        RECT 40.420 150.030 40.590 150.200 ;
        RECT 40.760 150.030 41.030 150.200 ;
        RECT 41.200 150.030 41.440 150.200 ;
        RECT 41.610 150.030 41.870 150.200 ;
        RECT 42.040 150.030 42.310 150.200 ;
        RECT 42.480 150.030 42.720 150.200 ;
        RECT 42.890 150.030 43.150 150.200 ;
        RECT 40.420 149.230 43.150 150.030 ;
        RECT 44.260 150.200 46.990 150.230 ;
        RECT 44.260 150.030 44.430 150.200 ;
        RECT 44.600 150.030 44.870 150.200 ;
        RECT 45.040 150.030 45.280 150.200 ;
        RECT 45.450 150.030 45.710 150.200 ;
        RECT 45.880 150.030 46.150 150.200 ;
        RECT 46.320 150.030 46.560 150.200 ;
        RECT 46.730 150.030 46.990 150.200 ;
        RECT 44.260 149.230 46.990 150.030 ;
        RECT 48.100 150.200 50.830 150.230 ;
        RECT 48.100 150.030 48.270 150.200 ;
        RECT 48.440 150.030 48.710 150.200 ;
        RECT 48.880 150.030 49.120 150.200 ;
        RECT 49.290 150.030 49.550 150.200 ;
        RECT 49.720 150.030 49.990 150.200 ;
        RECT 50.160 150.030 50.400 150.200 ;
        RECT 50.570 150.030 50.830 150.200 ;
        RECT 48.100 149.230 50.830 150.030 ;
        RECT 51.940 150.200 54.670 150.230 ;
        RECT 51.940 150.030 52.110 150.200 ;
        RECT 52.280 150.030 52.550 150.200 ;
        RECT 52.720 150.030 52.960 150.200 ;
        RECT 53.130 150.030 53.390 150.200 ;
        RECT 53.560 150.030 53.830 150.200 ;
        RECT 54.000 150.030 54.240 150.200 ;
        RECT 54.410 150.030 54.670 150.200 ;
        RECT 51.940 149.230 54.670 150.030 ;
        RECT 55.780 150.200 58.510 150.230 ;
        RECT 55.780 150.030 55.950 150.200 ;
        RECT 56.120 150.030 56.390 150.200 ;
        RECT 56.560 150.030 56.800 150.200 ;
        RECT 56.970 150.030 57.230 150.200 ;
        RECT 57.400 150.030 57.670 150.200 ;
        RECT 57.840 150.030 58.080 150.200 ;
        RECT 58.250 150.030 58.510 150.200 ;
        RECT 55.780 149.230 58.510 150.030 ;
        RECT 59.620 150.200 62.350 150.230 ;
        RECT 59.620 150.030 59.790 150.200 ;
        RECT 59.960 150.030 60.230 150.200 ;
        RECT 60.400 150.030 60.640 150.200 ;
        RECT 60.810 150.030 61.070 150.200 ;
        RECT 61.240 150.030 61.510 150.200 ;
        RECT 61.680 150.030 61.920 150.200 ;
        RECT 62.090 150.030 62.350 150.200 ;
        RECT 59.620 149.230 62.350 150.030 ;
        RECT 63.050 150.190 64.660 150.220 ;
        RECT 63.050 150.020 63.100 150.190 ;
        RECT 63.270 150.020 63.540 150.190 ;
        RECT 63.710 150.020 63.980 150.190 ;
        RECT 64.150 150.020 64.390 150.190 ;
        RECT 64.560 150.020 64.660 150.190 ;
        RECT 66.340 150.190 66.990 150.300 ;
        RECT 63.050 149.740 64.660 150.020 ;
        RECT 63.360 149.340 64.660 149.740 ;
      LAYER li1 ;
        RECT 22.700 148.400 23.410 148.650 ;
      LAYER li1 ;
        RECT 25.220 148.560 25.550 149.230 ;
        RECT 6.260 147.030 9.000 147.910 ;
        RECT 6.260 146.860 6.470 147.030 ;
        RECT 6.640 146.860 6.910 147.030 ;
        RECT 7.080 146.860 7.320 147.030 ;
        RECT 7.490 146.860 7.750 147.030 ;
        RECT 7.920 146.860 8.190 147.030 ;
        RECT 8.360 146.860 8.600 147.030 ;
        RECT 8.770 146.860 9.000 147.030 ;
        RECT 6.260 146.840 9.000 146.860 ;
        RECT 10.100 147.030 12.840 147.910 ;
        RECT 10.100 146.860 10.310 147.030 ;
        RECT 10.480 146.860 10.750 147.030 ;
        RECT 10.920 146.860 11.160 147.030 ;
        RECT 11.330 146.860 11.590 147.030 ;
        RECT 11.760 146.860 12.030 147.030 ;
        RECT 12.200 146.860 12.440 147.030 ;
        RECT 12.610 146.860 12.840 147.030 ;
        RECT 10.100 146.840 12.840 146.860 ;
        RECT 13.940 147.030 16.680 147.910 ;
        RECT 13.940 146.860 14.150 147.030 ;
        RECT 14.320 146.860 14.590 147.030 ;
        RECT 14.760 146.860 15.000 147.030 ;
        RECT 15.170 146.860 15.430 147.030 ;
        RECT 15.600 146.860 15.870 147.030 ;
        RECT 16.040 146.860 16.280 147.030 ;
        RECT 16.450 146.860 16.680 147.030 ;
        RECT 13.940 146.840 16.680 146.860 ;
        RECT 17.780 147.030 20.520 147.910 ;
        RECT 17.780 146.860 17.990 147.030 ;
        RECT 18.160 146.860 18.430 147.030 ;
        RECT 18.600 146.860 18.840 147.030 ;
        RECT 19.010 146.860 19.270 147.030 ;
        RECT 19.440 146.860 19.710 147.030 ;
        RECT 19.880 146.860 20.120 147.030 ;
        RECT 20.290 146.860 20.520 147.030 ;
        RECT 17.780 146.840 20.520 146.860 ;
        RECT 22.300 147.140 22.700 147.410 ;
        RECT 22.300 147.080 22.950 147.140 ;
        RECT 22.300 146.910 22.360 147.080 ;
        RECT 22.530 146.910 22.720 147.080 ;
        RECT 22.890 146.910 22.950 147.080 ;
      LAYER li1 ;
        RECT 23.160 147.060 23.410 148.400 ;
      LAYER li1 ;
        RECT 25.950 147.910 26.280 148.890 ;
        RECT 26.500 148.560 26.830 149.230 ;
        RECT 27.230 147.910 27.560 148.890 ;
        RECT 29.060 148.560 29.390 149.230 ;
        RECT 29.790 147.910 30.120 148.890 ;
        RECT 30.340 148.560 30.670 149.230 ;
        RECT 31.070 147.910 31.400 148.890 ;
        RECT 32.900 148.560 33.230 149.230 ;
        RECT 33.630 147.910 33.960 148.890 ;
        RECT 34.180 148.560 34.510 149.230 ;
        RECT 34.910 147.910 35.240 148.890 ;
        RECT 36.740 148.560 37.070 149.230 ;
        RECT 37.470 147.910 37.800 148.890 ;
        RECT 38.020 148.560 38.350 149.230 ;
        RECT 38.750 147.910 39.080 148.890 ;
        RECT 40.580 148.560 40.910 149.230 ;
        RECT 41.310 147.910 41.640 148.890 ;
        RECT 41.860 148.560 42.190 149.230 ;
        RECT 42.590 147.910 42.920 148.890 ;
        RECT 44.420 148.560 44.750 149.230 ;
        RECT 45.150 147.910 45.480 148.890 ;
        RECT 45.700 148.560 46.030 149.230 ;
        RECT 46.430 147.910 46.760 148.890 ;
        RECT 48.260 148.560 48.590 149.230 ;
        RECT 48.990 147.910 49.320 148.890 ;
        RECT 49.540 148.560 49.870 149.230 ;
        RECT 50.270 147.910 50.600 148.890 ;
        RECT 52.100 148.560 52.430 149.230 ;
        RECT 52.830 147.910 53.160 148.890 ;
        RECT 53.380 148.560 53.710 149.230 ;
        RECT 54.110 147.910 54.440 148.890 ;
        RECT 55.940 148.560 56.270 149.230 ;
        RECT 56.670 147.910 57.000 148.890 ;
        RECT 57.220 148.560 57.550 149.230 ;
        RECT 57.950 147.910 58.280 148.890 ;
        RECT 59.780 148.560 60.110 149.230 ;
        RECT 60.510 147.910 60.840 148.890 ;
        RECT 61.060 148.560 61.390 149.230 ;
        RECT 61.790 147.910 62.120 148.890 ;
        RECT 63.360 148.560 63.690 149.340 ;
      LAYER li1 ;
        RECT 65.840 149.090 66.170 150.090 ;
      LAYER li1 ;
        RECT 66.340 150.020 66.400 150.190 ;
        RECT 66.570 150.020 66.760 150.190 ;
        RECT 66.930 150.020 66.990 150.190 ;
        RECT 66.340 149.960 66.990 150.020 ;
        RECT 66.580 149.520 66.990 149.960 ;
        RECT 67.780 150.200 70.510 150.230 ;
        RECT 67.780 150.030 67.950 150.200 ;
        RECT 68.120 150.030 68.390 150.200 ;
        RECT 68.560 150.030 68.800 150.200 ;
        RECT 68.970 150.030 69.230 150.200 ;
        RECT 69.400 150.030 69.670 150.200 ;
        RECT 69.840 150.030 70.080 150.200 ;
        RECT 70.250 150.030 70.510 150.200 ;
        RECT 67.780 149.230 70.510 150.030 ;
        RECT 71.620 150.200 74.350 150.230 ;
        RECT 71.620 150.030 71.790 150.200 ;
        RECT 71.960 150.030 72.230 150.200 ;
        RECT 72.400 150.030 72.640 150.200 ;
        RECT 72.810 150.030 73.070 150.200 ;
        RECT 73.240 150.030 73.510 150.200 ;
        RECT 73.680 150.030 73.920 150.200 ;
        RECT 74.090 150.030 74.350 150.200 ;
        RECT 76.420 150.190 77.070 150.300 ;
        RECT 71.620 149.230 74.350 150.030 ;
        RECT 22.300 146.800 22.950 146.910 ;
        RECT 24.980 147.030 27.720 147.910 ;
        RECT 24.980 146.860 25.190 147.030 ;
        RECT 25.360 146.860 25.630 147.030 ;
        RECT 25.800 146.860 26.040 147.030 ;
        RECT 26.210 146.860 26.470 147.030 ;
        RECT 26.640 146.860 26.910 147.030 ;
        RECT 27.080 146.860 27.320 147.030 ;
        RECT 27.490 146.860 27.720 147.030 ;
        RECT 24.980 146.840 27.720 146.860 ;
        RECT 28.820 147.030 31.560 147.910 ;
        RECT 28.820 146.860 29.030 147.030 ;
        RECT 29.200 146.860 29.470 147.030 ;
        RECT 29.640 146.860 29.880 147.030 ;
        RECT 30.050 146.860 30.310 147.030 ;
        RECT 30.480 146.860 30.750 147.030 ;
        RECT 30.920 146.860 31.160 147.030 ;
        RECT 31.330 146.860 31.560 147.030 ;
        RECT 28.820 146.840 31.560 146.860 ;
        RECT 32.660 147.030 35.400 147.910 ;
        RECT 32.660 146.860 32.870 147.030 ;
        RECT 33.040 146.860 33.310 147.030 ;
        RECT 33.480 146.860 33.720 147.030 ;
        RECT 33.890 146.860 34.150 147.030 ;
        RECT 34.320 146.860 34.590 147.030 ;
        RECT 34.760 146.860 35.000 147.030 ;
        RECT 35.170 146.860 35.400 147.030 ;
        RECT 32.660 146.840 35.400 146.860 ;
        RECT 36.500 147.030 39.240 147.910 ;
        RECT 36.500 146.860 36.710 147.030 ;
        RECT 36.880 146.860 37.150 147.030 ;
        RECT 37.320 146.860 37.560 147.030 ;
        RECT 37.730 146.860 37.990 147.030 ;
        RECT 38.160 146.860 38.430 147.030 ;
        RECT 38.600 146.860 38.840 147.030 ;
        RECT 39.010 146.860 39.240 147.030 ;
        RECT 36.500 146.840 39.240 146.860 ;
        RECT 40.340 147.030 43.080 147.910 ;
        RECT 40.340 146.860 40.550 147.030 ;
        RECT 40.720 146.860 40.990 147.030 ;
        RECT 41.160 146.860 41.400 147.030 ;
        RECT 41.570 146.860 41.830 147.030 ;
        RECT 42.000 146.860 42.270 147.030 ;
        RECT 42.440 146.860 42.680 147.030 ;
        RECT 42.850 146.860 43.080 147.030 ;
        RECT 40.340 146.840 43.080 146.860 ;
        RECT 44.180 147.030 46.920 147.910 ;
        RECT 44.180 146.860 44.390 147.030 ;
        RECT 44.560 146.860 44.830 147.030 ;
        RECT 45.000 146.860 45.240 147.030 ;
        RECT 45.410 146.860 45.670 147.030 ;
        RECT 45.840 146.860 46.110 147.030 ;
        RECT 46.280 146.860 46.520 147.030 ;
        RECT 46.690 146.860 46.920 147.030 ;
        RECT 44.180 146.840 46.920 146.860 ;
        RECT 48.020 147.030 50.760 147.910 ;
        RECT 48.020 146.860 48.230 147.030 ;
        RECT 48.400 146.860 48.670 147.030 ;
        RECT 48.840 146.860 49.080 147.030 ;
        RECT 49.250 146.860 49.510 147.030 ;
        RECT 49.680 146.860 49.950 147.030 ;
        RECT 50.120 146.860 50.360 147.030 ;
        RECT 50.530 146.860 50.760 147.030 ;
        RECT 48.020 146.840 50.760 146.860 ;
        RECT 51.860 147.030 54.600 147.910 ;
        RECT 51.860 146.860 52.070 147.030 ;
        RECT 52.240 146.860 52.510 147.030 ;
        RECT 52.680 146.860 52.920 147.030 ;
        RECT 53.090 146.860 53.350 147.030 ;
        RECT 53.520 146.860 53.790 147.030 ;
        RECT 53.960 146.860 54.200 147.030 ;
        RECT 54.370 146.860 54.600 147.030 ;
        RECT 51.860 146.840 54.600 146.860 ;
        RECT 55.700 147.030 58.440 147.910 ;
        RECT 55.700 146.860 55.910 147.030 ;
        RECT 56.080 146.860 56.350 147.030 ;
        RECT 56.520 146.860 56.760 147.030 ;
        RECT 56.930 146.860 57.190 147.030 ;
        RECT 57.360 146.860 57.630 147.030 ;
        RECT 57.800 146.860 58.040 147.030 ;
        RECT 58.210 146.860 58.440 147.030 ;
        RECT 55.700 146.840 58.440 146.860 ;
        RECT 59.540 147.030 62.280 147.910 ;
        RECT 63.900 147.900 64.230 148.890 ;
      LAYER li1 ;
        RECT 65.840 148.820 66.600 149.090 ;
      LAYER li1 ;
        RECT 59.540 146.860 59.750 147.030 ;
        RECT 59.920 146.860 60.190 147.030 ;
        RECT 60.360 146.860 60.600 147.030 ;
        RECT 60.770 146.860 61.030 147.030 ;
        RECT 61.200 146.860 61.470 147.030 ;
        RECT 61.640 146.860 61.880 147.030 ;
        RECT 62.050 146.860 62.280 147.030 ;
        RECT 59.540 146.840 62.280 146.860 ;
        RECT 63.130 147.030 64.580 147.900 ;
      LAYER li1 ;
        RECT 66.330 147.410 66.600 148.820 ;
      LAYER li1 ;
        RECT 67.940 148.560 68.270 149.230 ;
        RECT 68.670 147.910 69.000 148.890 ;
        RECT 69.220 148.560 69.550 149.230 ;
        RECT 69.950 147.910 70.280 148.890 ;
        RECT 71.780 148.560 72.110 149.230 ;
        RECT 72.510 147.910 72.840 148.890 ;
        RECT 73.060 148.560 73.390 149.230 ;
      LAYER li1 ;
        RECT 75.920 149.090 76.250 150.090 ;
      LAYER li1 ;
        RECT 76.420 150.020 76.480 150.190 ;
        RECT 76.650 150.020 76.840 150.190 ;
        RECT 77.010 150.020 77.070 150.190 ;
        RECT 76.420 149.960 77.070 150.020 ;
        RECT 76.660 149.520 77.070 149.960 ;
        RECT 77.860 150.200 80.590 150.230 ;
        RECT 77.860 150.030 78.030 150.200 ;
        RECT 78.200 150.030 78.470 150.200 ;
        RECT 78.640 150.030 78.880 150.200 ;
        RECT 79.050 150.030 79.310 150.200 ;
        RECT 79.480 150.030 79.750 150.200 ;
        RECT 79.920 150.030 80.160 150.200 ;
        RECT 80.330 150.030 80.590 150.200 ;
        RECT 77.860 149.230 80.590 150.030 ;
        RECT 81.700 150.200 84.430 150.230 ;
        RECT 81.700 150.030 81.870 150.200 ;
        RECT 82.040 150.030 82.310 150.200 ;
        RECT 82.480 150.030 82.720 150.200 ;
        RECT 82.890 150.030 83.150 150.200 ;
        RECT 83.320 150.030 83.590 150.200 ;
        RECT 83.760 150.030 84.000 150.200 ;
        RECT 84.170 150.030 84.430 150.200 ;
        RECT 81.700 149.230 84.430 150.030 ;
        RECT 85.540 150.200 88.270 150.230 ;
        RECT 85.540 150.030 85.710 150.200 ;
        RECT 85.880 150.030 86.150 150.200 ;
        RECT 86.320 150.030 86.560 150.200 ;
        RECT 86.730 150.030 86.990 150.200 ;
        RECT 87.160 150.030 87.430 150.200 ;
        RECT 87.600 150.030 87.840 150.200 ;
        RECT 88.010 150.030 88.270 150.200 ;
        RECT 85.540 149.230 88.270 150.030 ;
        RECT 89.380 150.200 92.110 150.230 ;
        RECT 89.380 150.030 89.550 150.200 ;
        RECT 89.720 150.030 89.990 150.200 ;
        RECT 90.160 150.030 90.400 150.200 ;
        RECT 90.570 150.030 90.830 150.200 ;
        RECT 91.000 150.030 91.270 150.200 ;
        RECT 91.440 150.030 91.680 150.200 ;
        RECT 91.850 150.030 92.110 150.200 ;
        RECT 89.380 149.230 92.110 150.030 ;
        RECT 93.220 150.200 95.950 150.230 ;
        RECT 93.220 150.030 93.390 150.200 ;
        RECT 93.560 150.030 93.830 150.200 ;
        RECT 94.000 150.030 94.240 150.200 ;
        RECT 94.410 150.030 94.670 150.200 ;
        RECT 94.840 150.030 95.110 150.200 ;
        RECT 95.280 150.030 95.520 150.200 ;
        RECT 95.690 150.030 95.950 150.200 ;
        RECT 93.220 149.230 95.950 150.030 ;
        RECT 97.060 150.200 99.790 150.230 ;
        RECT 97.060 150.030 97.230 150.200 ;
        RECT 97.400 150.030 97.670 150.200 ;
        RECT 97.840 150.030 98.080 150.200 ;
        RECT 98.250 150.030 98.510 150.200 ;
        RECT 98.680 150.030 98.950 150.200 ;
        RECT 99.120 150.030 99.360 150.200 ;
        RECT 99.530 150.030 99.790 150.200 ;
        RECT 97.060 149.230 99.790 150.030 ;
        RECT 100.900 150.200 103.630 150.230 ;
        RECT 100.900 150.030 101.070 150.200 ;
        RECT 101.240 150.030 101.510 150.200 ;
        RECT 101.680 150.030 101.920 150.200 ;
        RECT 102.090 150.030 102.350 150.200 ;
        RECT 102.520 150.030 102.790 150.200 ;
        RECT 102.960 150.030 103.200 150.200 ;
        RECT 103.370 150.030 103.630 150.200 ;
        RECT 100.900 149.230 103.630 150.030 ;
        RECT 104.740 150.200 107.470 150.230 ;
        RECT 104.740 150.030 104.910 150.200 ;
        RECT 105.080 150.030 105.350 150.200 ;
        RECT 105.520 150.030 105.760 150.200 ;
        RECT 105.930 150.030 106.190 150.200 ;
        RECT 106.360 150.030 106.630 150.200 ;
        RECT 106.800 150.030 107.040 150.200 ;
        RECT 107.210 150.030 107.470 150.200 ;
        RECT 104.740 149.230 107.470 150.030 ;
        RECT 108.580 150.200 111.310 150.230 ;
        RECT 108.580 150.030 108.750 150.200 ;
        RECT 108.920 150.030 109.190 150.200 ;
        RECT 109.360 150.030 109.600 150.200 ;
        RECT 109.770 150.030 110.030 150.200 ;
        RECT 110.200 150.030 110.470 150.200 ;
        RECT 110.640 150.030 110.880 150.200 ;
        RECT 111.050 150.030 111.310 150.200 ;
        RECT 108.580 149.230 111.310 150.030 ;
        RECT 112.420 150.200 115.150 150.230 ;
        RECT 112.420 150.030 112.590 150.200 ;
        RECT 112.760 150.030 113.030 150.200 ;
        RECT 113.200 150.030 113.440 150.200 ;
        RECT 113.610 150.030 113.870 150.200 ;
        RECT 114.040 150.030 114.310 150.200 ;
        RECT 114.480 150.030 114.720 150.200 ;
        RECT 114.890 150.030 115.150 150.200 ;
        RECT 112.420 149.230 115.150 150.030 ;
        RECT 116.260 150.200 118.990 150.230 ;
        RECT 116.260 150.030 116.430 150.200 ;
        RECT 116.600 150.030 116.870 150.200 ;
        RECT 117.040 150.030 117.280 150.200 ;
        RECT 117.450 150.030 117.710 150.200 ;
        RECT 117.880 150.030 118.150 150.200 ;
        RECT 118.320 150.030 118.560 150.200 ;
        RECT 118.730 150.030 118.990 150.200 ;
        RECT 116.260 149.230 118.990 150.030 ;
        RECT 120.100 150.200 122.830 150.230 ;
        RECT 120.100 150.030 120.270 150.200 ;
        RECT 120.440 150.030 120.710 150.200 ;
        RECT 120.880 150.030 121.120 150.200 ;
        RECT 121.290 150.030 121.550 150.200 ;
        RECT 121.720 150.030 121.990 150.200 ;
        RECT 122.160 150.030 122.400 150.200 ;
        RECT 122.570 150.030 122.830 150.200 ;
        RECT 120.100 149.230 122.830 150.030 ;
        RECT 123.940 150.200 126.670 150.230 ;
        RECT 123.940 150.030 124.110 150.200 ;
        RECT 124.280 150.030 124.550 150.200 ;
        RECT 124.720 150.030 124.960 150.200 ;
        RECT 125.130 150.030 125.390 150.200 ;
        RECT 125.560 150.030 125.830 150.200 ;
        RECT 126.000 150.030 126.240 150.200 ;
        RECT 126.410 150.030 126.670 150.200 ;
        RECT 123.940 149.230 126.670 150.030 ;
        RECT 127.780 150.200 130.510 150.230 ;
        RECT 127.780 150.030 127.950 150.200 ;
        RECT 128.120 150.030 128.390 150.200 ;
        RECT 128.560 150.030 128.800 150.200 ;
        RECT 128.970 150.030 129.230 150.200 ;
        RECT 129.400 150.030 129.670 150.200 ;
        RECT 129.840 150.030 130.080 150.200 ;
        RECT 130.250 150.030 130.510 150.200 ;
        RECT 127.780 149.230 130.510 150.030 ;
        RECT 131.620 150.200 134.350 150.230 ;
        RECT 131.620 150.030 131.790 150.200 ;
        RECT 131.960 150.030 132.230 150.200 ;
        RECT 132.400 150.030 132.640 150.200 ;
        RECT 132.810 150.030 133.070 150.200 ;
        RECT 133.240 150.030 133.510 150.200 ;
        RECT 133.680 150.030 133.920 150.200 ;
        RECT 134.090 150.030 134.350 150.200 ;
        RECT 131.620 149.230 134.350 150.030 ;
        RECT 135.460 150.200 138.190 150.230 ;
        RECT 135.460 150.030 135.630 150.200 ;
        RECT 135.800 150.030 136.070 150.200 ;
        RECT 136.240 150.030 136.480 150.200 ;
        RECT 136.650 150.030 136.910 150.200 ;
        RECT 137.080 150.030 137.350 150.200 ;
        RECT 137.520 150.030 137.760 150.200 ;
        RECT 137.930 150.030 138.190 150.200 ;
        RECT 135.460 149.230 138.190 150.030 ;
        RECT 138.890 150.190 140.500 150.220 ;
        RECT 138.890 150.020 138.940 150.190 ;
        RECT 139.110 150.020 139.380 150.190 ;
        RECT 139.550 150.020 139.820 150.190 ;
        RECT 139.990 150.020 140.230 150.190 ;
        RECT 140.400 150.020 140.500 150.190 ;
        RECT 138.890 149.740 140.500 150.020 ;
        RECT 139.200 149.340 140.500 149.740 ;
        RECT 73.790 147.910 74.120 148.890 ;
      LAYER li1 ;
        RECT 75.920 148.820 76.680 149.090 ;
      LAYER li1 ;
        RECT 63.130 146.860 63.380 147.030 ;
        RECT 63.550 146.860 63.740 147.030 ;
        RECT 63.910 146.860 64.180 147.030 ;
        RECT 64.350 146.860 64.580 147.030 ;
        RECT 63.130 146.830 64.580 146.860 ;
        RECT 65.020 147.140 65.420 147.410 ;
        RECT 65.020 147.080 65.670 147.140 ;
        RECT 65.020 146.910 65.080 147.080 ;
        RECT 65.250 146.910 65.440 147.080 ;
        RECT 65.610 146.910 65.670 147.080 ;
        RECT 65.020 146.800 65.670 146.910 ;
      LAYER li1 ;
        RECT 66.330 146.770 66.910 147.410 ;
      LAYER li1 ;
        RECT 67.700 147.030 70.440 147.910 ;
        RECT 67.700 146.860 67.910 147.030 ;
        RECT 68.080 146.860 68.350 147.030 ;
        RECT 68.520 146.860 68.760 147.030 ;
        RECT 68.930 146.860 69.190 147.030 ;
        RECT 69.360 146.860 69.630 147.030 ;
        RECT 69.800 146.860 70.040 147.030 ;
        RECT 70.210 146.860 70.440 147.030 ;
        RECT 67.700 146.840 70.440 146.860 ;
        RECT 71.540 147.030 74.280 147.910 ;
      LAYER li1 ;
        RECT 76.410 147.410 76.680 148.820 ;
      LAYER li1 ;
        RECT 78.020 148.560 78.350 149.230 ;
        RECT 78.750 147.910 79.080 148.890 ;
        RECT 79.300 148.560 79.630 149.230 ;
        RECT 80.030 147.910 80.360 148.890 ;
        RECT 81.860 148.560 82.190 149.230 ;
        RECT 82.590 147.910 82.920 148.890 ;
        RECT 83.140 148.560 83.470 149.230 ;
        RECT 83.870 147.910 84.200 148.890 ;
        RECT 85.700 148.560 86.030 149.230 ;
        RECT 86.430 147.910 86.760 148.890 ;
        RECT 86.980 148.560 87.310 149.230 ;
        RECT 87.710 147.910 88.040 148.890 ;
        RECT 89.540 148.560 89.870 149.230 ;
        RECT 90.270 147.910 90.600 148.890 ;
        RECT 90.820 148.560 91.150 149.230 ;
        RECT 91.550 147.910 91.880 148.890 ;
        RECT 93.380 148.560 93.710 149.230 ;
        RECT 94.110 147.910 94.440 148.890 ;
        RECT 94.660 148.560 94.990 149.230 ;
        RECT 95.390 147.910 95.720 148.890 ;
        RECT 97.220 148.560 97.550 149.230 ;
        RECT 97.950 147.910 98.280 148.890 ;
        RECT 98.500 148.560 98.830 149.230 ;
        RECT 99.230 147.910 99.560 148.890 ;
        RECT 101.060 148.560 101.390 149.230 ;
        RECT 101.790 147.910 102.120 148.890 ;
        RECT 102.340 148.560 102.670 149.230 ;
        RECT 103.070 147.910 103.400 148.890 ;
        RECT 104.900 148.560 105.230 149.230 ;
        RECT 105.630 147.910 105.960 148.890 ;
        RECT 106.180 148.560 106.510 149.230 ;
        RECT 106.910 147.910 107.240 148.890 ;
        RECT 108.740 148.560 109.070 149.230 ;
        RECT 109.470 147.910 109.800 148.890 ;
        RECT 110.020 148.560 110.350 149.230 ;
        RECT 110.750 147.910 111.080 148.890 ;
        RECT 112.580 148.560 112.910 149.230 ;
        RECT 113.310 147.910 113.640 148.890 ;
        RECT 113.860 148.560 114.190 149.230 ;
        RECT 114.590 147.910 114.920 148.890 ;
        RECT 116.420 148.560 116.750 149.230 ;
        RECT 117.150 147.910 117.480 148.890 ;
        RECT 117.700 148.560 118.030 149.230 ;
        RECT 118.430 147.910 118.760 148.890 ;
        RECT 120.260 148.560 120.590 149.230 ;
        RECT 120.990 147.910 121.320 148.890 ;
        RECT 121.540 148.560 121.870 149.230 ;
        RECT 122.270 147.910 122.600 148.890 ;
        RECT 124.100 148.560 124.430 149.230 ;
        RECT 124.830 147.910 125.160 148.890 ;
        RECT 125.380 148.560 125.710 149.230 ;
        RECT 126.110 147.910 126.440 148.890 ;
        RECT 127.940 148.560 128.270 149.230 ;
        RECT 128.670 147.910 129.000 148.890 ;
        RECT 129.220 148.560 129.550 149.230 ;
        RECT 129.950 147.910 130.280 148.890 ;
        RECT 131.780 148.560 132.110 149.230 ;
        RECT 132.510 147.910 132.840 148.890 ;
        RECT 133.060 148.560 133.390 149.230 ;
        RECT 133.790 147.910 134.120 148.890 ;
        RECT 135.620 148.560 135.950 149.230 ;
        RECT 136.350 147.910 136.680 148.890 ;
        RECT 136.900 148.560 137.230 149.230 ;
        RECT 137.630 147.910 137.960 148.890 ;
        RECT 139.200 148.560 139.530 149.340 ;
        RECT 71.540 146.860 71.750 147.030 ;
        RECT 71.920 146.860 72.190 147.030 ;
        RECT 72.360 146.860 72.600 147.030 ;
        RECT 72.770 146.860 73.030 147.030 ;
        RECT 73.200 146.860 73.470 147.030 ;
        RECT 73.640 146.860 73.880 147.030 ;
        RECT 74.050 146.860 74.280 147.030 ;
        RECT 71.540 146.840 74.280 146.860 ;
        RECT 75.100 147.140 75.500 147.410 ;
        RECT 75.100 147.080 75.750 147.140 ;
        RECT 75.100 146.910 75.160 147.080 ;
        RECT 75.330 146.910 75.520 147.080 ;
        RECT 75.690 146.910 75.750 147.080 ;
        RECT 75.100 146.800 75.750 146.910 ;
      LAYER li1 ;
        RECT 76.410 146.770 76.990 147.410 ;
      LAYER li1 ;
        RECT 77.780 147.030 80.520 147.910 ;
        RECT 77.780 146.860 77.990 147.030 ;
        RECT 78.160 146.860 78.430 147.030 ;
        RECT 78.600 146.860 78.840 147.030 ;
        RECT 79.010 146.860 79.270 147.030 ;
        RECT 79.440 146.860 79.710 147.030 ;
        RECT 79.880 146.860 80.120 147.030 ;
        RECT 80.290 146.860 80.520 147.030 ;
        RECT 77.780 146.840 80.520 146.860 ;
        RECT 81.620 147.030 84.360 147.910 ;
        RECT 81.620 146.860 81.830 147.030 ;
        RECT 82.000 146.860 82.270 147.030 ;
        RECT 82.440 146.860 82.680 147.030 ;
        RECT 82.850 146.860 83.110 147.030 ;
        RECT 83.280 146.860 83.550 147.030 ;
        RECT 83.720 146.860 83.960 147.030 ;
        RECT 84.130 146.860 84.360 147.030 ;
        RECT 81.620 146.840 84.360 146.860 ;
        RECT 85.460 147.030 88.200 147.910 ;
        RECT 85.460 146.860 85.670 147.030 ;
        RECT 85.840 146.860 86.110 147.030 ;
        RECT 86.280 146.860 86.520 147.030 ;
        RECT 86.690 146.860 86.950 147.030 ;
        RECT 87.120 146.860 87.390 147.030 ;
        RECT 87.560 146.860 87.800 147.030 ;
        RECT 87.970 146.860 88.200 147.030 ;
        RECT 85.460 146.840 88.200 146.860 ;
        RECT 89.300 147.030 92.040 147.910 ;
        RECT 89.300 146.860 89.510 147.030 ;
        RECT 89.680 146.860 89.950 147.030 ;
        RECT 90.120 146.860 90.360 147.030 ;
        RECT 90.530 146.860 90.790 147.030 ;
        RECT 90.960 146.860 91.230 147.030 ;
        RECT 91.400 146.860 91.640 147.030 ;
        RECT 91.810 146.860 92.040 147.030 ;
        RECT 89.300 146.840 92.040 146.860 ;
        RECT 93.140 147.030 95.880 147.910 ;
        RECT 93.140 146.860 93.350 147.030 ;
        RECT 93.520 146.860 93.790 147.030 ;
        RECT 93.960 146.860 94.200 147.030 ;
        RECT 94.370 146.860 94.630 147.030 ;
        RECT 94.800 146.860 95.070 147.030 ;
        RECT 95.240 146.860 95.480 147.030 ;
        RECT 95.650 146.860 95.880 147.030 ;
        RECT 93.140 146.840 95.880 146.860 ;
        RECT 96.980 147.030 99.720 147.910 ;
        RECT 96.980 146.860 97.190 147.030 ;
        RECT 97.360 146.860 97.630 147.030 ;
        RECT 97.800 146.860 98.040 147.030 ;
        RECT 98.210 146.860 98.470 147.030 ;
        RECT 98.640 146.860 98.910 147.030 ;
        RECT 99.080 146.860 99.320 147.030 ;
        RECT 99.490 146.860 99.720 147.030 ;
        RECT 96.980 146.840 99.720 146.860 ;
        RECT 100.820 147.030 103.560 147.910 ;
        RECT 100.820 146.860 101.030 147.030 ;
        RECT 101.200 146.860 101.470 147.030 ;
        RECT 101.640 146.860 101.880 147.030 ;
        RECT 102.050 146.860 102.310 147.030 ;
        RECT 102.480 146.860 102.750 147.030 ;
        RECT 102.920 146.860 103.160 147.030 ;
        RECT 103.330 146.860 103.560 147.030 ;
        RECT 100.820 146.840 103.560 146.860 ;
        RECT 104.660 147.030 107.400 147.910 ;
        RECT 104.660 146.860 104.870 147.030 ;
        RECT 105.040 146.860 105.310 147.030 ;
        RECT 105.480 146.860 105.720 147.030 ;
        RECT 105.890 146.860 106.150 147.030 ;
        RECT 106.320 146.860 106.590 147.030 ;
        RECT 106.760 146.860 107.000 147.030 ;
        RECT 107.170 146.860 107.400 147.030 ;
        RECT 104.660 146.840 107.400 146.860 ;
        RECT 108.500 147.030 111.240 147.910 ;
        RECT 108.500 146.860 108.710 147.030 ;
        RECT 108.880 146.860 109.150 147.030 ;
        RECT 109.320 146.860 109.560 147.030 ;
        RECT 109.730 146.860 109.990 147.030 ;
        RECT 110.160 146.860 110.430 147.030 ;
        RECT 110.600 146.860 110.840 147.030 ;
        RECT 111.010 146.860 111.240 147.030 ;
        RECT 108.500 146.840 111.240 146.860 ;
        RECT 112.340 147.030 115.080 147.910 ;
        RECT 112.340 146.860 112.550 147.030 ;
        RECT 112.720 146.860 112.990 147.030 ;
        RECT 113.160 146.860 113.400 147.030 ;
        RECT 113.570 146.860 113.830 147.030 ;
        RECT 114.000 146.860 114.270 147.030 ;
        RECT 114.440 146.860 114.680 147.030 ;
        RECT 114.850 146.860 115.080 147.030 ;
        RECT 112.340 146.840 115.080 146.860 ;
        RECT 116.180 147.030 118.920 147.910 ;
        RECT 116.180 146.860 116.390 147.030 ;
        RECT 116.560 146.860 116.830 147.030 ;
        RECT 117.000 146.860 117.240 147.030 ;
        RECT 117.410 146.860 117.670 147.030 ;
        RECT 117.840 146.860 118.110 147.030 ;
        RECT 118.280 146.860 118.520 147.030 ;
        RECT 118.690 146.860 118.920 147.030 ;
        RECT 116.180 146.840 118.920 146.860 ;
        RECT 120.020 147.030 122.760 147.910 ;
        RECT 120.020 146.860 120.230 147.030 ;
        RECT 120.400 146.860 120.670 147.030 ;
        RECT 120.840 146.860 121.080 147.030 ;
        RECT 121.250 146.860 121.510 147.030 ;
        RECT 121.680 146.860 121.950 147.030 ;
        RECT 122.120 146.860 122.360 147.030 ;
        RECT 122.530 146.860 122.760 147.030 ;
        RECT 120.020 146.840 122.760 146.860 ;
        RECT 123.860 147.030 126.600 147.910 ;
        RECT 123.860 146.860 124.070 147.030 ;
        RECT 124.240 146.860 124.510 147.030 ;
        RECT 124.680 146.860 124.920 147.030 ;
        RECT 125.090 146.860 125.350 147.030 ;
        RECT 125.520 146.860 125.790 147.030 ;
        RECT 125.960 146.860 126.200 147.030 ;
        RECT 126.370 146.860 126.600 147.030 ;
        RECT 123.860 146.840 126.600 146.860 ;
        RECT 127.700 147.030 130.440 147.910 ;
        RECT 127.700 146.860 127.910 147.030 ;
        RECT 128.080 146.860 128.350 147.030 ;
        RECT 128.520 146.860 128.760 147.030 ;
        RECT 128.930 146.860 129.190 147.030 ;
        RECT 129.360 146.860 129.630 147.030 ;
        RECT 129.800 146.860 130.040 147.030 ;
        RECT 130.210 146.860 130.440 147.030 ;
        RECT 127.700 146.840 130.440 146.860 ;
        RECT 131.540 147.030 134.280 147.910 ;
        RECT 131.540 146.860 131.750 147.030 ;
        RECT 131.920 146.860 132.190 147.030 ;
        RECT 132.360 146.860 132.600 147.030 ;
        RECT 132.770 146.860 133.030 147.030 ;
        RECT 133.200 146.860 133.470 147.030 ;
        RECT 133.640 146.860 133.880 147.030 ;
        RECT 134.050 146.860 134.280 147.030 ;
        RECT 131.540 146.840 134.280 146.860 ;
        RECT 135.380 147.030 138.120 147.910 ;
        RECT 139.740 147.900 140.070 148.890 ;
        RECT 135.380 146.860 135.590 147.030 ;
        RECT 135.760 146.860 136.030 147.030 ;
        RECT 136.200 146.860 136.440 147.030 ;
        RECT 136.610 146.860 136.870 147.030 ;
        RECT 137.040 146.860 137.310 147.030 ;
        RECT 137.480 146.860 137.720 147.030 ;
        RECT 137.890 146.860 138.120 147.030 ;
        RECT 135.380 146.840 138.120 146.860 ;
        RECT 138.970 147.030 140.420 147.900 ;
        RECT 138.970 146.860 139.220 147.030 ;
        RECT 139.390 146.860 139.580 147.030 ;
        RECT 139.750 146.860 140.020 147.030 ;
        RECT 140.190 146.860 140.420 147.030 ;
        RECT 138.970 146.830 140.420 146.860 ;
        RECT 5.760 146.430 5.920 146.610 ;
        RECT 6.090 146.430 6.400 146.610 ;
        RECT 6.570 146.430 6.880 146.610 ;
        RECT 7.050 146.430 7.360 146.610 ;
        RECT 7.530 146.430 7.840 146.610 ;
        RECT 8.010 146.430 8.320 146.610 ;
        RECT 8.490 146.430 8.800 146.610 ;
        RECT 8.970 146.430 9.280 146.610 ;
        RECT 9.450 146.430 9.760 146.610 ;
        RECT 9.930 146.430 10.240 146.610 ;
        RECT 10.410 146.430 10.720 146.610 ;
        RECT 10.890 146.430 11.200 146.610 ;
        RECT 11.370 146.430 11.680 146.610 ;
        RECT 11.850 146.430 12.160 146.610 ;
        RECT 12.330 146.430 12.640 146.610 ;
        RECT 12.810 146.430 13.120 146.610 ;
        RECT 13.290 146.430 13.600 146.610 ;
        RECT 13.770 146.430 14.080 146.610 ;
        RECT 14.250 146.430 14.560 146.610 ;
        RECT 14.730 146.430 15.040 146.610 ;
        RECT 15.210 146.430 15.520 146.610 ;
        RECT 15.690 146.430 16.000 146.610 ;
        RECT 16.170 146.430 16.480 146.610 ;
        RECT 16.650 146.430 16.960 146.610 ;
        RECT 17.130 146.430 17.440 146.610 ;
        RECT 17.610 146.600 17.760 146.610 ;
        RECT 18.240 146.600 18.400 146.610 ;
        RECT 17.610 146.430 17.920 146.600 ;
        RECT 18.090 146.430 18.400 146.600 ;
        RECT 18.570 146.430 18.880 146.610 ;
        RECT 19.050 146.430 19.360 146.610 ;
        RECT 19.530 146.430 19.840 146.610 ;
        RECT 20.010 146.430 20.320 146.610 ;
        RECT 20.490 146.430 20.800 146.610 ;
        RECT 20.970 146.430 21.280 146.610 ;
        RECT 21.450 146.430 21.760 146.610 ;
        RECT 21.930 146.430 22.240 146.610 ;
        RECT 22.410 146.430 22.720 146.610 ;
        RECT 22.890 146.430 23.200 146.610 ;
        RECT 23.370 146.430 23.680 146.610 ;
        RECT 23.850 146.430 24.160 146.610 ;
        RECT 24.330 146.430 24.640 146.610 ;
        RECT 24.810 146.430 25.120 146.610 ;
        RECT 25.290 146.430 25.600 146.610 ;
        RECT 25.770 146.430 26.080 146.610 ;
        RECT 26.250 146.430 26.560 146.610 ;
        RECT 26.730 146.430 27.040 146.610 ;
        RECT 27.210 146.430 27.520 146.610 ;
        RECT 27.690 146.430 28.000 146.610 ;
        RECT 28.170 146.430 28.480 146.610 ;
        RECT 28.650 146.430 28.960 146.610 ;
        RECT 29.130 146.430 29.440 146.610 ;
        RECT 29.610 146.430 29.920 146.610 ;
        RECT 30.090 146.430 30.400 146.610 ;
        RECT 30.570 146.430 30.880 146.610 ;
        RECT 31.050 146.430 31.360 146.610 ;
        RECT 31.530 146.430 31.840 146.610 ;
        RECT 32.010 146.430 32.320 146.610 ;
        RECT 32.490 146.430 32.800 146.610 ;
        RECT 32.970 146.430 33.280 146.610 ;
        RECT 33.450 146.430 33.760 146.610 ;
        RECT 33.930 146.430 34.240 146.610 ;
        RECT 34.410 146.430 34.720 146.610 ;
        RECT 34.890 146.430 35.200 146.610 ;
        RECT 35.370 146.430 35.680 146.610 ;
        RECT 35.850 146.600 36.000 146.610 ;
        RECT 36.480 146.600 36.640 146.610 ;
        RECT 35.850 146.430 36.160 146.600 ;
        RECT 36.330 146.430 36.640 146.600 ;
        RECT 36.810 146.430 37.120 146.610 ;
        RECT 37.290 146.430 37.600 146.610 ;
        RECT 37.770 146.430 38.080 146.610 ;
        RECT 38.250 146.430 38.560 146.610 ;
        RECT 38.730 146.430 39.040 146.610 ;
        RECT 39.210 146.430 39.520 146.610 ;
        RECT 39.690 146.430 40.000 146.610 ;
        RECT 40.170 146.430 40.480 146.610 ;
        RECT 40.650 146.430 40.960 146.610 ;
        RECT 41.130 146.430 41.440 146.610 ;
        RECT 41.610 146.430 41.920 146.610 ;
        RECT 42.090 146.430 42.400 146.610 ;
        RECT 42.570 146.430 42.880 146.610 ;
        RECT 43.050 146.430 43.360 146.610 ;
        RECT 43.530 146.600 43.680 146.610 ;
        RECT 44.160 146.600 44.320 146.610 ;
        RECT 43.530 146.430 43.840 146.600 ;
        RECT 44.010 146.430 44.320 146.600 ;
        RECT 44.490 146.430 44.800 146.610 ;
        RECT 44.970 146.430 45.280 146.610 ;
        RECT 45.450 146.430 45.760 146.610 ;
        RECT 45.930 146.430 46.240 146.610 ;
        RECT 46.410 146.430 46.720 146.610 ;
        RECT 46.890 146.430 47.200 146.610 ;
        RECT 47.370 146.430 47.680 146.610 ;
        RECT 47.850 146.430 48.160 146.610 ;
        RECT 48.330 146.430 48.640 146.610 ;
        RECT 48.810 146.430 49.120 146.610 ;
        RECT 49.290 146.430 49.600 146.610 ;
        RECT 49.770 146.430 50.080 146.610 ;
        RECT 50.250 146.430 50.560 146.610 ;
        RECT 50.730 146.430 51.040 146.610 ;
        RECT 51.210 146.430 51.520 146.610 ;
        RECT 51.690 146.430 52.000 146.610 ;
        RECT 52.170 146.430 52.480 146.610 ;
        RECT 52.650 146.430 52.960 146.610 ;
        RECT 53.130 146.430 53.440 146.610 ;
        RECT 53.610 146.430 53.920 146.610 ;
        RECT 54.090 146.430 54.400 146.610 ;
        RECT 54.570 146.430 54.880 146.610 ;
        RECT 55.050 146.430 55.360 146.610 ;
        RECT 55.530 146.430 55.840 146.610 ;
        RECT 56.010 146.430 56.320 146.610 ;
        RECT 56.490 146.430 56.800 146.610 ;
        RECT 56.970 146.430 57.280 146.610 ;
        RECT 57.450 146.430 57.760 146.610 ;
        RECT 57.930 146.430 58.240 146.610 ;
        RECT 58.410 146.430 58.720 146.610 ;
        RECT 58.890 146.430 59.200 146.610 ;
        RECT 59.370 146.430 59.680 146.610 ;
        RECT 59.850 146.430 60.160 146.610 ;
        RECT 60.330 146.430 60.640 146.610 ;
        RECT 60.810 146.430 61.120 146.610 ;
        RECT 61.290 146.430 61.600 146.610 ;
        RECT 61.770 146.430 62.080 146.610 ;
        RECT 62.250 146.430 62.560 146.610 ;
        RECT 62.730 146.430 63.040 146.610 ;
        RECT 63.210 146.430 63.520 146.610 ;
        RECT 63.690 146.430 64.000 146.610 ;
        RECT 64.170 146.430 64.480 146.610 ;
        RECT 64.650 146.430 64.960 146.610 ;
        RECT 65.130 146.430 65.440 146.610 ;
        RECT 65.610 146.430 65.920 146.610 ;
        RECT 66.090 146.430 66.400 146.610 ;
        RECT 66.570 146.430 66.880 146.610 ;
        RECT 67.050 146.430 67.360 146.610 ;
        RECT 67.530 146.430 67.840 146.610 ;
        RECT 68.010 146.430 68.320 146.610 ;
        RECT 68.490 146.430 68.800 146.610 ;
        RECT 68.970 146.430 69.280 146.610 ;
        RECT 69.450 146.430 69.760 146.610 ;
        RECT 69.930 146.430 70.240 146.610 ;
        RECT 70.410 146.430 70.720 146.610 ;
        RECT 70.890 146.430 71.200 146.610 ;
        RECT 71.370 146.430 71.680 146.610 ;
        RECT 71.850 146.430 72.160 146.610 ;
        RECT 72.330 146.430 72.640 146.610 ;
        RECT 72.810 146.430 73.120 146.610 ;
        RECT 73.290 146.430 73.600 146.610 ;
        RECT 73.770 146.430 74.080 146.610 ;
        RECT 74.250 146.430 74.560 146.610 ;
        RECT 74.730 146.430 75.040 146.610 ;
        RECT 75.210 146.430 75.520 146.610 ;
        RECT 75.690 146.430 76.000 146.610 ;
        RECT 76.170 146.430 76.480 146.610 ;
        RECT 76.650 146.430 76.960 146.610 ;
        RECT 77.130 146.430 77.440 146.610 ;
        RECT 77.610 146.430 77.920 146.610 ;
        RECT 78.090 146.430 78.400 146.610 ;
        RECT 78.570 146.430 78.880 146.610 ;
        RECT 79.050 146.430 79.360 146.610 ;
        RECT 79.530 146.430 79.840 146.610 ;
        RECT 80.010 146.430 80.320 146.610 ;
        RECT 80.490 146.430 80.800 146.610 ;
        RECT 80.970 146.430 81.280 146.610 ;
        RECT 81.450 146.430 81.760 146.610 ;
        RECT 81.930 146.430 82.240 146.610 ;
        RECT 82.410 146.430 82.720 146.610 ;
        RECT 82.890 146.430 83.200 146.610 ;
        RECT 83.370 146.430 83.680 146.610 ;
        RECT 83.850 146.430 84.160 146.610 ;
        RECT 84.330 146.430 84.640 146.610 ;
        RECT 84.810 146.430 85.120 146.610 ;
        RECT 85.290 146.600 85.440 146.610 ;
        RECT 85.920 146.600 86.080 146.610 ;
        RECT 85.290 146.430 85.600 146.600 ;
        RECT 85.770 146.430 86.080 146.600 ;
        RECT 86.250 146.430 86.560 146.610 ;
        RECT 86.730 146.430 87.040 146.610 ;
        RECT 87.210 146.430 87.520 146.610 ;
        RECT 87.690 146.430 88.000 146.610 ;
        RECT 88.170 146.430 88.480 146.610 ;
        RECT 88.650 146.430 88.960 146.610 ;
        RECT 89.130 146.430 89.440 146.610 ;
        RECT 89.610 146.430 89.920 146.610 ;
        RECT 90.090 146.430 90.400 146.610 ;
        RECT 90.570 146.430 90.880 146.610 ;
        RECT 91.050 146.430 91.360 146.610 ;
        RECT 91.530 146.430 91.840 146.610 ;
        RECT 92.010 146.430 92.320 146.610 ;
        RECT 92.490 146.430 92.800 146.610 ;
        RECT 92.970 146.430 93.280 146.610 ;
        RECT 93.450 146.430 93.760 146.610 ;
        RECT 93.930 146.430 94.240 146.610 ;
        RECT 94.410 146.430 94.720 146.610 ;
        RECT 94.890 146.430 95.200 146.610 ;
        RECT 95.370 146.430 95.680 146.610 ;
        RECT 95.850 146.430 96.160 146.610 ;
        RECT 96.330 146.430 96.640 146.610 ;
        RECT 96.810 146.430 97.120 146.610 ;
        RECT 97.290 146.430 97.600 146.610 ;
        RECT 97.770 146.430 98.080 146.610 ;
        RECT 98.250 146.430 98.560 146.610 ;
        RECT 98.730 146.430 99.040 146.610 ;
        RECT 99.210 146.430 99.520 146.610 ;
        RECT 99.690 146.430 100.000 146.610 ;
        RECT 100.170 146.430 100.480 146.610 ;
        RECT 100.650 146.430 100.960 146.610 ;
        RECT 101.130 146.430 101.440 146.610 ;
        RECT 101.610 146.430 101.920 146.610 ;
        RECT 102.090 146.430 102.400 146.610 ;
        RECT 102.570 146.430 102.880 146.610 ;
        RECT 103.050 146.430 103.360 146.610 ;
        RECT 103.530 146.430 103.840 146.610 ;
        RECT 104.010 146.430 104.320 146.610 ;
        RECT 104.490 146.430 104.800 146.610 ;
        RECT 104.970 146.430 105.280 146.610 ;
        RECT 105.450 146.430 105.760 146.610 ;
        RECT 105.930 146.430 106.240 146.610 ;
        RECT 106.410 146.430 106.720 146.610 ;
        RECT 106.890 146.430 107.200 146.610 ;
        RECT 107.370 146.430 107.680 146.610 ;
        RECT 107.850 146.430 108.160 146.610 ;
        RECT 108.330 146.430 108.640 146.610 ;
        RECT 108.810 146.430 109.120 146.610 ;
        RECT 109.290 146.430 109.600 146.610 ;
        RECT 109.770 146.430 110.080 146.610 ;
        RECT 110.250 146.430 110.560 146.610 ;
        RECT 110.730 146.430 111.040 146.610 ;
        RECT 111.210 146.430 111.520 146.610 ;
        RECT 111.690 146.430 112.000 146.610 ;
        RECT 112.170 146.430 112.480 146.610 ;
        RECT 112.650 146.430 112.960 146.610 ;
        RECT 113.130 146.430 113.440 146.610 ;
        RECT 113.610 146.430 113.920 146.610 ;
        RECT 114.090 146.430 114.400 146.610 ;
        RECT 114.570 146.430 114.880 146.610 ;
        RECT 115.050 146.430 115.360 146.610 ;
        RECT 115.530 146.430 115.840 146.610 ;
        RECT 116.010 146.430 116.320 146.610 ;
        RECT 116.490 146.430 116.800 146.610 ;
        RECT 116.970 146.430 117.280 146.610 ;
        RECT 117.450 146.430 117.760 146.610 ;
        RECT 117.930 146.430 118.240 146.610 ;
        RECT 118.410 146.430 118.720 146.610 ;
        RECT 118.890 146.430 119.200 146.610 ;
        RECT 119.370 146.430 119.680 146.610 ;
        RECT 119.850 146.430 120.160 146.610 ;
        RECT 120.330 146.430 120.640 146.610 ;
        RECT 120.810 146.430 121.120 146.610 ;
        RECT 121.290 146.430 121.600 146.610 ;
        RECT 121.770 146.430 122.080 146.610 ;
        RECT 122.250 146.430 122.560 146.610 ;
        RECT 122.730 146.430 123.040 146.610 ;
        RECT 123.210 146.430 123.520 146.610 ;
        RECT 123.690 146.430 124.000 146.610 ;
        RECT 124.170 146.430 124.480 146.610 ;
        RECT 124.650 146.430 124.960 146.610 ;
        RECT 125.130 146.430 125.440 146.610 ;
        RECT 125.610 146.430 125.920 146.610 ;
        RECT 126.090 146.430 126.400 146.610 ;
        RECT 126.570 146.430 126.880 146.610 ;
        RECT 127.050 146.430 127.360 146.610 ;
        RECT 127.530 146.430 127.840 146.610 ;
        RECT 128.010 146.430 128.320 146.610 ;
        RECT 128.490 146.430 128.800 146.610 ;
        RECT 128.970 146.430 129.280 146.610 ;
        RECT 129.450 146.430 129.760 146.610 ;
        RECT 129.930 146.430 130.240 146.610 ;
        RECT 130.410 146.430 130.720 146.610 ;
        RECT 130.890 146.430 131.200 146.610 ;
        RECT 131.370 146.430 131.680 146.610 ;
        RECT 131.850 146.430 132.160 146.610 ;
        RECT 132.330 146.430 132.640 146.610 ;
        RECT 132.810 146.430 133.120 146.610 ;
        RECT 133.290 146.430 133.600 146.610 ;
        RECT 133.770 146.430 134.080 146.610 ;
        RECT 134.250 146.430 134.560 146.610 ;
        RECT 134.730 146.430 135.040 146.610 ;
        RECT 135.210 146.430 135.520 146.610 ;
        RECT 135.690 146.430 136.000 146.610 ;
        RECT 136.170 146.430 136.480 146.610 ;
        RECT 136.650 146.430 136.960 146.610 ;
        RECT 137.130 146.430 137.440 146.610 ;
        RECT 137.610 146.430 137.920 146.610 ;
        RECT 138.090 146.430 138.400 146.610 ;
        RECT 138.570 146.430 138.880 146.610 ;
        RECT 139.050 146.430 139.360 146.610 ;
        RECT 139.530 146.430 139.840 146.610 ;
        RECT 140.010 146.430 140.320 146.610 ;
        RECT 140.490 146.430 140.800 146.610 ;
        RECT 140.970 146.430 141.280 146.610 ;
        RECT 141.450 146.430 141.600 146.610 ;
        RECT 6.260 146.180 9.000 146.200 ;
        RECT 6.260 146.010 6.470 146.180 ;
        RECT 6.640 146.010 6.910 146.180 ;
        RECT 7.080 146.010 7.320 146.180 ;
        RECT 7.490 146.010 7.750 146.180 ;
        RECT 7.920 146.010 8.190 146.180 ;
        RECT 8.360 146.010 8.600 146.180 ;
        RECT 8.770 146.010 9.000 146.180 ;
        RECT 6.260 145.130 9.000 146.010 ;
        RECT 10.780 146.130 11.430 146.240 ;
        RECT 10.780 145.960 10.840 146.130 ;
        RECT 11.010 145.960 11.200 146.130 ;
        RECT 11.370 145.960 11.430 146.130 ;
        RECT 10.780 145.900 11.430 145.960 ;
        RECT 10.780 145.630 11.180 145.900 ;
      LAYER li1 ;
        RECT 12.090 145.630 12.670 146.270 ;
      LAYER li1 ;
        RECT 13.460 146.180 16.200 146.200 ;
        RECT 13.460 146.010 13.670 146.180 ;
        RECT 13.840 146.010 14.110 146.180 ;
        RECT 14.280 146.010 14.520 146.180 ;
        RECT 14.690 146.010 14.950 146.180 ;
        RECT 15.120 146.010 15.390 146.180 ;
        RECT 15.560 146.010 15.800 146.180 ;
        RECT 15.970 146.010 16.200 146.180 ;
        RECT 6.500 143.810 6.830 144.480 ;
        RECT 7.230 144.150 7.560 145.130 ;
        RECT 7.780 143.810 8.110 144.480 ;
        RECT 8.510 144.150 8.840 145.130 ;
      LAYER li1 ;
        RECT 12.090 144.220 12.360 145.630 ;
      LAYER li1 ;
        RECT 13.460 145.130 16.200 146.010 ;
      LAYER li1 ;
        RECT 11.600 143.950 12.360 144.220 ;
      LAYER li1 ;
        RECT 6.340 142.810 9.070 143.810 ;
      LAYER li1 ;
        RECT 11.600 142.950 11.930 143.950 ;
      LAYER li1 ;
        RECT 13.700 143.810 14.030 144.480 ;
        RECT 14.430 144.150 14.760 145.130 ;
        RECT 14.980 143.810 15.310 144.480 ;
        RECT 15.710 144.150 16.040 145.130 ;
        RECT 18.360 143.920 18.610 146.190 ;
        RECT 18.790 146.130 19.740 146.210 ;
        RECT 18.790 145.960 18.820 146.130 ;
        RECT 18.990 145.960 19.180 146.130 ;
        RECT 19.350 145.960 19.540 146.130 ;
        RECT 19.710 145.960 19.740 146.130 ;
        RECT 18.790 145.380 19.740 145.960 ;
        RECT 19.920 145.400 20.250 146.190 ;
        RECT 19.930 144.900 20.250 145.400 ;
        RECT 20.480 146.130 20.730 146.160 ;
        RECT 20.480 145.960 20.510 146.130 ;
        RECT 20.680 145.960 20.730 146.130 ;
        RECT 20.480 145.080 20.730 145.960 ;
        RECT 20.910 144.900 21.080 146.210 ;
        RECT 23.850 146.130 24.180 146.160 ;
        RECT 19.930 144.730 21.080 144.900 ;
        RECT 21.260 145.740 23.250 146.070 ;
        RECT 19.420 143.920 19.750 144.350 ;
        RECT 12.340 143.080 12.750 143.520 ;
        RECT 12.100 142.740 12.750 143.080 ;
        RECT 13.540 142.810 16.270 143.810 ;
        RECT 18.360 143.750 19.750 143.920 ;
        RECT 18.360 143.070 18.620 143.750 ;
        RECT 18.810 142.820 19.400 143.570 ;
        RECT 19.580 142.890 19.750 143.750 ;
        RECT 19.930 143.070 20.180 144.730 ;
      LAYER li1 ;
        RECT 20.750 143.980 21.080 144.550 ;
      LAYER li1 ;
        RECT 21.260 143.800 21.430 145.740 ;
        RECT 20.360 143.630 21.430 143.800 ;
        RECT 20.360 142.890 20.530 143.630 ;
        RECT 21.610 143.450 21.780 145.560 ;
        RECT 21.960 143.540 22.130 145.740 ;
        RECT 22.310 145.060 22.640 145.560 ;
        RECT 22.310 143.590 22.480 145.060 ;
        RECT 23.080 144.780 23.250 145.740 ;
        RECT 23.430 145.130 23.670 146.010 ;
        RECT 23.850 145.960 23.880 146.130 ;
        RECT 24.050 145.960 24.180 146.130 ;
        RECT 23.850 145.310 24.180 145.960 ;
        RECT 25.320 146.130 26.270 146.160 ;
        RECT 25.320 145.960 25.350 146.130 ;
        RECT 25.520 145.960 25.710 146.130 ;
        RECT 25.880 145.960 26.070 146.130 ;
        RECT 26.240 145.960 26.270 146.130 ;
        RECT 24.810 145.300 25.140 145.560 ;
        RECT 24.360 145.130 25.140 145.300 ;
        RECT 25.320 145.130 26.270 145.960 ;
        RECT 26.940 146.050 28.070 146.260 ;
        RECT 28.250 146.130 29.200 146.160 ;
        RECT 26.940 145.300 27.110 146.050 ;
        RECT 28.250 145.960 28.280 146.130 ;
        RECT 28.450 145.960 28.640 146.130 ;
        RECT 28.810 145.960 29.000 146.130 ;
        RECT 29.170 145.960 29.200 146.130 ;
        RECT 27.290 145.480 27.900 145.870 ;
        RECT 26.940 145.130 27.550 145.300 ;
        RECT 23.430 144.960 24.530 145.130 ;
        RECT 24.710 144.780 27.200 144.950 ;
        RECT 22.660 144.430 22.900 144.620 ;
        RECT 23.080 144.610 24.880 144.780 ;
        RECT 25.060 144.430 26.690 144.600 ;
        RECT 26.870 144.540 27.200 144.780 ;
        RECT 22.660 144.260 25.230 144.430 ;
        RECT 26.520 144.330 26.690 144.430 ;
        RECT 27.380 144.330 27.550 145.130 ;
        RECT 22.660 143.950 22.900 144.260 ;
        RECT 23.380 143.770 24.110 144.080 ;
      LAYER li1 ;
        RECT 25.410 144.010 26.340 144.250 ;
      LAYER li1 ;
        RECT 19.580 142.720 20.530 142.890 ;
        RECT 20.710 142.820 21.250 143.450 ;
        RECT 21.430 142.950 21.780 143.450 ;
        RECT 22.310 143.420 24.560 143.590 ;
        RECT 22.310 142.950 22.560 143.420 ;
        RECT 23.100 142.820 24.050 143.240 ;
        RECT 24.230 142.720 24.560 143.420 ;
        RECT 25.040 142.820 25.990 143.830 ;
      LAYER li1 ;
        RECT 26.170 143.460 26.340 144.010 ;
      LAYER li1 ;
        RECT 26.520 144.160 27.550 144.330 ;
        RECT 27.730 144.940 27.900 145.480 ;
        RECT 28.250 145.120 29.200 145.960 ;
        RECT 29.540 145.710 29.790 146.210 ;
        RECT 29.970 146.130 30.920 146.190 ;
        RECT 33.370 146.180 34.820 146.210 ;
        RECT 29.970 145.960 30.000 146.130 ;
        RECT 30.170 145.960 30.360 146.130 ;
        RECT 30.530 145.960 30.720 146.130 ;
        RECT 30.890 145.960 30.920 146.130 ;
        RECT 29.970 145.810 30.920 145.960 ;
        RECT 31.540 146.130 32.480 146.160 ;
        RECT 31.540 145.960 31.560 146.130 ;
        RECT 31.730 145.960 31.920 146.130 ;
        RECT 32.090 145.960 32.280 146.130 ;
        RECT 32.450 145.960 32.480 146.130 ;
        RECT 29.620 145.630 29.790 145.710 ;
        RECT 29.620 145.460 30.800 145.630 ;
        RECT 29.650 145.130 29.980 145.280 ;
        RECT 29.650 144.940 30.450 145.130 ;
        RECT 27.730 144.770 30.450 144.940 ;
        RECT 26.520 144.000 27.030 144.160 ;
        RECT 27.730 143.930 27.900 144.770 ;
        RECT 28.550 144.280 28.880 144.590 ;
        RECT 30.120 144.460 30.450 144.770 ;
        RECT 30.630 144.280 30.800 145.460 ;
        RECT 28.550 144.110 30.800 144.280 ;
        RECT 31.110 144.850 31.360 145.820 ;
        RECT 31.540 145.030 32.480 145.960 ;
        RECT 33.370 146.010 33.620 146.180 ;
        RECT 33.790 146.010 33.980 146.180 ;
        RECT 34.150 146.010 34.420 146.180 ;
        RECT 34.590 146.010 34.820 146.180 ;
        RECT 33.370 145.140 34.820 146.010 ;
        RECT 31.110 144.680 32.480 144.850 ;
        RECT 28.550 144.000 28.880 144.110 ;
        RECT 27.270 143.640 27.900 143.930 ;
      LAYER li1 ;
        RECT 29.130 143.460 29.400 143.490 ;
        RECT 26.170 143.290 29.400 143.460 ;
        RECT 26.530 143.010 29.400 143.290 ;
      LAYER li1 ;
        RECT 29.580 142.820 30.170 143.930 ;
        RECT 30.360 143.430 30.690 144.110 ;
        RECT 31.110 143.930 31.320 144.680 ;
        RECT 32.150 144.180 32.480 144.680 ;
        RECT 30.990 143.430 31.320 143.930 ;
        RECT 31.500 142.820 32.450 143.930 ;
        RECT 33.600 143.700 33.930 144.480 ;
        RECT 34.140 144.150 34.470 145.140 ;
      LAYER li1 ;
        RECT 36.600 144.630 37.030 146.210 ;
      LAYER li1 ;
        RECT 37.210 146.130 37.770 146.210 ;
        RECT 37.210 145.960 37.220 146.130 ;
        RECT 37.390 145.960 37.580 146.130 ;
        RECT 37.750 145.960 37.770 146.130 ;
        RECT 37.210 144.630 37.770 145.960 ;
        RECT 39.380 146.180 42.120 146.200 ;
        RECT 39.380 146.010 39.590 146.180 ;
        RECT 39.760 146.010 40.030 146.180 ;
        RECT 40.200 146.010 40.440 146.180 ;
        RECT 40.610 146.010 40.870 146.180 ;
        RECT 41.040 146.010 41.310 146.180 ;
        RECT 41.480 146.010 41.720 146.180 ;
        RECT 41.890 146.010 42.120 146.180 ;
        RECT 33.600 143.300 34.900 143.700 ;
        RECT 33.290 142.820 34.900 143.300 ;
      LAYER li1 ;
        RECT 36.600 142.950 36.850 144.630 ;
      LAYER li1 ;
        RECT 37.160 143.740 37.490 144.200 ;
      LAYER li1 ;
        RECT 37.950 143.920 38.280 145.710 ;
      LAYER li1 ;
        RECT 38.460 143.740 38.710 145.460 ;
        RECT 39.380 145.130 42.120 146.010 ;
        RECT 44.380 146.130 45.030 146.240 ;
        RECT 44.380 145.960 44.440 146.130 ;
        RECT 44.610 145.960 44.800 146.130 ;
        RECT 44.970 145.960 45.030 146.130 ;
        RECT 47.060 146.180 49.800 146.200 ;
        RECT 47.060 146.010 47.270 146.180 ;
        RECT 47.440 146.010 47.710 146.180 ;
        RECT 47.880 146.010 48.120 146.180 ;
        RECT 48.290 146.010 48.550 146.180 ;
        RECT 48.720 146.010 48.990 146.180 ;
        RECT 49.160 146.010 49.400 146.180 ;
        RECT 49.570 146.010 49.800 146.180 ;
        RECT 44.380 145.900 45.030 145.960 ;
        RECT 44.380 145.630 44.780 145.900 ;
        RECT 39.620 143.810 39.950 144.480 ;
        RECT 40.350 144.150 40.680 145.130 ;
        RECT 40.900 143.810 41.230 144.480 ;
        RECT 41.630 144.150 41.960 145.130 ;
      LAYER li1 ;
        RECT 45.240 144.640 45.490 145.980 ;
      LAYER li1 ;
        RECT 47.060 145.130 49.800 146.010 ;
      LAYER li1 ;
        RECT 44.780 144.390 45.490 144.640 ;
      LAYER li1 ;
        RECT 37.160 143.570 38.710 143.740 ;
        RECT 37.030 142.820 38.280 143.390 ;
        RECT 38.460 142.950 38.710 143.570 ;
        RECT 39.460 142.810 42.190 143.810 ;
      LAYER li1 ;
        RECT 44.780 143.520 45.030 144.390 ;
      LAYER li1 ;
        RECT 47.300 143.810 47.630 144.480 ;
        RECT 48.030 144.150 48.360 145.130 ;
        RECT 48.580 143.810 48.910 144.480 ;
        RECT 49.310 144.150 49.640 145.130 ;
      LAYER li1 ;
        RECT 50.520 144.630 50.950 146.210 ;
      LAYER li1 ;
        RECT 51.130 146.130 51.690 146.210 ;
        RECT 51.130 145.960 51.140 146.130 ;
        RECT 51.310 145.960 51.500 146.130 ;
        RECT 51.670 145.960 51.690 146.130 ;
        RECT 51.130 144.630 51.690 145.960 ;
        RECT 53.300 146.180 56.040 146.200 ;
        RECT 53.300 146.010 53.510 146.180 ;
        RECT 53.680 146.010 53.950 146.180 ;
        RECT 54.120 146.010 54.360 146.180 ;
        RECT 54.530 146.010 54.790 146.180 ;
        RECT 54.960 146.010 55.230 146.180 ;
        RECT 55.400 146.010 55.640 146.180 ;
        RECT 55.810 146.010 56.040 146.180 ;
      LAYER li1 ;
        RECT 44.450 142.880 45.030 143.520 ;
      LAYER li1 ;
        RECT 45.940 143.080 46.350 143.520 ;
        RECT 45.700 142.740 46.350 143.080 ;
        RECT 47.140 142.810 49.870 143.810 ;
      LAYER li1 ;
        RECT 50.520 142.950 50.770 144.630 ;
      LAYER li1 ;
        RECT 51.080 143.740 51.410 144.200 ;
      LAYER li1 ;
        RECT 51.870 143.920 52.200 145.710 ;
      LAYER li1 ;
        RECT 52.380 143.740 52.630 145.460 ;
        RECT 53.300 145.130 56.040 146.010 ;
        RECT 57.140 146.180 59.880 146.200 ;
        RECT 57.140 146.010 57.350 146.180 ;
        RECT 57.520 146.010 57.790 146.180 ;
        RECT 57.960 146.010 58.200 146.180 ;
        RECT 58.370 146.010 58.630 146.180 ;
        RECT 58.800 146.010 59.070 146.180 ;
        RECT 59.240 146.010 59.480 146.180 ;
        RECT 59.650 146.010 59.880 146.180 ;
        RECT 57.140 145.130 59.880 146.010 ;
        RECT 61.110 146.130 61.700 146.160 ;
        RECT 61.110 145.960 61.140 146.130 ;
        RECT 61.310 145.960 61.500 146.130 ;
        RECT 61.670 145.960 61.700 146.130 ;
        RECT 53.540 143.810 53.870 144.480 ;
        RECT 54.270 144.150 54.600 145.130 ;
        RECT 54.820 143.810 55.150 144.480 ;
        RECT 55.550 144.150 55.880 145.130 ;
        RECT 57.380 143.810 57.710 144.480 ;
        RECT 58.110 144.150 58.440 145.130 ;
        RECT 58.660 143.810 58.990 144.480 ;
        RECT 59.390 144.150 59.720 145.130 ;
        RECT 60.590 144.980 60.920 145.910 ;
        RECT 61.110 145.180 61.700 145.960 ;
        RECT 61.880 146.090 63.320 146.260 ;
        RECT 61.880 144.980 62.050 146.090 ;
        RECT 60.590 144.810 62.050 144.980 ;
        RECT 51.080 143.570 52.630 143.740 ;
        RECT 50.950 142.820 52.200 143.390 ;
        RECT 52.380 142.950 52.630 143.570 ;
        RECT 53.380 142.810 56.110 143.810 ;
        RECT 57.220 142.810 59.950 143.810 ;
        RECT 60.590 142.950 60.860 144.810 ;
      LAYER li1 ;
        RECT 61.040 143.630 61.370 144.600 ;
      LAYER li1 ;
        RECT 61.720 144.310 62.050 144.810 ;
        RECT 62.230 144.600 62.480 145.910 ;
        RECT 62.720 145.290 62.970 145.910 ;
        RECT 63.150 145.640 63.320 146.090 ;
        RECT 63.500 146.130 63.830 146.160 ;
        RECT 63.500 145.960 63.530 146.130 ;
        RECT 63.700 145.960 63.830 146.130 ;
        RECT 63.500 145.820 63.830 145.960 ;
        RECT 64.010 146.090 65.750 146.260 ;
        RECT 64.010 145.640 64.180 146.090 ;
        RECT 63.150 145.470 64.180 145.640 ;
        RECT 64.360 145.290 64.530 145.910 ;
        RECT 65.060 145.650 65.390 145.910 ;
        RECT 62.720 145.120 64.530 145.290 ;
        RECT 64.710 145.120 64.930 145.450 ;
        RECT 64.360 144.940 64.530 145.120 ;
        RECT 62.230 144.370 62.760 144.600 ;
        RECT 62.230 143.450 62.500 144.370 ;
      LAYER li1 ;
        RECT 63.180 144.070 63.720 144.940 ;
      LAYER li1 ;
        RECT 64.360 144.770 64.580 144.940 ;
        RECT 61.040 142.820 61.990 143.450 ;
        RECT 62.170 142.950 62.500 143.450 ;
        RECT 62.680 142.820 63.270 143.700 ;
      LAYER li1 ;
        RECT 63.550 143.080 63.720 144.070 ;
        RECT 63.900 143.260 64.230 144.560 ;
      LAYER li1 ;
        RECT 64.410 143.780 64.580 144.770 ;
        RECT 64.760 144.600 64.930 145.120 ;
        RECT 65.110 144.950 65.280 145.650 ;
        RECT 65.580 145.500 65.750 146.090 ;
        RECT 65.930 146.130 66.880 146.160 ;
        RECT 65.930 145.960 65.960 146.130 ;
        RECT 66.130 145.960 66.320 146.130 ;
        RECT 66.490 145.960 66.680 146.130 ;
        RECT 66.850 145.960 66.880 146.130 ;
        RECT 65.930 145.680 66.880 145.960 ;
        RECT 67.060 146.090 68.090 146.260 ;
        RECT 67.060 145.500 67.230 146.090 ;
        RECT 65.580 145.450 67.230 145.500 ;
        RECT 65.460 145.330 67.230 145.450 ;
        RECT 65.460 145.130 65.790 145.330 ;
        RECT 67.410 145.150 67.740 145.910 ;
        RECT 67.920 145.730 68.090 146.090 ;
        RECT 68.270 146.130 69.220 146.210 ;
        RECT 68.270 145.960 68.300 146.130 ;
        RECT 68.470 145.960 68.660 146.130 ;
        RECT 68.830 145.960 69.020 146.130 ;
        RECT 69.190 145.960 69.220 146.130 ;
        RECT 68.270 145.910 69.220 145.960 ;
        RECT 67.920 145.560 69.730 145.730 ;
        RECT 65.970 144.980 67.740 145.150 ;
        RECT 65.970 144.950 66.140 144.980 ;
        RECT 65.110 144.780 66.140 144.950 ;
        RECT 69.050 144.800 69.380 145.380 ;
        RECT 64.760 144.370 65.790 144.600 ;
        RECT 65.460 143.880 65.790 144.370 ;
        RECT 65.970 144.100 66.140 144.780 ;
        RECT 66.320 144.630 69.380 144.800 ;
        RECT 66.320 144.280 66.650 144.630 ;
      LAYER li1 ;
        RECT 67.090 144.280 68.940 144.450 ;
      LAYER li1 ;
        RECT 65.970 143.930 68.590 144.100 ;
        RECT 64.410 143.280 64.680 143.780 ;
        RECT 65.970 143.700 66.140 143.930 ;
      LAYER li1 ;
        RECT 68.770 143.750 68.940 144.280 ;
      LAYER li1 ;
        RECT 65.130 143.530 66.140 143.700 ;
      LAYER li1 ;
        RECT 66.320 143.580 68.940 143.750 ;
      LAYER li1 ;
        RECT 65.130 143.280 65.460 143.530 ;
      LAYER li1 ;
        RECT 66.320 143.080 66.490 143.580 ;
        RECT 63.550 142.910 66.490 143.080 ;
      LAYER li1 ;
        RECT 67.640 142.820 68.590 143.400 ;
      LAYER li1 ;
        RECT 68.770 142.890 68.940 143.580 ;
      LAYER li1 ;
        RECT 69.120 143.780 69.380 144.630 ;
        RECT 69.560 144.210 69.730 145.560 ;
        RECT 69.910 145.300 70.160 146.210 ;
        RECT 70.970 146.130 71.920 146.160 ;
        RECT 72.750 146.130 73.650 146.160 ;
        RECT 70.970 145.960 71.000 146.130 ;
        RECT 71.170 145.960 71.360 146.130 ;
        RECT 71.530 145.960 71.720 146.130 ;
        RECT 71.890 145.960 71.920 146.130 ;
        RECT 72.920 145.960 73.110 146.130 ;
        RECT 73.280 145.960 73.470 146.130 ;
        RECT 73.640 145.960 73.650 146.130 ;
        RECT 69.910 145.130 70.790 145.300 ;
        RECT 70.970 145.130 71.920 145.960 ;
        RECT 72.320 145.160 72.570 145.630 ;
        RECT 72.750 145.340 73.650 145.960 ;
        RECT 74.260 146.130 75.200 146.190 ;
        RECT 74.260 145.960 74.280 146.130 ;
        RECT 74.450 145.960 74.640 146.130 ;
        RECT 74.810 145.960 75.000 146.130 ;
        RECT 75.170 145.960 75.200 146.130 ;
        RECT 70.110 144.390 70.440 144.890 ;
        RECT 70.620 144.810 70.790 145.130 ;
        RECT 72.320 144.990 73.330 145.160 ;
        RECT 70.620 144.640 72.980 144.810 ;
        RECT 69.560 144.040 70.730 144.210 ;
        RECT 69.120 143.070 69.450 143.780 ;
        RECT 69.910 143.240 70.240 143.780 ;
        RECT 70.450 143.540 70.730 144.040 ;
        RECT 70.910 143.240 71.080 144.640 ;
        RECT 73.160 144.460 73.330 144.990 ;
        RECT 71.290 144.290 73.330 144.460 ;
        RECT 71.290 143.900 71.620 144.290 ;
      LAYER li1 ;
        RECT 71.940 143.830 72.270 144.110 ;
        RECT 71.940 143.720 72.320 143.830 ;
      LAYER li1 ;
        RECT 69.910 143.070 71.080 143.240 ;
      LAYER li1 ;
        RECT 71.260 143.660 72.320 143.720 ;
        RECT 71.260 143.550 72.270 143.660 ;
        RECT 71.260 142.890 71.430 143.550 ;
      LAYER li1 ;
        RECT 73.100 143.450 73.330 144.290 ;
        RECT 73.830 144.460 74.080 145.460 ;
        RECT 74.260 144.650 75.200 145.960 ;
        RECT 76.090 146.180 77.540 146.210 ;
        RECT 76.090 146.010 76.340 146.180 ;
        RECT 76.510 146.010 76.700 146.180 ;
        RECT 76.870 146.010 77.140 146.180 ;
        RECT 77.310 146.010 77.540 146.180 ;
        RECT 76.090 145.140 77.540 146.010 ;
        RECT 77.850 146.130 78.800 146.210 ;
        RECT 77.850 145.960 77.880 146.130 ;
        RECT 78.050 145.960 78.240 146.130 ;
        RECT 78.410 145.960 78.600 146.130 ;
        RECT 78.770 145.960 78.800 146.130 ;
        RECT 73.830 144.130 75.200 144.460 ;
        RECT 73.830 143.950 74.040 144.130 ;
        RECT 73.710 143.450 74.040 143.950 ;
      LAYER li1 ;
        RECT 68.770 142.720 71.430 142.890 ;
      LAYER li1 ;
        RECT 71.610 142.820 72.560 143.370 ;
        RECT 73.100 142.950 73.430 143.450 ;
        RECT 74.220 142.820 75.170 143.950 ;
        RECT 76.320 143.700 76.650 144.480 ;
        RECT 76.860 144.150 77.190 145.140 ;
        RECT 77.850 144.630 78.800 145.960 ;
      LAYER li1 ;
        RECT 78.980 144.530 79.230 146.210 ;
      LAYER li1 ;
        RECT 79.410 146.130 80.360 146.210 ;
        RECT 79.410 145.960 79.440 146.130 ;
        RECT 79.610 145.960 79.800 146.130 ;
        RECT 79.970 145.960 80.160 146.130 ;
        RECT 80.330 145.960 80.360 146.130 ;
        RECT 79.410 144.710 80.360 145.960 ;
      LAYER li1 ;
        RECT 80.540 144.530 80.870 146.210 ;
      LAYER li1 ;
        RECT 81.050 146.130 82.000 146.210 ;
        RECT 81.050 145.960 81.080 146.130 ;
        RECT 81.250 145.960 81.440 146.130 ;
        RECT 81.610 145.960 81.800 146.130 ;
        RECT 81.970 145.960 82.000 146.130 ;
        RECT 81.050 144.750 82.000 145.960 ;
      LAYER li1 ;
        RECT 78.980 144.360 80.870 144.530 ;
        RECT 78.980 144.230 79.150 144.360 ;
        RECT 77.890 144.000 79.150 144.230 ;
      LAYER li1 ;
        RECT 79.330 144.050 81.360 144.180 ;
        RECT 82.180 144.050 82.430 146.210 ;
        RECT 82.810 146.180 84.260 146.210 ;
        RECT 82.810 146.010 83.060 146.180 ;
        RECT 83.230 146.010 83.420 146.180 ;
        RECT 83.590 146.010 83.860 146.180 ;
        RECT 84.030 146.010 84.260 146.180 ;
        RECT 82.810 145.140 84.260 146.010 ;
        RECT 79.330 144.010 82.430 144.050 ;
      LAYER li1 ;
        RECT 78.980 143.830 79.150 144.000 ;
      LAYER li1 ;
        RECT 81.190 143.880 82.430 144.010 ;
        RECT 76.320 143.300 77.620 143.700 ;
        RECT 76.010 142.820 77.620 143.300 ;
        RECT 77.850 142.820 78.800 143.780 ;
      LAYER li1 ;
        RECT 78.980 143.660 80.790 143.830 ;
        RECT 78.980 142.950 79.230 143.660 ;
      LAYER li1 ;
        RECT 79.410 142.820 80.360 143.480 ;
      LAYER li1 ;
        RECT 80.540 142.950 80.790 143.660 ;
      LAYER li1 ;
        RECT 80.970 142.820 81.920 143.700 ;
        RECT 82.100 142.950 82.430 143.880 ;
        RECT 83.040 143.700 83.370 144.480 ;
        RECT 83.580 144.150 83.910 145.140 ;
      LAYER li1 ;
        RECT 86.040 144.630 86.470 146.210 ;
      LAYER li1 ;
        RECT 86.650 146.130 87.210 146.210 ;
        RECT 86.650 145.960 86.660 146.130 ;
        RECT 86.830 145.960 87.020 146.130 ;
        RECT 87.190 145.960 87.210 146.130 ;
        RECT 86.650 144.630 87.210 145.960 ;
        RECT 88.820 146.180 91.560 146.200 ;
        RECT 88.820 146.010 89.030 146.180 ;
        RECT 89.200 146.010 89.470 146.180 ;
        RECT 89.640 146.010 89.880 146.180 ;
        RECT 90.050 146.010 90.310 146.180 ;
        RECT 90.480 146.010 90.750 146.180 ;
        RECT 90.920 146.010 91.160 146.180 ;
        RECT 91.330 146.010 91.560 146.180 ;
        RECT 83.040 143.300 84.340 143.700 ;
        RECT 82.730 142.820 84.340 143.300 ;
      LAYER li1 ;
        RECT 86.040 142.950 86.290 144.630 ;
      LAYER li1 ;
        RECT 86.600 143.740 86.930 144.200 ;
      LAYER li1 ;
        RECT 87.390 143.920 87.720 145.710 ;
      LAYER li1 ;
        RECT 87.900 143.740 88.150 145.460 ;
        RECT 88.820 145.130 91.560 146.010 ;
        RECT 92.660 146.180 95.400 146.200 ;
        RECT 92.660 146.010 92.870 146.180 ;
        RECT 93.040 146.010 93.310 146.180 ;
        RECT 93.480 146.010 93.720 146.180 ;
        RECT 93.890 146.010 94.150 146.180 ;
        RECT 94.320 146.010 94.590 146.180 ;
        RECT 94.760 146.010 95.000 146.180 ;
        RECT 95.170 146.010 95.400 146.180 ;
        RECT 92.660 145.130 95.400 146.010 ;
        RECT 96.250 146.180 97.700 146.210 ;
        RECT 96.250 146.010 96.500 146.180 ;
        RECT 96.670 146.010 96.860 146.180 ;
        RECT 97.030 146.010 97.300 146.180 ;
        RECT 97.470 146.010 97.700 146.180 ;
        RECT 96.250 145.140 97.700 146.010 ;
        RECT 89.060 143.810 89.390 144.480 ;
        RECT 89.790 144.150 90.120 145.130 ;
        RECT 90.340 143.810 90.670 144.480 ;
        RECT 91.070 144.150 91.400 145.130 ;
        RECT 92.900 143.810 93.230 144.480 ;
        RECT 93.630 144.150 93.960 145.130 ;
        RECT 94.180 143.810 94.510 144.480 ;
        RECT 94.910 144.150 95.240 145.130 ;
        RECT 86.600 143.570 88.150 143.740 ;
        RECT 86.470 142.820 87.720 143.390 ;
        RECT 87.900 142.950 88.150 143.570 ;
        RECT 88.900 142.810 91.630 143.810 ;
        RECT 92.740 142.810 95.470 143.810 ;
        RECT 96.480 143.700 96.810 144.480 ;
        RECT 97.020 144.150 97.350 145.140 ;
      LAYER li1 ;
        RECT 98.040 144.630 98.470 146.210 ;
      LAYER li1 ;
        RECT 98.650 146.130 99.210 146.210 ;
        RECT 98.650 145.960 98.660 146.130 ;
        RECT 98.830 145.960 99.020 146.130 ;
        RECT 99.190 145.960 99.210 146.130 ;
        RECT 98.650 144.630 99.210 145.960 ;
        RECT 100.570 146.180 102.020 146.210 ;
        RECT 100.570 146.010 100.820 146.180 ;
        RECT 100.990 146.010 101.180 146.180 ;
        RECT 101.350 146.010 101.620 146.180 ;
        RECT 101.790 146.010 102.020 146.180 ;
        RECT 96.480 143.300 97.780 143.700 ;
        RECT 96.170 142.820 97.780 143.300 ;
      LAYER li1 ;
        RECT 98.040 142.950 98.290 144.630 ;
      LAYER li1 ;
        RECT 98.600 143.740 98.930 144.200 ;
      LAYER li1 ;
        RECT 99.390 143.920 99.720 145.710 ;
      LAYER li1 ;
        RECT 99.900 143.740 100.150 145.460 ;
        RECT 100.570 145.140 102.020 146.010 ;
        RECT 102.970 146.130 103.530 146.210 ;
        RECT 102.970 145.960 102.980 146.130 ;
        RECT 103.150 145.960 103.340 146.130 ;
        RECT 103.510 145.960 103.530 146.130 ;
        RECT 98.600 143.570 100.150 143.740 ;
        RECT 98.470 142.820 99.720 143.390 ;
        RECT 99.900 142.950 100.150 143.570 ;
        RECT 100.800 143.700 101.130 144.480 ;
        RECT 101.340 144.150 101.670 145.140 ;
        RECT 102.970 144.630 103.530 145.960 ;
        RECT 104.890 146.180 106.340 146.210 ;
        RECT 104.890 146.010 105.140 146.180 ;
        RECT 105.310 146.010 105.500 146.180 ;
        RECT 105.670 146.010 105.940 146.180 ;
        RECT 106.110 146.010 106.340 146.180 ;
        RECT 102.920 143.740 103.250 144.200 ;
        RECT 104.220 143.740 104.470 145.460 ;
        RECT 104.890 145.140 106.340 146.010 ;
        RECT 100.800 143.300 102.100 143.700 ;
        RECT 102.920 143.570 104.470 143.740 ;
        RECT 100.490 142.820 102.100 143.300 ;
        RECT 102.790 142.820 104.040 143.390 ;
        RECT 104.220 142.950 104.470 143.570 ;
        RECT 105.120 143.700 105.450 144.480 ;
        RECT 105.660 144.150 105.990 145.140 ;
      LAYER li1 ;
        RECT 106.680 144.630 107.110 146.210 ;
      LAYER li1 ;
        RECT 107.290 146.130 107.850 146.210 ;
        RECT 107.290 145.960 107.300 146.130 ;
        RECT 107.470 145.960 107.660 146.130 ;
        RECT 107.830 145.960 107.850 146.130 ;
        RECT 107.290 144.630 107.850 145.960 ;
        RECT 109.460 146.180 112.200 146.200 ;
        RECT 109.460 146.010 109.670 146.180 ;
        RECT 109.840 146.010 110.110 146.180 ;
        RECT 110.280 146.010 110.520 146.180 ;
        RECT 110.690 146.010 110.950 146.180 ;
        RECT 111.120 146.010 111.390 146.180 ;
        RECT 111.560 146.010 111.800 146.180 ;
        RECT 111.970 146.010 112.200 146.180 ;
        RECT 105.120 143.300 106.420 143.700 ;
        RECT 104.810 142.820 106.420 143.300 ;
      LAYER li1 ;
        RECT 106.680 142.950 106.930 144.630 ;
      LAYER li1 ;
        RECT 107.240 143.740 107.570 144.200 ;
      LAYER li1 ;
        RECT 108.030 143.920 108.360 145.710 ;
      LAYER li1 ;
        RECT 108.540 143.740 108.790 145.460 ;
        RECT 109.460 145.130 112.200 146.010 ;
        RECT 113.300 146.180 116.040 146.200 ;
        RECT 113.300 146.010 113.510 146.180 ;
        RECT 113.680 146.010 113.950 146.180 ;
        RECT 114.120 146.010 114.360 146.180 ;
        RECT 114.530 146.010 114.790 146.180 ;
        RECT 114.960 146.010 115.230 146.180 ;
        RECT 115.400 146.010 115.640 146.180 ;
        RECT 115.810 146.010 116.040 146.180 ;
        RECT 113.300 145.130 116.040 146.010 ;
        RECT 117.140 146.180 119.880 146.200 ;
        RECT 117.140 146.010 117.350 146.180 ;
        RECT 117.520 146.010 117.790 146.180 ;
        RECT 117.960 146.010 118.200 146.180 ;
        RECT 118.370 146.010 118.630 146.180 ;
        RECT 118.800 146.010 119.070 146.180 ;
        RECT 119.240 146.010 119.480 146.180 ;
        RECT 119.650 146.010 119.880 146.180 ;
        RECT 117.140 145.130 119.880 146.010 ;
        RECT 120.980 146.180 123.720 146.200 ;
        RECT 120.980 146.010 121.190 146.180 ;
        RECT 121.360 146.010 121.630 146.180 ;
        RECT 121.800 146.010 122.040 146.180 ;
        RECT 122.210 146.010 122.470 146.180 ;
        RECT 122.640 146.010 122.910 146.180 ;
        RECT 123.080 146.010 123.320 146.180 ;
        RECT 123.490 146.010 123.720 146.180 ;
        RECT 120.980 145.130 123.720 146.010 ;
        RECT 124.570 146.180 126.020 146.210 ;
        RECT 124.570 146.010 124.820 146.180 ;
        RECT 124.990 146.010 125.180 146.180 ;
        RECT 125.350 146.010 125.620 146.180 ;
        RECT 125.790 146.010 126.020 146.180 ;
        RECT 124.570 145.140 126.020 146.010 ;
        RECT 127.420 146.130 128.070 146.240 ;
        RECT 127.420 145.960 127.480 146.130 ;
        RECT 127.650 145.960 127.840 146.130 ;
        RECT 128.010 145.960 128.070 146.130 ;
        RECT 130.100 146.180 132.840 146.200 ;
        RECT 130.100 146.010 130.310 146.180 ;
        RECT 130.480 146.010 130.750 146.180 ;
        RECT 130.920 146.010 131.160 146.180 ;
        RECT 131.330 146.010 131.590 146.180 ;
        RECT 131.760 146.010 132.030 146.180 ;
        RECT 132.200 146.010 132.440 146.180 ;
        RECT 132.610 146.010 132.840 146.180 ;
        RECT 127.420 145.900 128.070 145.960 ;
        RECT 127.420 145.630 127.820 145.900 ;
        RECT 109.700 143.810 110.030 144.480 ;
        RECT 110.430 144.150 110.760 145.130 ;
        RECT 110.980 143.810 111.310 144.480 ;
        RECT 111.710 144.150 112.040 145.130 ;
        RECT 113.540 143.810 113.870 144.480 ;
        RECT 114.270 144.150 114.600 145.130 ;
        RECT 114.820 143.810 115.150 144.480 ;
        RECT 115.550 144.150 115.880 145.130 ;
        RECT 117.380 143.810 117.710 144.480 ;
        RECT 118.110 144.150 118.440 145.130 ;
        RECT 118.660 143.810 118.990 144.480 ;
        RECT 119.390 144.150 119.720 145.130 ;
        RECT 121.220 143.810 121.550 144.480 ;
        RECT 121.950 144.150 122.280 145.130 ;
        RECT 122.500 143.810 122.830 144.480 ;
        RECT 123.230 144.150 123.560 145.130 ;
        RECT 107.240 143.570 108.790 143.740 ;
        RECT 107.110 142.820 108.360 143.390 ;
        RECT 108.540 142.950 108.790 143.570 ;
        RECT 109.540 142.810 112.270 143.810 ;
        RECT 113.380 142.810 116.110 143.810 ;
        RECT 117.220 142.810 119.950 143.810 ;
        RECT 121.060 142.810 123.790 143.810 ;
        RECT 124.800 143.700 125.130 144.480 ;
        RECT 125.340 144.150 125.670 145.140 ;
      LAYER li1 ;
        RECT 128.280 144.640 128.530 145.980 ;
      LAYER li1 ;
        RECT 130.100 145.130 132.840 146.010 ;
        RECT 134.170 146.130 134.730 146.210 ;
        RECT 134.170 145.960 134.180 146.130 ;
        RECT 134.350 145.960 134.540 146.130 ;
        RECT 134.710 145.960 134.730 146.130 ;
      LAYER li1 ;
        RECT 127.820 144.390 128.530 144.640 ;
      LAYER li1 ;
        RECT 124.800 143.300 126.100 143.700 ;
      LAYER li1 ;
        RECT 127.820 143.520 128.070 144.390 ;
      LAYER li1 ;
        RECT 130.340 143.810 130.670 144.480 ;
        RECT 131.070 144.150 131.400 145.130 ;
        RECT 131.620 143.810 131.950 144.480 ;
        RECT 132.350 144.150 132.680 145.130 ;
        RECT 134.170 144.630 134.730 145.960 ;
        RECT 136.340 146.180 139.080 146.200 ;
        RECT 136.340 146.010 136.550 146.180 ;
        RECT 136.720 146.010 136.990 146.180 ;
        RECT 137.160 146.010 137.400 146.180 ;
        RECT 137.570 146.010 137.830 146.180 ;
        RECT 138.000 146.010 138.270 146.180 ;
        RECT 138.440 146.010 138.680 146.180 ;
        RECT 138.850 146.010 139.080 146.180 ;
        RECT 124.490 142.820 126.100 143.300 ;
      LAYER li1 ;
        RECT 127.490 142.880 128.070 143.520 ;
      LAYER li1 ;
        RECT 128.980 143.080 129.390 143.520 ;
        RECT 128.740 142.740 129.390 143.080 ;
        RECT 130.180 142.810 132.910 143.810 ;
        RECT 134.120 143.740 134.450 144.200 ;
        RECT 135.420 143.740 135.670 145.460 ;
        RECT 136.340 145.130 139.080 146.010 ;
        RECT 139.930 146.180 141.380 146.210 ;
        RECT 139.930 146.010 140.180 146.180 ;
        RECT 140.350 146.010 140.540 146.180 ;
        RECT 140.710 146.010 140.980 146.180 ;
        RECT 141.150 146.010 141.380 146.180 ;
        RECT 139.930 145.140 141.380 146.010 ;
        RECT 136.580 143.810 136.910 144.480 ;
        RECT 137.310 144.150 137.640 145.130 ;
        RECT 137.860 143.810 138.190 144.480 ;
        RECT 138.590 144.150 138.920 145.130 ;
        RECT 134.120 143.570 135.670 143.740 ;
        RECT 133.990 142.820 135.240 143.390 ;
        RECT 135.420 142.950 135.670 143.570 ;
        RECT 136.420 142.810 139.150 143.810 ;
        RECT 140.160 143.700 140.490 144.480 ;
        RECT 140.700 144.150 141.030 145.140 ;
        RECT 140.160 143.300 141.460 143.700 ;
        RECT 139.850 142.820 141.460 143.300 ;
        RECT 5.760 142.360 5.920 142.540 ;
        RECT 6.090 142.360 6.400 142.540 ;
        RECT 6.570 142.360 6.880 142.540 ;
        RECT 7.050 142.360 7.360 142.540 ;
        RECT 7.530 142.360 7.840 142.540 ;
        RECT 8.010 142.360 8.320 142.540 ;
        RECT 8.490 142.360 8.800 142.540 ;
        RECT 8.970 142.360 9.280 142.540 ;
        RECT 9.450 142.360 9.760 142.540 ;
        RECT 9.930 142.360 10.240 142.540 ;
        RECT 10.410 142.360 10.720 142.540 ;
        RECT 10.890 142.360 11.200 142.540 ;
        RECT 11.370 142.360 11.680 142.540 ;
        RECT 11.850 142.360 12.160 142.540 ;
        RECT 12.330 142.360 12.640 142.540 ;
        RECT 12.810 142.360 13.120 142.540 ;
        RECT 13.290 142.360 13.600 142.540 ;
        RECT 13.770 142.360 14.080 142.540 ;
        RECT 14.250 142.360 14.560 142.540 ;
        RECT 14.730 142.360 15.040 142.540 ;
        RECT 15.210 142.360 15.520 142.540 ;
        RECT 15.690 142.360 16.000 142.540 ;
        RECT 16.170 142.360 16.480 142.540 ;
        RECT 16.650 142.360 16.960 142.540 ;
        RECT 17.130 142.360 17.440 142.540 ;
        RECT 17.610 142.360 17.760 142.540 ;
        RECT 18.240 142.360 18.400 142.540 ;
        RECT 18.570 142.360 18.880 142.540 ;
        RECT 19.050 142.360 19.360 142.540 ;
        RECT 19.530 142.360 19.840 142.540 ;
        RECT 20.010 142.360 20.320 142.540 ;
        RECT 20.490 142.360 20.800 142.540 ;
        RECT 20.970 142.360 21.280 142.540 ;
        RECT 21.450 142.360 21.760 142.540 ;
        RECT 21.930 142.360 22.240 142.540 ;
        RECT 22.410 142.360 22.720 142.540 ;
        RECT 22.890 142.360 23.200 142.540 ;
        RECT 23.370 142.360 23.680 142.540 ;
        RECT 23.850 142.360 24.160 142.540 ;
        RECT 24.330 142.360 24.640 142.540 ;
        RECT 24.810 142.360 25.120 142.540 ;
        RECT 25.290 142.360 25.600 142.540 ;
        RECT 25.770 142.360 26.080 142.540 ;
        RECT 26.250 142.360 26.560 142.540 ;
        RECT 26.730 142.360 27.040 142.540 ;
        RECT 27.210 142.360 27.520 142.540 ;
        RECT 27.690 142.360 28.000 142.540 ;
        RECT 28.170 142.360 28.480 142.540 ;
        RECT 28.650 142.360 28.960 142.540 ;
        RECT 29.130 142.360 29.440 142.540 ;
        RECT 29.610 142.360 29.920 142.540 ;
        RECT 30.090 142.360 30.400 142.540 ;
        RECT 30.570 142.360 30.880 142.540 ;
        RECT 31.050 142.360 31.360 142.540 ;
        RECT 31.530 142.360 31.840 142.540 ;
        RECT 32.010 142.360 32.320 142.540 ;
        RECT 32.490 142.360 32.800 142.540 ;
        RECT 32.970 142.360 33.280 142.540 ;
        RECT 33.450 142.360 33.760 142.540 ;
        RECT 33.930 142.360 34.240 142.540 ;
        RECT 34.410 142.360 34.720 142.540 ;
        RECT 34.890 142.360 35.200 142.540 ;
        RECT 35.370 142.360 35.680 142.540 ;
        RECT 35.850 142.360 36.000 142.540 ;
        RECT 36.480 142.360 36.640 142.540 ;
        RECT 36.810 142.360 37.120 142.540 ;
        RECT 37.290 142.360 37.600 142.540 ;
        RECT 37.770 142.360 38.080 142.540 ;
        RECT 38.250 142.360 38.560 142.540 ;
        RECT 38.730 142.360 39.040 142.540 ;
        RECT 39.210 142.360 39.520 142.540 ;
        RECT 39.690 142.360 40.000 142.540 ;
        RECT 40.170 142.360 40.480 142.540 ;
        RECT 40.650 142.360 40.960 142.540 ;
        RECT 41.130 142.360 41.440 142.540 ;
        RECT 41.610 142.360 41.920 142.540 ;
        RECT 42.090 142.360 42.400 142.540 ;
        RECT 42.570 142.360 42.880 142.540 ;
        RECT 43.050 142.360 43.360 142.540 ;
        RECT 43.530 142.360 43.680 142.540 ;
        RECT 44.160 142.360 44.320 142.540 ;
        RECT 44.490 142.360 44.800 142.540 ;
        RECT 44.970 142.360 45.280 142.540 ;
        RECT 45.450 142.360 45.760 142.540 ;
        RECT 45.930 142.360 46.240 142.540 ;
        RECT 46.410 142.360 46.720 142.540 ;
        RECT 46.890 142.360 47.200 142.540 ;
        RECT 47.370 142.360 47.680 142.540 ;
        RECT 47.850 142.360 48.160 142.540 ;
        RECT 48.330 142.360 48.640 142.540 ;
        RECT 48.810 142.360 49.120 142.540 ;
        RECT 49.290 142.360 49.600 142.540 ;
        RECT 49.770 142.360 50.080 142.540 ;
        RECT 50.250 142.360 50.560 142.540 ;
        RECT 50.730 142.360 51.040 142.540 ;
        RECT 51.210 142.360 51.520 142.540 ;
        RECT 51.690 142.360 52.000 142.540 ;
        RECT 52.170 142.360 52.480 142.540 ;
        RECT 52.650 142.360 52.960 142.540 ;
        RECT 53.130 142.360 53.440 142.540 ;
        RECT 53.610 142.360 53.920 142.540 ;
        RECT 54.090 142.360 54.400 142.540 ;
        RECT 54.570 142.360 54.880 142.540 ;
        RECT 55.050 142.360 55.360 142.540 ;
        RECT 55.530 142.360 55.840 142.540 ;
        RECT 56.010 142.360 56.320 142.540 ;
        RECT 56.490 142.360 56.800 142.540 ;
        RECT 56.970 142.360 57.280 142.540 ;
        RECT 57.450 142.360 57.760 142.540 ;
        RECT 57.930 142.360 58.240 142.540 ;
        RECT 58.410 142.360 58.720 142.540 ;
        RECT 58.890 142.360 59.200 142.540 ;
        RECT 59.370 142.360 59.680 142.540 ;
        RECT 59.850 142.360 60.160 142.540 ;
        RECT 60.330 142.360 60.640 142.540 ;
        RECT 60.810 142.360 61.120 142.540 ;
        RECT 61.290 142.360 61.600 142.540 ;
        RECT 61.770 142.360 62.080 142.540 ;
        RECT 62.250 142.360 62.560 142.540 ;
        RECT 62.730 142.360 63.040 142.540 ;
        RECT 63.210 142.360 63.520 142.540 ;
        RECT 63.690 142.360 64.000 142.540 ;
        RECT 64.170 142.360 64.480 142.540 ;
        RECT 64.650 142.360 64.960 142.540 ;
        RECT 65.130 142.360 65.440 142.540 ;
        RECT 65.610 142.360 65.920 142.540 ;
        RECT 66.090 142.360 66.400 142.540 ;
        RECT 66.570 142.360 66.880 142.540 ;
        RECT 67.050 142.360 67.360 142.540 ;
        RECT 67.530 142.360 67.840 142.540 ;
        RECT 68.010 142.360 68.320 142.540 ;
        RECT 68.490 142.360 68.800 142.540 ;
        RECT 68.970 142.360 69.280 142.540 ;
        RECT 69.450 142.360 69.760 142.540 ;
        RECT 69.930 142.360 70.240 142.540 ;
        RECT 70.410 142.360 70.720 142.540 ;
        RECT 70.890 142.360 71.200 142.540 ;
        RECT 71.370 142.360 71.680 142.540 ;
        RECT 71.850 142.360 72.160 142.540 ;
        RECT 72.330 142.360 72.640 142.540 ;
        RECT 72.810 142.360 73.120 142.540 ;
        RECT 73.290 142.360 73.600 142.540 ;
        RECT 73.770 142.360 74.080 142.540 ;
        RECT 74.250 142.360 74.560 142.540 ;
        RECT 74.730 142.360 75.040 142.540 ;
        RECT 75.210 142.360 75.520 142.540 ;
        RECT 75.690 142.360 76.000 142.540 ;
        RECT 76.170 142.360 76.480 142.540 ;
        RECT 76.650 142.360 76.960 142.540 ;
        RECT 77.130 142.360 77.440 142.540 ;
        RECT 77.610 142.360 77.920 142.540 ;
        RECT 78.090 142.360 78.400 142.540 ;
        RECT 78.570 142.360 78.880 142.540 ;
        RECT 79.050 142.360 79.360 142.540 ;
        RECT 79.530 142.360 79.840 142.540 ;
        RECT 80.010 142.360 80.320 142.540 ;
        RECT 80.490 142.360 80.800 142.540 ;
        RECT 80.970 142.360 81.280 142.540 ;
        RECT 81.450 142.360 81.760 142.540 ;
        RECT 81.930 142.360 82.240 142.540 ;
        RECT 82.410 142.360 82.720 142.540 ;
        RECT 82.890 142.360 83.200 142.540 ;
        RECT 83.370 142.360 83.680 142.540 ;
        RECT 83.850 142.360 84.160 142.540 ;
        RECT 84.330 142.360 84.640 142.540 ;
        RECT 84.810 142.360 85.120 142.540 ;
        RECT 85.290 142.360 85.440 142.540 ;
        RECT 85.920 142.360 86.080 142.540 ;
        RECT 86.250 142.360 86.560 142.540 ;
        RECT 86.730 142.360 87.040 142.540 ;
        RECT 87.210 142.360 87.520 142.540 ;
        RECT 87.690 142.360 88.000 142.540 ;
        RECT 88.170 142.360 88.480 142.540 ;
        RECT 88.650 142.360 88.960 142.540 ;
        RECT 89.130 142.360 89.440 142.540 ;
        RECT 89.610 142.360 89.920 142.540 ;
        RECT 90.090 142.360 90.400 142.540 ;
        RECT 90.570 142.360 90.880 142.540 ;
        RECT 91.050 142.360 91.360 142.540 ;
        RECT 91.530 142.360 91.840 142.540 ;
        RECT 92.010 142.360 92.320 142.540 ;
        RECT 92.490 142.360 92.800 142.540 ;
        RECT 92.970 142.360 93.280 142.540 ;
        RECT 93.450 142.360 93.760 142.540 ;
        RECT 93.930 142.360 94.240 142.540 ;
        RECT 94.410 142.360 94.720 142.540 ;
        RECT 94.890 142.360 95.200 142.540 ;
        RECT 95.370 142.360 95.680 142.540 ;
        RECT 95.850 142.360 96.160 142.540 ;
        RECT 96.330 142.360 96.640 142.540 ;
        RECT 96.810 142.360 97.120 142.540 ;
        RECT 97.290 142.360 97.600 142.540 ;
        RECT 97.770 142.360 98.080 142.540 ;
        RECT 98.250 142.360 98.560 142.540 ;
        RECT 98.730 142.360 99.040 142.540 ;
        RECT 99.210 142.360 99.520 142.540 ;
        RECT 99.690 142.360 100.000 142.540 ;
        RECT 100.170 142.360 100.480 142.540 ;
        RECT 100.650 142.360 100.960 142.540 ;
        RECT 101.130 142.360 101.440 142.540 ;
        RECT 101.610 142.360 101.920 142.540 ;
        RECT 102.090 142.360 102.400 142.540 ;
        RECT 102.570 142.360 102.880 142.540 ;
        RECT 103.050 142.360 103.360 142.540 ;
        RECT 103.530 142.360 103.840 142.540 ;
        RECT 104.010 142.360 104.320 142.540 ;
        RECT 104.490 142.360 104.800 142.540 ;
        RECT 104.970 142.360 105.280 142.540 ;
        RECT 105.450 142.360 105.760 142.540 ;
        RECT 105.930 142.360 106.240 142.540 ;
        RECT 106.410 142.360 106.720 142.540 ;
        RECT 106.890 142.360 107.200 142.540 ;
        RECT 107.370 142.360 107.680 142.540 ;
        RECT 107.850 142.360 108.160 142.540 ;
        RECT 108.330 142.360 108.640 142.540 ;
        RECT 108.810 142.360 109.120 142.540 ;
        RECT 109.290 142.360 109.600 142.540 ;
        RECT 109.770 142.360 110.080 142.540 ;
        RECT 110.250 142.360 110.560 142.540 ;
        RECT 110.730 142.360 111.040 142.540 ;
        RECT 111.210 142.360 111.520 142.540 ;
        RECT 111.690 142.360 112.000 142.540 ;
        RECT 112.170 142.360 112.480 142.540 ;
        RECT 112.650 142.360 112.960 142.540 ;
        RECT 113.130 142.360 113.440 142.540 ;
        RECT 113.610 142.360 113.920 142.540 ;
        RECT 114.090 142.360 114.400 142.540 ;
        RECT 114.570 142.360 114.880 142.540 ;
        RECT 115.050 142.360 115.360 142.540 ;
        RECT 115.530 142.360 115.840 142.540 ;
        RECT 116.010 142.360 116.320 142.540 ;
        RECT 116.490 142.360 116.800 142.540 ;
        RECT 116.970 142.360 117.280 142.540 ;
        RECT 117.450 142.360 117.760 142.540 ;
        RECT 117.930 142.360 118.240 142.540 ;
        RECT 118.410 142.360 118.720 142.540 ;
        RECT 118.890 142.360 119.200 142.540 ;
        RECT 119.370 142.360 119.680 142.540 ;
        RECT 119.850 142.360 120.160 142.540 ;
        RECT 120.330 142.360 120.640 142.540 ;
        RECT 120.810 142.360 121.120 142.540 ;
        RECT 121.290 142.360 121.600 142.540 ;
        RECT 121.770 142.360 122.080 142.540 ;
        RECT 122.250 142.360 122.560 142.540 ;
        RECT 122.730 142.360 123.040 142.540 ;
        RECT 123.210 142.360 123.520 142.540 ;
        RECT 123.690 142.360 124.000 142.540 ;
        RECT 124.170 142.360 124.480 142.540 ;
        RECT 124.650 142.360 124.960 142.540 ;
        RECT 125.130 142.360 125.440 142.540 ;
        RECT 125.610 142.360 125.920 142.540 ;
        RECT 126.090 142.360 126.400 142.540 ;
        RECT 126.570 142.360 126.880 142.540 ;
        RECT 127.050 142.360 127.360 142.540 ;
        RECT 127.530 142.360 127.840 142.540 ;
        RECT 128.010 142.360 128.320 142.540 ;
        RECT 128.490 142.360 128.800 142.540 ;
        RECT 128.970 142.360 129.280 142.540 ;
        RECT 129.450 142.360 129.760 142.540 ;
        RECT 129.930 142.360 130.240 142.540 ;
        RECT 130.410 142.360 130.720 142.540 ;
        RECT 130.890 142.360 131.200 142.540 ;
        RECT 131.370 142.360 131.680 142.540 ;
        RECT 131.850 142.360 132.160 142.540 ;
        RECT 132.330 142.360 132.640 142.540 ;
        RECT 132.810 142.360 133.120 142.540 ;
        RECT 133.290 142.360 133.600 142.540 ;
        RECT 133.770 142.360 134.080 142.540 ;
        RECT 134.250 142.360 134.560 142.540 ;
        RECT 134.730 142.360 135.040 142.540 ;
        RECT 135.210 142.360 135.520 142.540 ;
        RECT 135.690 142.360 136.000 142.540 ;
        RECT 136.170 142.360 136.480 142.540 ;
        RECT 136.650 142.360 136.960 142.540 ;
        RECT 137.130 142.360 137.440 142.540 ;
        RECT 137.610 142.360 137.920 142.540 ;
        RECT 138.090 142.360 138.400 142.540 ;
        RECT 138.570 142.360 138.880 142.540 ;
        RECT 139.050 142.360 139.360 142.540 ;
        RECT 139.530 142.360 139.840 142.540 ;
        RECT 140.010 142.360 140.320 142.540 ;
        RECT 140.490 142.360 140.800 142.540 ;
        RECT 140.970 142.360 141.280 142.540 ;
        RECT 141.450 142.360 141.600 142.540 ;
        RECT 6.340 142.060 9.070 142.090 ;
        RECT 6.340 141.890 6.510 142.060 ;
        RECT 6.680 141.890 6.950 142.060 ;
        RECT 7.120 141.890 7.360 142.060 ;
        RECT 7.530 141.890 7.790 142.060 ;
        RECT 7.960 141.890 8.230 142.060 ;
        RECT 8.400 141.890 8.640 142.060 ;
        RECT 8.810 141.890 9.070 142.060 ;
        RECT 6.340 141.090 9.070 141.890 ;
        RECT 10.180 142.060 12.910 142.090 ;
        RECT 10.180 141.890 10.350 142.060 ;
        RECT 10.520 141.890 10.790 142.060 ;
        RECT 10.960 141.890 11.200 142.060 ;
        RECT 11.370 141.890 11.630 142.060 ;
        RECT 11.800 141.890 12.070 142.060 ;
        RECT 12.240 141.890 12.480 142.060 ;
        RECT 12.650 141.890 12.910 142.060 ;
        RECT 10.180 141.090 12.910 141.890 ;
        RECT 14.020 142.060 16.750 142.090 ;
        RECT 14.020 141.890 14.190 142.060 ;
        RECT 14.360 141.890 14.630 142.060 ;
        RECT 14.800 141.890 15.040 142.060 ;
        RECT 15.210 141.890 15.470 142.060 ;
        RECT 15.640 141.890 15.910 142.060 ;
        RECT 16.080 141.890 16.320 142.060 ;
        RECT 16.490 141.890 16.750 142.060 ;
        RECT 14.020 141.090 16.750 141.890 ;
        RECT 17.860 142.060 20.590 142.090 ;
        RECT 17.860 141.890 18.030 142.060 ;
        RECT 18.200 141.890 18.470 142.060 ;
        RECT 18.640 141.890 18.880 142.060 ;
        RECT 19.050 141.890 19.310 142.060 ;
        RECT 19.480 141.890 19.750 142.060 ;
        RECT 19.920 141.890 20.160 142.060 ;
        RECT 20.330 141.890 20.590 142.060 ;
        RECT 17.860 141.090 20.590 141.890 ;
        RECT 21.700 142.060 24.430 142.090 ;
        RECT 21.700 141.890 21.870 142.060 ;
        RECT 22.040 141.890 22.310 142.060 ;
        RECT 22.480 141.890 22.720 142.060 ;
        RECT 22.890 141.890 23.150 142.060 ;
        RECT 23.320 141.890 23.590 142.060 ;
        RECT 23.760 141.890 24.000 142.060 ;
        RECT 24.170 141.890 24.430 142.060 ;
        RECT 21.700 141.090 24.430 141.890 ;
        RECT 25.540 142.060 28.270 142.090 ;
        RECT 25.540 141.890 25.710 142.060 ;
        RECT 25.880 141.890 26.150 142.060 ;
        RECT 26.320 141.890 26.560 142.060 ;
        RECT 26.730 141.890 26.990 142.060 ;
        RECT 27.160 141.890 27.430 142.060 ;
        RECT 27.600 141.890 27.840 142.060 ;
        RECT 28.010 141.890 28.270 142.060 ;
        RECT 30.800 142.050 31.750 142.080 ;
        RECT 25.540 141.090 28.270 141.890 ;
        RECT 6.500 140.420 6.830 141.090 ;
        RECT 7.230 139.770 7.560 140.750 ;
        RECT 7.780 140.420 8.110 141.090 ;
        RECT 8.510 139.770 8.840 140.750 ;
        RECT 10.340 140.420 10.670 141.090 ;
        RECT 11.070 139.770 11.400 140.750 ;
        RECT 11.620 140.420 11.950 141.090 ;
        RECT 12.350 139.770 12.680 140.750 ;
        RECT 14.180 140.420 14.510 141.090 ;
        RECT 14.910 139.770 15.240 140.750 ;
        RECT 15.460 140.420 15.790 141.090 ;
        RECT 16.190 139.770 16.520 140.750 ;
        RECT 18.020 140.420 18.350 141.090 ;
        RECT 18.750 139.770 19.080 140.750 ;
        RECT 19.300 140.420 19.630 141.090 ;
        RECT 20.030 139.770 20.360 140.750 ;
        RECT 21.860 140.420 22.190 141.090 ;
        RECT 22.590 139.770 22.920 140.750 ;
        RECT 23.140 140.420 23.470 141.090 ;
        RECT 23.870 139.770 24.200 140.750 ;
        RECT 25.700 140.420 26.030 141.090 ;
        RECT 26.430 139.770 26.760 140.750 ;
        RECT 26.980 140.420 27.310 141.090 ;
        RECT 27.710 139.770 28.040 140.750 ;
        RECT 30.350 140.090 30.620 141.950 ;
        RECT 30.800 141.880 30.830 142.050 ;
        RECT 31.000 141.880 31.190 142.050 ;
        RECT 31.360 141.880 31.550 142.050 ;
        RECT 31.720 141.880 31.750 142.050 ;
        RECT 32.440 142.050 33.030 142.080 ;
        RECT 30.800 141.450 31.750 141.880 ;
        RECT 31.930 141.450 32.260 141.950 ;
        RECT 31.480 140.090 31.810 140.590 ;
        RECT 30.350 139.920 31.810 140.090 ;
        RECT 6.260 138.890 9.000 139.770 ;
        RECT 6.260 138.720 6.470 138.890 ;
        RECT 6.640 138.720 6.910 138.890 ;
        RECT 7.080 138.720 7.320 138.890 ;
        RECT 7.490 138.720 7.750 138.890 ;
        RECT 7.920 138.720 8.190 138.890 ;
        RECT 8.360 138.720 8.600 138.890 ;
        RECT 8.770 138.720 9.000 138.890 ;
        RECT 6.260 138.700 9.000 138.720 ;
        RECT 10.100 138.890 12.840 139.770 ;
        RECT 10.100 138.720 10.310 138.890 ;
        RECT 10.480 138.720 10.750 138.890 ;
        RECT 10.920 138.720 11.160 138.890 ;
        RECT 11.330 138.720 11.590 138.890 ;
        RECT 11.760 138.720 12.030 138.890 ;
        RECT 12.200 138.720 12.440 138.890 ;
        RECT 12.610 138.720 12.840 138.890 ;
        RECT 10.100 138.700 12.840 138.720 ;
        RECT 13.940 138.890 16.680 139.770 ;
        RECT 13.940 138.720 14.150 138.890 ;
        RECT 14.320 138.720 14.590 138.890 ;
        RECT 14.760 138.720 15.000 138.890 ;
        RECT 15.170 138.720 15.430 138.890 ;
        RECT 15.600 138.720 15.870 138.890 ;
        RECT 16.040 138.720 16.280 138.890 ;
        RECT 16.450 138.720 16.680 138.890 ;
        RECT 13.940 138.700 16.680 138.720 ;
        RECT 17.780 138.890 20.520 139.770 ;
        RECT 17.780 138.720 17.990 138.890 ;
        RECT 18.160 138.720 18.430 138.890 ;
        RECT 18.600 138.720 18.840 138.890 ;
        RECT 19.010 138.720 19.270 138.890 ;
        RECT 19.440 138.720 19.710 138.890 ;
        RECT 19.880 138.720 20.120 138.890 ;
        RECT 20.290 138.720 20.520 138.890 ;
        RECT 17.780 138.700 20.520 138.720 ;
        RECT 21.620 138.890 24.360 139.770 ;
        RECT 21.620 138.720 21.830 138.890 ;
        RECT 22.000 138.720 22.270 138.890 ;
        RECT 22.440 138.720 22.680 138.890 ;
        RECT 22.850 138.720 23.110 138.890 ;
        RECT 23.280 138.720 23.550 138.890 ;
        RECT 23.720 138.720 23.960 138.890 ;
        RECT 24.130 138.720 24.360 138.890 ;
        RECT 21.620 138.700 24.360 138.720 ;
        RECT 25.460 138.890 28.200 139.770 ;
        RECT 30.350 138.990 30.680 139.920 ;
        RECT 25.460 138.720 25.670 138.890 ;
        RECT 25.840 138.720 26.110 138.890 ;
        RECT 26.280 138.720 26.520 138.890 ;
        RECT 26.690 138.720 26.950 138.890 ;
        RECT 27.120 138.720 27.390 138.890 ;
        RECT 27.560 138.720 27.800 138.890 ;
        RECT 27.970 138.720 28.200 138.890 ;
        RECT 30.870 138.940 31.460 139.720 ;
        RECT 30.870 138.770 30.900 138.940 ;
        RECT 31.070 138.770 31.260 138.940 ;
        RECT 31.430 138.770 31.460 138.940 ;
        RECT 30.870 138.740 31.460 138.770 ;
        RECT 31.640 138.810 31.810 139.920 ;
        RECT 31.990 140.530 32.260 141.450 ;
        RECT 32.440 141.880 32.470 142.050 ;
        RECT 32.640 141.880 32.830 142.050 ;
        RECT 33.000 141.880 33.030 142.050 ;
        RECT 37.400 142.050 38.350 142.080 ;
        RECT 32.440 141.200 33.030 141.880 ;
      LAYER li1 ;
        RECT 33.310 141.820 36.250 141.990 ;
        RECT 33.310 141.610 33.480 141.820 ;
        RECT 33.270 141.440 33.480 141.610 ;
        RECT 33.310 140.830 33.480 141.440 ;
      LAYER li1 ;
        RECT 31.990 140.300 32.520 140.530 ;
        RECT 31.990 138.990 32.240 140.300 ;
      LAYER li1 ;
        RECT 32.940 139.960 33.480 140.830 ;
        RECT 33.660 140.340 33.990 141.640 ;
      LAYER li1 ;
        RECT 34.170 141.120 34.440 141.620 ;
        RECT 34.890 141.370 35.220 141.620 ;
        RECT 34.890 141.200 35.900 141.370 ;
        RECT 34.170 140.130 34.340 141.120 ;
        RECT 35.220 140.530 35.550 141.020 ;
        RECT 34.120 139.960 34.340 140.130 ;
        RECT 34.520 140.300 35.550 140.530 ;
        RECT 35.730 140.970 35.900 141.200 ;
      LAYER li1 ;
        RECT 36.080 141.320 36.250 141.820 ;
      LAYER li1 ;
        RECT 37.400 141.880 37.430 142.050 ;
        RECT 37.600 141.880 37.790 142.050 ;
        RECT 37.960 141.880 38.150 142.050 ;
        RECT 38.320 141.880 38.350 142.050 ;
        RECT 37.400 141.500 38.350 141.880 ;
      LAYER li1 ;
        RECT 38.530 142.010 41.190 142.180 ;
        RECT 38.530 141.320 38.700 142.010 ;
        RECT 36.080 141.150 38.700 141.320 ;
      LAYER li1 ;
        RECT 35.730 140.800 38.350 140.970 ;
        RECT 34.120 139.780 34.290 139.960 ;
        RECT 34.520 139.780 34.690 140.300 ;
        RECT 35.730 140.120 35.900 140.800 ;
      LAYER li1 ;
        RECT 38.530 140.620 38.700 141.150 ;
      LAYER li1 ;
        RECT 32.480 139.610 34.290 139.780 ;
        RECT 32.480 138.990 32.730 139.610 ;
        RECT 32.910 139.260 33.940 139.430 ;
        RECT 32.910 138.810 33.080 139.260 ;
        RECT 25.460 138.700 28.200 138.720 ;
        RECT 31.640 138.640 33.080 138.810 ;
        RECT 33.260 138.940 33.590 139.080 ;
        RECT 33.260 138.770 33.290 138.940 ;
        RECT 33.460 138.770 33.590 138.940 ;
        RECT 33.260 138.740 33.590 138.770 ;
        RECT 33.770 138.810 33.940 139.260 ;
        RECT 34.120 138.990 34.290 139.610 ;
        RECT 34.470 139.450 34.690 139.780 ;
        RECT 34.870 139.950 35.900 140.120 ;
        RECT 36.080 140.270 36.410 140.620 ;
      LAYER li1 ;
        RECT 36.850 140.450 38.700 140.620 ;
      LAYER li1 ;
        RECT 38.880 141.120 39.210 141.830 ;
        RECT 39.670 141.660 40.840 141.830 ;
        RECT 39.670 141.120 40.000 141.660 ;
        RECT 38.880 140.270 39.140 141.120 ;
        RECT 40.210 140.860 40.490 141.360 ;
        RECT 36.080 140.100 39.140 140.270 ;
        RECT 34.870 139.250 35.040 139.950 ;
        RECT 35.730 139.920 35.900 139.950 ;
        RECT 35.220 139.570 35.550 139.770 ;
        RECT 35.730 139.750 37.500 139.920 ;
        RECT 35.220 139.450 36.990 139.570 ;
        RECT 35.340 139.400 36.990 139.450 ;
        RECT 34.820 138.990 35.150 139.250 ;
        RECT 35.340 138.810 35.510 139.400 ;
        RECT 33.770 138.640 35.510 138.810 ;
        RECT 35.690 138.940 36.640 139.220 ;
        RECT 35.690 138.770 35.720 138.940 ;
        RECT 35.890 138.770 36.080 138.940 ;
        RECT 36.250 138.770 36.440 138.940 ;
        RECT 36.610 138.770 36.640 138.940 ;
        RECT 35.690 138.740 36.640 138.770 ;
        RECT 36.820 138.810 36.990 139.400 ;
        RECT 37.170 138.990 37.500 139.750 ;
        RECT 38.810 139.520 39.140 140.100 ;
        RECT 39.320 140.690 40.490 140.860 ;
        RECT 39.320 139.340 39.490 140.690 ;
        RECT 39.870 140.010 40.200 140.510 ;
        RECT 40.670 140.260 40.840 141.660 ;
      LAYER li1 ;
        RECT 41.020 141.350 41.190 142.010 ;
      LAYER li1 ;
        RECT 41.370 142.050 42.320 142.080 ;
        RECT 41.370 141.880 41.400 142.050 ;
        RECT 41.570 141.880 41.760 142.050 ;
        RECT 41.930 141.880 42.120 142.050 ;
        RECT 42.290 141.880 42.320 142.050 ;
        RECT 43.980 142.050 44.930 142.080 ;
        RECT 41.370 141.530 42.320 141.880 ;
        RECT 42.860 141.450 43.190 141.950 ;
        RECT 43.980 141.880 44.010 142.050 ;
        RECT 44.180 141.880 44.370 142.050 ;
        RECT 44.540 141.880 44.730 142.050 ;
        RECT 44.900 141.880 44.930 142.050 ;
      LAYER li1 ;
        RECT 41.020 141.180 42.030 141.350 ;
      LAYER li1 ;
        RECT 41.050 140.610 41.380 141.000 ;
      LAYER li1 ;
        RECT 41.700 140.790 42.030 141.180 ;
      LAYER li1 ;
        RECT 42.860 140.610 43.090 141.450 ;
        RECT 43.470 140.950 43.800 141.450 ;
        RECT 43.980 140.950 44.930 141.880 ;
        RECT 45.770 142.050 47.380 142.080 ;
        RECT 45.770 141.880 45.820 142.050 ;
        RECT 45.990 141.880 46.260 142.050 ;
        RECT 46.430 141.880 46.700 142.050 ;
        RECT 46.870 141.880 47.110 142.050 ;
        RECT 47.280 141.880 47.380 142.050 ;
        RECT 48.080 142.050 49.030 142.080 ;
        RECT 45.770 141.600 47.380 141.880 ;
        RECT 46.080 141.200 47.380 141.600 ;
        RECT 41.050 140.440 43.090 140.610 ;
        RECT 40.380 140.090 42.740 140.260 ;
        RECT 40.380 139.770 40.550 140.090 ;
        RECT 42.920 139.910 43.090 140.440 ;
        RECT 37.680 139.170 39.490 139.340 ;
        RECT 39.670 139.600 40.550 139.770 ;
        RECT 37.680 138.810 37.850 139.170 ;
        RECT 36.820 138.640 37.850 138.810 ;
        RECT 38.030 138.940 38.980 138.990 ;
        RECT 38.030 138.770 38.060 138.940 ;
        RECT 38.230 138.770 38.420 138.940 ;
        RECT 38.590 138.770 38.780 138.940 ;
        RECT 38.950 138.770 38.980 138.940 ;
        RECT 38.030 138.690 38.980 138.770 ;
        RECT 39.670 138.690 39.920 139.600 ;
        RECT 40.730 138.940 41.680 139.770 ;
        RECT 42.080 139.740 43.090 139.910 ;
        RECT 43.590 140.770 43.800 140.950 ;
        RECT 43.590 140.440 44.960 140.770 ;
        RECT 42.080 139.270 42.330 139.740 ;
        RECT 42.510 138.940 43.410 139.560 ;
        RECT 43.590 139.440 43.840 140.440 ;
        RECT 46.080 140.420 46.410 141.200 ;
        RECT 40.730 138.770 40.760 138.940 ;
        RECT 40.930 138.770 41.120 138.940 ;
        RECT 41.290 138.770 41.480 138.940 ;
        RECT 41.650 138.770 41.680 138.940 ;
        RECT 42.680 138.770 42.870 138.940 ;
        RECT 43.040 138.770 43.230 138.940 ;
        RECT 43.400 138.770 43.410 138.940 ;
        RECT 40.730 138.740 41.680 138.770 ;
        RECT 42.510 138.740 43.410 138.770 ;
        RECT 44.020 138.940 44.960 140.250 ;
        RECT 46.620 139.760 46.950 140.750 ;
        RECT 47.630 140.090 47.900 141.950 ;
        RECT 48.080 141.880 48.110 142.050 ;
        RECT 48.280 141.880 48.470 142.050 ;
        RECT 48.640 141.880 48.830 142.050 ;
        RECT 49.000 141.880 49.030 142.050 ;
        RECT 49.720 142.050 50.310 142.080 ;
        RECT 48.080 141.450 49.030 141.880 ;
        RECT 49.210 141.450 49.540 141.950 ;
        RECT 48.760 140.090 49.090 140.590 ;
        RECT 47.630 139.920 49.090 140.090 ;
        RECT 44.020 138.770 44.040 138.940 ;
        RECT 44.210 138.770 44.400 138.940 ;
        RECT 44.570 138.770 44.760 138.940 ;
        RECT 44.930 138.770 44.960 138.940 ;
        RECT 44.020 138.710 44.960 138.770 ;
        RECT 45.850 138.890 47.300 139.760 ;
        RECT 47.630 138.990 47.960 139.920 ;
        RECT 45.850 138.720 46.100 138.890 ;
        RECT 46.270 138.720 46.460 138.890 ;
        RECT 46.630 138.720 46.900 138.890 ;
        RECT 47.070 138.720 47.300 138.890 ;
        RECT 48.150 138.940 48.740 139.720 ;
        RECT 48.150 138.770 48.180 138.940 ;
        RECT 48.350 138.770 48.540 138.940 ;
        RECT 48.710 138.770 48.740 138.940 ;
        RECT 48.150 138.740 48.740 138.770 ;
        RECT 48.920 138.810 49.090 139.920 ;
        RECT 49.270 140.530 49.540 141.450 ;
        RECT 49.720 141.880 49.750 142.050 ;
        RECT 49.920 141.880 50.110 142.050 ;
        RECT 50.280 141.880 50.310 142.050 ;
        RECT 54.680 142.050 55.630 142.080 ;
        RECT 49.720 141.200 50.310 141.880 ;
      LAYER li1 ;
        RECT 50.590 141.820 53.530 141.990 ;
        RECT 50.590 141.610 50.760 141.820 ;
        RECT 50.550 141.440 50.760 141.610 ;
        RECT 50.590 140.830 50.760 141.440 ;
      LAYER li1 ;
        RECT 49.270 140.300 49.800 140.530 ;
        RECT 49.270 138.990 49.520 140.300 ;
      LAYER li1 ;
        RECT 50.220 139.960 50.760 140.830 ;
        RECT 50.940 140.340 51.270 141.640 ;
      LAYER li1 ;
        RECT 51.450 141.120 51.720 141.620 ;
        RECT 52.170 141.370 52.500 141.620 ;
        RECT 52.170 141.200 53.180 141.370 ;
        RECT 51.450 140.130 51.620 141.120 ;
        RECT 52.500 140.530 52.830 141.020 ;
        RECT 51.400 139.960 51.620 140.130 ;
        RECT 51.800 140.300 52.830 140.530 ;
        RECT 53.010 140.970 53.180 141.200 ;
      LAYER li1 ;
        RECT 53.360 141.320 53.530 141.820 ;
      LAYER li1 ;
        RECT 54.680 141.880 54.710 142.050 ;
        RECT 54.880 141.880 55.070 142.050 ;
        RECT 55.240 141.880 55.430 142.050 ;
        RECT 55.600 141.880 55.630 142.050 ;
        RECT 54.680 141.500 55.630 141.880 ;
      LAYER li1 ;
        RECT 55.810 142.010 58.470 142.180 ;
        RECT 55.810 141.320 55.980 142.010 ;
        RECT 53.360 141.150 55.980 141.320 ;
      LAYER li1 ;
        RECT 53.010 140.800 55.630 140.970 ;
        RECT 51.400 139.780 51.570 139.960 ;
        RECT 51.800 139.780 51.970 140.300 ;
        RECT 53.010 140.120 53.180 140.800 ;
      LAYER li1 ;
        RECT 55.810 140.620 55.980 141.150 ;
      LAYER li1 ;
        RECT 49.760 139.610 51.570 139.780 ;
        RECT 49.760 138.990 50.010 139.610 ;
        RECT 50.190 139.260 51.220 139.430 ;
        RECT 50.190 138.810 50.360 139.260 ;
        RECT 45.850 138.690 47.300 138.720 ;
        RECT 48.920 138.640 50.360 138.810 ;
        RECT 50.540 138.940 50.870 139.080 ;
        RECT 50.540 138.770 50.570 138.940 ;
        RECT 50.740 138.770 50.870 138.940 ;
        RECT 50.540 138.740 50.870 138.770 ;
        RECT 51.050 138.810 51.220 139.260 ;
        RECT 51.400 138.990 51.570 139.610 ;
        RECT 51.750 139.450 51.970 139.780 ;
        RECT 52.150 139.950 53.180 140.120 ;
        RECT 53.360 140.270 53.690 140.620 ;
      LAYER li1 ;
        RECT 54.130 140.450 55.980 140.620 ;
      LAYER li1 ;
        RECT 56.160 141.120 56.490 141.830 ;
        RECT 56.950 141.660 58.120 141.830 ;
        RECT 56.950 141.120 57.280 141.660 ;
        RECT 56.160 140.270 56.420 141.120 ;
        RECT 57.490 140.860 57.770 141.360 ;
        RECT 53.360 140.100 56.420 140.270 ;
        RECT 52.150 139.250 52.320 139.950 ;
        RECT 53.010 139.920 53.180 139.950 ;
        RECT 52.500 139.570 52.830 139.770 ;
        RECT 53.010 139.750 54.780 139.920 ;
        RECT 52.500 139.450 54.270 139.570 ;
        RECT 52.620 139.400 54.270 139.450 ;
        RECT 52.100 138.990 52.430 139.250 ;
        RECT 52.620 138.810 52.790 139.400 ;
        RECT 51.050 138.640 52.790 138.810 ;
        RECT 52.970 138.940 53.920 139.220 ;
        RECT 52.970 138.770 53.000 138.940 ;
        RECT 53.170 138.770 53.360 138.940 ;
        RECT 53.530 138.770 53.720 138.940 ;
        RECT 53.890 138.770 53.920 138.940 ;
        RECT 52.970 138.740 53.920 138.770 ;
        RECT 54.100 138.810 54.270 139.400 ;
        RECT 54.450 138.990 54.780 139.750 ;
        RECT 56.090 139.520 56.420 140.100 ;
        RECT 56.600 140.690 57.770 140.860 ;
        RECT 56.600 139.340 56.770 140.690 ;
        RECT 57.150 140.010 57.480 140.510 ;
        RECT 57.950 140.260 58.120 141.660 ;
      LAYER li1 ;
        RECT 58.300 141.350 58.470 142.010 ;
      LAYER li1 ;
        RECT 58.650 142.050 59.600 142.080 ;
        RECT 58.650 141.880 58.680 142.050 ;
        RECT 58.850 141.880 59.040 142.050 ;
        RECT 59.210 141.880 59.400 142.050 ;
        RECT 59.570 141.880 59.600 142.050 ;
        RECT 61.260 142.050 62.210 142.080 ;
        RECT 58.650 141.530 59.600 141.880 ;
        RECT 60.140 141.450 60.470 141.950 ;
        RECT 61.260 141.880 61.290 142.050 ;
        RECT 61.460 141.880 61.650 142.050 ;
        RECT 61.820 141.880 62.010 142.050 ;
        RECT 62.180 141.880 62.210 142.050 ;
      LAYER li1 ;
        RECT 58.300 141.180 59.310 141.350 ;
      LAYER li1 ;
        RECT 58.330 140.610 58.660 141.000 ;
      LAYER li1 ;
        RECT 58.980 140.790 59.310 141.180 ;
      LAYER li1 ;
        RECT 60.140 140.610 60.370 141.450 ;
        RECT 60.750 140.950 61.080 141.450 ;
        RECT 61.260 140.950 62.210 141.880 ;
        RECT 63.050 142.050 64.660 142.080 ;
        RECT 65.350 142.050 66.600 142.080 ;
        RECT 67.780 142.060 70.510 142.090 ;
        RECT 63.050 141.880 63.100 142.050 ;
        RECT 63.270 141.880 63.540 142.050 ;
        RECT 63.710 141.880 63.980 142.050 ;
        RECT 64.150 141.880 64.390 142.050 ;
        RECT 64.560 141.880 64.660 142.050 ;
        RECT 63.050 141.600 64.660 141.880 ;
        RECT 63.360 141.200 64.660 141.600 ;
        RECT 58.330 140.440 60.370 140.610 ;
        RECT 57.660 140.090 60.020 140.260 ;
        RECT 57.660 139.770 57.830 140.090 ;
        RECT 60.200 139.910 60.370 140.440 ;
        RECT 54.960 139.170 56.770 139.340 ;
        RECT 56.950 139.600 57.830 139.770 ;
        RECT 54.960 138.810 55.130 139.170 ;
        RECT 54.100 138.640 55.130 138.810 ;
        RECT 55.310 138.940 56.260 138.990 ;
        RECT 55.310 138.770 55.340 138.940 ;
        RECT 55.510 138.770 55.700 138.940 ;
        RECT 55.870 138.770 56.060 138.940 ;
        RECT 56.230 138.770 56.260 138.940 ;
        RECT 55.310 138.690 56.260 138.770 ;
        RECT 56.950 138.690 57.200 139.600 ;
        RECT 58.010 138.940 58.960 139.770 ;
        RECT 59.360 139.740 60.370 139.910 ;
        RECT 60.870 140.770 61.080 140.950 ;
        RECT 60.870 140.440 62.240 140.770 ;
        RECT 59.360 139.270 59.610 139.740 ;
        RECT 59.790 138.940 60.690 139.560 ;
        RECT 60.870 139.440 61.120 140.440 ;
        RECT 63.360 140.420 63.690 141.200 ;
        RECT 58.010 138.770 58.040 138.940 ;
        RECT 58.210 138.770 58.400 138.940 ;
        RECT 58.570 138.770 58.760 138.940 ;
        RECT 58.930 138.770 58.960 138.940 ;
        RECT 59.960 138.770 60.150 138.940 ;
        RECT 60.320 138.770 60.510 138.940 ;
        RECT 60.680 138.770 60.690 138.940 ;
        RECT 58.010 138.740 58.960 138.770 ;
        RECT 59.790 138.740 60.690 138.770 ;
        RECT 61.300 138.940 62.240 140.250 ;
        RECT 63.900 139.760 64.230 140.750 ;
      LAYER li1 ;
        RECT 64.920 140.270 65.170 141.950 ;
      LAYER li1 ;
        RECT 65.520 141.880 65.710 142.050 ;
        RECT 65.880 141.880 66.070 142.050 ;
        RECT 66.240 141.880 66.430 142.050 ;
        RECT 65.350 141.510 66.600 141.880 ;
        RECT 66.780 141.330 67.030 141.950 ;
        RECT 65.480 141.160 67.030 141.330 ;
        RECT 65.480 140.700 65.810 141.160 ;
        RECT 61.300 138.770 61.320 138.940 ;
        RECT 61.490 138.770 61.680 138.940 ;
        RECT 61.850 138.770 62.040 138.940 ;
        RECT 62.210 138.770 62.240 138.940 ;
        RECT 61.300 138.710 62.240 138.770 ;
        RECT 63.130 138.890 64.580 139.760 ;
        RECT 63.130 138.720 63.380 138.890 ;
        RECT 63.550 138.720 63.740 138.890 ;
        RECT 63.910 138.720 64.180 138.890 ;
        RECT 64.350 138.720 64.580 138.890 ;
        RECT 63.130 138.690 64.580 138.720 ;
      LAYER li1 ;
        RECT 64.920 138.690 65.350 140.270 ;
      LAYER li1 ;
        RECT 65.530 138.940 66.090 140.270 ;
      LAYER li1 ;
        RECT 66.270 139.190 66.600 140.980 ;
      LAYER li1 ;
        RECT 66.780 139.440 67.030 141.160 ;
        RECT 67.780 141.890 67.950 142.060 ;
        RECT 68.120 141.890 68.390 142.060 ;
        RECT 68.560 141.890 68.800 142.060 ;
        RECT 68.970 141.890 69.230 142.060 ;
        RECT 69.400 141.890 69.670 142.060 ;
        RECT 69.840 141.890 70.080 142.060 ;
        RECT 70.250 141.890 70.510 142.060 ;
        RECT 67.780 141.090 70.510 141.890 ;
        RECT 71.130 142.050 71.720 142.080 ;
        RECT 71.130 141.880 71.160 142.050 ;
        RECT 71.330 141.880 71.520 142.050 ;
        RECT 71.690 141.880 71.720 142.050 ;
        RECT 72.650 142.050 74.260 142.080 ;
        RECT 74.950 142.050 76.200 142.080 ;
        RECT 76.970 142.050 78.580 142.080 ;
        RECT 71.130 141.120 71.720 141.880 ;
        RECT 67.940 140.420 68.270 141.090 ;
        RECT 68.670 139.770 69.000 140.750 ;
        RECT 69.220 140.420 69.550 141.090 ;
        RECT 69.950 139.770 70.280 140.750 ;
      LAYER li1 ;
        RECT 71.170 140.510 71.880 140.900 ;
        RECT 72.060 140.270 72.390 141.950 ;
      LAYER li1 ;
        RECT 72.650 141.880 72.700 142.050 ;
        RECT 72.870 141.880 73.140 142.050 ;
        RECT 73.310 141.880 73.580 142.050 ;
        RECT 73.750 141.880 73.990 142.050 ;
        RECT 74.160 141.880 74.260 142.050 ;
        RECT 72.650 141.600 74.260 141.880 ;
        RECT 72.960 141.200 74.260 141.600 ;
        RECT 72.960 140.420 73.290 141.200 ;
        RECT 65.530 138.770 65.540 138.940 ;
        RECT 65.710 138.770 65.900 138.940 ;
        RECT 66.070 138.770 66.090 138.940 ;
        RECT 65.530 138.690 66.090 138.770 ;
        RECT 67.700 138.890 70.440 139.770 ;
        RECT 67.700 138.720 67.910 138.890 ;
        RECT 68.080 138.720 68.350 138.890 ;
        RECT 68.520 138.720 68.760 138.890 ;
        RECT 68.930 138.720 69.190 138.890 ;
        RECT 69.360 138.720 69.630 138.890 ;
        RECT 69.800 138.720 70.040 138.890 ;
        RECT 70.210 138.720 70.440 138.890 ;
        RECT 67.700 138.700 70.440 138.720 ;
        RECT 71.130 138.940 71.720 140.270 ;
        RECT 71.130 138.770 71.160 138.940 ;
        RECT 71.330 138.770 71.520 138.940 ;
        RECT 71.690 138.770 71.720 138.940 ;
        RECT 71.130 138.690 71.720 138.770 ;
      LAYER li1 ;
        RECT 72.000 138.690 72.390 140.270 ;
      LAYER li1 ;
        RECT 73.500 139.760 73.830 140.750 ;
      LAYER li1 ;
        RECT 74.520 140.270 74.770 141.950 ;
      LAYER li1 ;
        RECT 75.120 141.880 75.310 142.050 ;
        RECT 75.480 141.880 75.670 142.050 ;
        RECT 75.840 141.880 76.030 142.050 ;
        RECT 74.950 141.510 76.200 141.880 ;
        RECT 76.380 141.330 76.630 141.950 ;
        RECT 76.970 141.880 77.020 142.050 ;
        RECT 77.190 141.880 77.460 142.050 ;
        RECT 77.630 141.880 77.900 142.050 ;
        RECT 78.070 141.880 78.310 142.050 ;
        RECT 78.480 141.880 78.580 142.050 ;
        RECT 79.280 142.050 80.230 142.080 ;
        RECT 76.970 141.600 78.580 141.880 ;
        RECT 75.080 141.160 76.630 141.330 ;
        RECT 75.080 140.700 75.410 141.160 ;
        RECT 72.730 138.890 74.180 139.760 ;
        RECT 72.730 138.720 72.980 138.890 ;
        RECT 73.150 138.720 73.340 138.890 ;
        RECT 73.510 138.720 73.780 138.890 ;
        RECT 73.950 138.720 74.180 138.890 ;
        RECT 72.730 138.690 74.180 138.720 ;
      LAYER li1 ;
        RECT 74.520 138.690 74.950 140.270 ;
      LAYER li1 ;
        RECT 75.130 138.940 75.690 140.270 ;
      LAYER li1 ;
        RECT 75.870 139.190 76.200 140.980 ;
      LAYER li1 ;
        RECT 76.380 139.440 76.630 141.160 ;
        RECT 77.280 141.200 78.580 141.600 ;
        RECT 77.280 140.420 77.610 141.200 ;
        RECT 77.820 139.760 78.150 140.750 ;
        RECT 78.830 140.090 79.100 141.950 ;
        RECT 79.280 141.880 79.310 142.050 ;
        RECT 79.480 141.880 79.670 142.050 ;
        RECT 79.840 141.880 80.030 142.050 ;
        RECT 80.200 141.880 80.230 142.050 ;
        RECT 80.920 142.050 81.510 142.080 ;
        RECT 79.280 141.450 80.230 141.880 ;
        RECT 80.410 141.450 80.740 141.950 ;
      LAYER li1 ;
        RECT 79.280 140.300 79.610 141.270 ;
      LAYER li1 ;
        RECT 79.960 140.090 80.290 140.590 ;
        RECT 78.830 139.920 80.290 140.090 ;
        RECT 75.130 138.770 75.140 138.940 ;
        RECT 75.310 138.770 75.500 138.940 ;
        RECT 75.670 138.770 75.690 138.940 ;
        RECT 75.130 138.690 75.690 138.770 ;
        RECT 77.050 138.890 78.500 139.760 ;
        RECT 78.830 138.990 79.160 139.920 ;
        RECT 77.050 138.720 77.300 138.890 ;
        RECT 77.470 138.720 77.660 138.890 ;
        RECT 77.830 138.720 78.100 138.890 ;
        RECT 78.270 138.720 78.500 138.890 ;
        RECT 79.350 138.940 79.940 139.720 ;
        RECT 79.350 138.770 79.380 138.940 ;
        RECT 79.550 138.770 79.740 138.940 ;
        RECT 79.910 138.770 79.940 138.940 ;
        RECT 79.350 138.740 79.940 138.770 ;
        RECT 80.120 138.810 80.290 139.920 ;
        RECT 80.470 140.530 80.740 141.450 ;
        RECT 80.920 141.880 80.950 142.050 ;
        RECT 81.120 141.880 81.310 142.050 ;
        RECT 81.480 141.880 81.510 142.050 ;
        RECT 85.880 142.050 86.830 142.080 ;
        RECT 80.920 141.200 81.510 141.880 ;
      LAYER li1 ;
        RECT 81.790 141.820 84.730 141.990 ;
        RECT 81.790 141.610 81.960 141.820 ;
        RECT 81.750 141.440 81.960 141.610 ;
        RECT 81.790 140.830 81.960 141.440 ;
      LAYER li1 ;
        RECT 80.470 140.300 81.000 140.530 ;
        RECT 80.470 138.990 80.720 140.300 ;
      LAYER li1 ;
        RECT 81.420 139.960 81.960 140.830 ;
        RECT 82.140 140.340 82.470 141.640 ;
      LAYER li1 ;
        RECT 82.650 141.120 82.920 141.620 ;
        RECT 83.370 141.370 83.700 141.620 ;
        RECT 83.370 141.200 84.380 141.370 ;
        RECT 82.650 140.130 82.820 141.120 ;
        RECT 83.700 140.530 84.030 141.020 ;
        RECT 82.600 139.960 82.820 140.130 ;
        RECT 83.000 140.300 84.030 140.530 ;
        RECT 84.210 140.970 84.380 141.200 ;
      LAYER li1 ;
        RECT 84.560 141.320 84.730 141.820 ;
      LAYER li1 ;
        RECT 85.880 141.880 85.910 142.050 ;
        RECT 86.080 141.880 86.270 142.050 ;
        RECT 86.440 141.880 86.630 142.050 ;
        RECT 86.800 141.880 86.830 142.050 ;
        RECT 85.880 141.500 86.830 141.880 ;
      LAYER li1 ;
        RECT 87.010 142.010 89.670 142.180 ;
        RECT 87.010 141.320 87.180 142.010 ;
        RECT 84.560 141.150 87.180 141.320 ;
      LAYER li1 ;
        RECT 84.210 140.800 86.830 140.970 ;
        RECT 82.600 139.780 82.770 139.960 ;
        RECT 83.000 139.780 83.170 140.300 ;
        RECT 84.210 140.120 84.380 140.800 ;
      LAYER li1 ;
        RECT 87.010 140.620 87.180 141.150 ;
      LAYER li1 ;
        RECT 80.960 139.610 82.770 139.780 ;
        RECT 80.960 138.990 81.210 139.610 ;
        RECT 81.390 139.260 82.420 139.430 ;
        RECT 81.390 138.810 81.560 139.260 ;
        RECT 77.050 138.690 78.500 138.720 ;
        RECT 80.120 138.640 81.560 138.810 ;
        RECT 81.740 138.940 82.070 139.080 ;
        RECT 81.740 138.770 81.770 138.940 ;
        RECT 81.940 138.770 82.070 138.940 ;
        RECT 81.740 138.740 82.070 138.770 ;
        RECT 82.250 138.810 82.420 139.260 ;
        RECT 82.600 138.990 82.770 139.610 ;
        RECT 82.950 139.450 83.170 139.780 ;
        RECT 83.350 139.950 84.380 140.120 ;
        RECT 84.560 140.270 84.890 140.620 ;
      LAYER li1 ;
        RECT 85.330 140.450 87.180 140.620 ;
      LAYER li1 ;
        RECT 87.360 141.120 87.690 141.830 ;
        RECT 88.150 141.660 89.320 141.830 ;
        RECT 88.150 141.120 88.480 141.660 ;
        RECT 87.360 140.270 87.620 141.120 ;
        RECT 88.690 140.860 88.970 141.360 ;
        RECT 84.560 140.100 87.620 140.270 ;
        RECT 83.350 139.250 83.520 139.950 ;
        RECT 84.210 139.920 84.380 139.950 ;
        RECT 83.700 139.570 84.030 139.770 ;
        RECT 84.210 139.750 85.980 139.920 ;
        RECT 83.700 139.450 85.470 139.570 ;
        RECT 83.820 139.400 85.470 139.450 ;
        RECT 83.300 138.990 83.630 139.250 ;
        RECT 83.820 138.810 83.990 139.400 ;
        RECT 82.250 138.640 83.990 138.810 ;
        RECT 84.170 138.940 85.120 139.220 ;
        RECT 84.170 138.770 84.200 138.940 ;
        RECT 84.370 138.770 84.560 138.940 ;
        RECT 84.730 138.770 84.920 138.940 ;
        RECT 85.090 138.770 85.120 138.940 ;
        RECT 84.170 138.740 85.120 138.770 ;
        RECT 85.300 138.810 85.470 139.400 ;
        RECT 85.650 138.990 85.980 139.750 ;
        RECT 87.290 139.520 87.620 140.100 ;
        RECT 87.800 140.690 88.970 140.860 ;
        RECT 87.800 139.340 87.970 140.690 ;
        RECT 88.350 140.010 88.680 140.510 ;
        RECT 89.150 140.260 89.320 141.660 ;
      LAYER li1 ;
        RECT 89.500 141.350 89.670 142.010 ;
      LAYER li1 ;
        RECT 89.850 142.050 90.800 142.080 ;
        RECT 89.850 141.880 89.880 142.050 ;
        RECT 90.050 141.880 90.240 142.050 ;
        RECT 90.410 141.880 90.600 142.050 ;
        RECT 90.770 141.880 90.800 142.050 ;
        RECT 92.460 142.050 93.410 142.080 ;
        RECT 89.850 141.530 90.800 141.880 ;
        RECT 91.340 141.450 91.670 141.950 ;
        RECT 92.460 141.880 92.490 142.050 ;
        RECT 92.660 141.880 92.850 142.050 ;
        RECT 93.020 141.880 93.210 142.050 ;
        RECT 93.380 141.880 93.410 142.050 ;
      LAYER li1 ;
        RECT 89.500 141.180 90.510 141.350 ;
      LAYER li1 ;
        RECT 89.530 140.610 89.860 141.000 ;
      LAYER li1 ;
        RECT 90.180 140.790 90.510 141.180 ;
      LAYER li1 ;
        RECT 91.340 140.610 91.570 141.450 ;
        RECT 91.950 140.950 92.280 141.450 ;
        RECT 92.460 140.950 93.410 141.880 ;
        RECT 94.660 142.060 97.390 142.090 ;
        RECT 94.660 141.890 94.830 142.060 ;
        RECT 95.000 141.890 95.270 142.060 ;
        RECT 95.440 141.890 95.680 142.060 ;
        RECT 95.850 141.890 96.110 142.060 ;
        RECT 96.280 141.890 96.550 142.060 ;
        RECT 96.720 141.890 96.960 142.060 ;
        RECT 97.130 141.890 97.390 142.060 ;
        RECT 98.480 142.050 99.430 142.080 ;
        RECT 89.530 140.440 91.570 140.610 ;
        RECT 88.860 140.090 91.220 140.260 ;
        RECT 88.860 139.770 89.030 140.090 ;
        RECT 91.400 139.910 91.570 140.440 ;
        RECT 86.160 139.170 87.970 139.340 ;
        RECT 88.150 139.600 89.030 139.770 ;
        RECT 86.160 138.810 86.330 139.170 ;
        RECT 85.300 138.640 86.330 138.810 ;
        RECT 86.510 138.940 87.460 138.990 ;
        RECT 86.510 138.770 86.540 138.940 ;
        RECT 86.710 138.770 86.900 138.940 ;
        RECT 87.070 138.770 87.260 138.940 ;
        RECT 87.430 138.770 87.460 138.940 ;
        RECT 86.510 138.690 87.460 138.770 ;
        RECT 88.150 138.690 88.400 139.600 ;
        RECT 89.210 138.940 90.160 139.770 ;
        RECT 90.560 139.740 91.570 139.910 ;
        RECT 92.070 140.770 92.280 140.950 ;
        RECT 92.070 140.440 93.440 140.770 ;
        RECT 90.560 139.270 90.810 139.740 ;
        RECT 90.990 138.940 91.890 139.560 ;
        RECT 92.070 139.440 92.320 140.440 ;
        RECT 89.210 138.770 89.240 138.940 ;
        RECT 89.410 138.770 89.600 138.940 ;
        RECT 89.770 138.770 89.960 138.940 ;
        RECT 90.130 138.770 90.160 138.940 ;
        RECT 91.160 138.770 91.350 138.940 ;
        RECT 91.520 138.770 91.710 138.940 ;
        RECT 91.880 138.770 91.890 138.940 ;
        RECT 89.210 138.740 90.160 138.770 ;
        RECT 90.990 138.740 91.890 138.770 ;
        RECT 92.500 138.940 93.440 140.250 ;
        RECT 92.500 138.770 92.520 138.940 ;
        RECT 92.690 138.770 92.880 138.940 ;
        RECT 93.050 138.770 93.240 138.940 ;
        RECT 93.410 138.770 93.440 138.940 ;
        RECT 92.500 138.710 93.440 138.770 ;
      LAYER li1 ;
        RECT 93.620 138.710 93.960 141.780 ;
      LAYER li1 ;
        RECT 94.660 141.090 97.390 141.890 ;
        RECT 94.820 140.420 95.150 141.090 ;
        RECT 95.550 139.770 95.880 140.750 ;
        RECT 96.100 140.420 96.430 141.090 ;
        RECT 96.830 139.770 97.160 140.750 ;
        RECT 98.030 140.090 98.300 141.950 ;
        RECT 98.480 141.880 98.510 142.050 ;
        RECT 98.680 141.880 98.870 142.050 ;
        RECT 99.040 141.880 99.230 142.050 ;
        RECT 99.400 141.880 99.430 142.050 ;
        RECT 100.120 142.050 100.710 142.080 ;
        RECT 98.480 141.450 99.430 141.880 ;
        RECT 99.610 141.450 99.940 141.950 ;
      LAYER li1 ;
        RECT 98.480 140.300 98.810 141.270 ;
      LAYER li1 ;
        RECT 99.160 140.090 99.490 140.590 ;
        RECT 98.030 139.920 99.490 140.090 ;
        RECT 94.580 138.890 97.320 139.770 ;
        RECT 98.030 138.990 98.360 139.920 ;
        RECT 94.580 138.720 94.790 138.890 ;
        RECT 94.960 138.720 95.230 138.890 ;
        RECT 95.400 138.720 95.640 138.890 ;
        RECT 95.810 138.720 96.070 138.890 ;
        RECT 96.240 138.720 96.510 138.890 ;
        RECT 96.680 138.720 96.920 138.890 ;
        RECT 97.090 138.720 97.320 138.890 ;
        RECT 98.550 138.940 99.140 139.720 ;
        RECT 98.550 138.770 98.580 138.940 ;
        RECT 98.750 138.770 98.940 138.940 ;
        RECT 99.110 138.770 99.140 138.940 ;
        RECT 98.550 138.740 99.140 138.770 ;
        RECT 99.320 138.810 99.490 139.920 ;
        RECT 99.670 140.530 99.940 141.450 ;
        RECT 100.120 141.880 100.150 142.050 ;
        RECT 100.320 141.880 100.510 142.050 ;
        RECT 100.680 141.880 100.710 142.050 ;
        RECT 105.080 142.050 106.030 142.080 ;
        RECT 100.120 141.200 100.710 141.880 ;
      LAYER li1 ;
        RECT 100.990 141.820 103.930 141.990 ;
        RECT 100.990 140.830 101.160 141.820 ;
      LAYER li1 ;
        RECT 99.670 140.300 100.200 140.530 ;
        RECT 99.670 138.990 99.920 140.300 ;
      LAYER li1 ;
        RECT 100.620 139.960 101.160 140.830 ;
        RECT 101.340 140.340 101.670 141.640 ;
      LAYER li1 ;
        RECT 101.850 141.120 102.120 141.620 ;
        RECT 102.570 141.370 102.900 141.620 ;
        RECT 102.570 141.200 103.580 141.370 ;
        RECT 101.850 140.130 102.020 141.120 ;
        RECT 102.900 140.530 103.230 141.020 ;
        RECT 101.800 139.960 102.020 140.130 ;
        RECT 102.200 140.300 103.230 140.530 ;
        RECT 103.410 140.970 103.580 141.200 ;
      LAYER li1 ;
        RECT 103.760 141.320 103.930 141.820 ;
      LAYER li1 ;
        RECT 105.080 141.880 105.110 142.050 ;
        RECT 105.280 141.880 105.470 142.050 ;
        RECT 105.640 141.880 105.830 142.050 ;
        RECT 106.000 141.880 106.030 142.050 ;
        RECT 105.080 141.500 106.030 141.880 ;
      LAYER li1 ;
        RECT 106.210 142.010 108.870 142.180 ;
        RECT 106.210 141.320 106.380 142.010 ;
        RECT 103.760 141.150 106.380 141.320 ;
      LAYER li1 ;
        RECT 103.410 140.800 106.030 140.970 ;
        RECT 101.800 139.780 101.970 139.960 ;
        RECT 102.200 139.780 102.370 140.300 ;
        RECT 103.410 140.120 103.580 140.800 ;
      LAYER li1 ;
        RECT 106.210 140.620 106.380 141.150 ;
      LAYER li1 ;
        RECT 100.160 139.610 101.970 139.780 ;
        RECT 100.160 138.990 100.410 139.610 ;
        RECT 100.590 139.260 101.620 139.430 ;
        RECT 100.590 138.810 100.760 139.260 ;
        RECT 94.580 138.700 97.320 138.720 ;
        RECT 99.320 138.640 100.760 138.810 ;
        RECT 100.940 138.940 101.270 139.080 ;
        RECT 100.940 138.770 100.970 138.940 ;
        RECT 101.140 138.770 101.270 138.940 ;
        RECT 100.940 138.740 101.270 138.770 ;
        RECT 101.450 138.810 101.620 139.260 ;
        RECT 101.800 138.990 101.970 139.610 ;
        RECT 102.150 139.450 102.370 139.780 ;
        RECT 102.550 139.950 103.580 140.120 ;
        RECT 103.760 140.270 104.090 140.620 ;
      LAYER li1 ;
        RECT 104.530 140.450 106.380 140.620 ;
      LAYER li1 ;
        RECT 106.560 141.120 106.890 141.830 ;
        RECT 107.350 141.660 108.520 141.830 ;
        RECT 107.350 141.120 107.680 141.660 ;
        RECT 106.560 140.270 106.820 141.120 ;
        RECT 107.890 140.860 108.170 141.360 ;
        RECT 103.760 140.100 106.820 140.270 ;
        RECT 102.550 139.250 102.720 139.950 ;
        RECT 103.410 139.920 103.580 139.950 ;
        RECT 102.900 139.570 103.230 139.770 ;
        RECT 103.410 139.750 105.180 139.920 ;
        RECT 102.900 139.450 104.670 139.570 ;
        RECT 103.020 139.400 104.670 139.450 ;
        RECT 102.500 138.990 102.830 139.250 ;
        RECT 103.020 138.810 103.190 139.400 ;
        RECT 101.450 138.640 103.190 138.810 ;
        RECT 103.370 138.940 104.320 139.220 ;
        RECT 103.370 138.770 103.400 138.940 ;
        RECT 103.570 138.770 103.760 138.940 ;
        RECT 103.930 138.770 104.120 138.940 ;
        RECT 104.290 138.770 104.320 138.940 ;
        RECT 103.370 138.740 104.320 138.770 ;
        RECT 104.500 138.810 104.670 139.400 ;
        RECT 104.850 138.990 105.180 139.750 ;
        RECT 106.490 139.520 106.820 140.100 ;
        RECT 107.000 140.690 108.170 140.860 ;
        RECT 107.000 139.340 107.170 140.690 ;
        RECT 107.550 140.010 107.880 140.510 ;
        RECT 108.350 140.260 108.520 141.660 ;
      LAYER li1 ;
        RECT 108.700 141.350 108.870 142.010 ;
      LAYER li1 ;
        RECT 109.050 142.050 110.000 142.080 ;
        RECT 109.050 141.880 109.080 142.050 ;
        RECT 109.250 141.880 109.440 142.050 ;
        RECT 109.610 141.880 109.800 142.050 ;
        RECT 109.970 141.880 110.000 142.050 ;
        RECT 111.660 142.050 112.610 142.080 ;
        RECT 109.050 141.530 110.000 141.880 ;
        RECT 110.540 141.450 110.870 141.950 ;
        RECT 111.660 141.880 111.690 142.050 ;
        RECT 111.860 141.880 112.050 142.050 ;
        RECT 112.220 141.880 112.410 142.050 ;
        RECT 112.580 141.880 112.610 142.050 ;
      LAYER li1 ;
        RECT 108.700 141.240 109.710 141.350 ;
        RECT 108.700 141.180 109.760 141.240 ;
        RECT 109.380 141.070 109.760 141.180 ;
      LAYER li1 ;
        RECT 108.730 140.610 109.060 141.000 ;
      LAYER li1 ;
        RECT 109.380 140.790 109.710 141.070 ;
      LAYER li1 ;
        RECT 110.540 140.610 110.770 141.450 ;
        RECT 111.150 140.950 111.480 141.450 ;
        RECT 111.660 140.950 112.610 141.880 ;
        RECT 113.860 142.060 116.590 142.090 ;
        RECT 113.860 141.890 114.030 142.060 ;
        RECT 114.200 141.890 114.470 142.060 ;
        RECT 114.640 141.890 114.880 142.060 ;
        RECT 115.050 141.890 115.310 142.060 ;
        RECT 115.480 141.890 115.750 142.060 ;
        RECT 115.920 141.890 116.160 142.060 ;
        RECT 116.330 141.890 116.590 142.060 ;
        RECT 108.730 140.440 110.770 140.610 ;
        RECT 108.060 140.090 110.420 140.260 ;
        RECT 108.060 139.770 108.230 140.090 ;
        RECT 110.600 139.910 110.770 140.440 ;
        RECT 105.360 139.170 107.170 139.340 ;
        RECT 107.350 139.600 108.230 139.770 ;
        RECT 105.360 138.810 105.530 139.170 ;
        RECT 104.500 138.640 105.530 138.810 ;
        RECT 105.710 138.940 106.660 138.990 ;
        RECT 105.710 138.770 105.740 138.940 ;
        RECT 105.910 138.770 106.100 138.940 ;
        RECT 106.270 138.770 106.460 138.940 ;
        RECT 106.630 138.770 106.660 138.940 ;
        RECT 105.710 138.690 106.660 138.770 ;
        RECT 107.350 138.690 107.600 139.600 ;
        RECT 108.410 138.940 109.360 139.770 ;
        RECT 109.760 139.740 110.770 139.910 ;
        RECT 111.270 140.770 111.480 140.950 ;
        RECT 111.270 140.440 112.640 140.770 ;
        RECT 109.760 139.270 110.010 139.740 ;
        RECT 110.190 138.940 111.090 139.560 ;
        RECT 111.270 139.440 111.520 140.440 ;
        RECT 108.410 138.770 108.440 138.940 ;
        RECT 108.610 138.770 108.800 138.940 ;
        RECT 108.970 138.770 109.160 138.940 ;
        RECT 109.330 138.770 109.360 138.940 ;
        RECT 110.360 138.770 110.550 138.940 ;
        RECT 110.720 138.770 110.910 138.940 ;
        RECT 111.080 138.770 111.090 138.940 ;
        RECT 108.410 138.740 109.360 138.770 ;
        RECT 110.190 138.740 111.090 138.770 ;
        RECT 111.700 138.940 112.640 140.250 ;
        RECT 111.700 138.770 111.720 138.940 ;
        RECT 111.890 138.770 112.080 138.940 ;
        RECT 112.250 138.770 112.440 138.940 ;
        RECT 112.610 138.770 112.640 138.940 ;
        RECT 111.700 138.710 112.640 138.770 ;
      LAYER li1 ;
        RECT 112.820 138.710 113.160 141.780 ;
      LAYER li1 ;
        RECT 113.860 141.090 116.590 141.890 ;
        RECT 117.700 142.060 120.430 142.090 ;
        RECT 117.700 141.890 117.870 142.060 ;
        RECT 118.040 141.890 118.310 142.060 ;
        RECT 118.480 141.890 118.720 142.060 ;
        RECT 118.890 141.890 119.150 142.060 ;
        RECT 119.320 141.890 119.590 142.060 ;
        RECT 119.760 141.890 120.000 142.060 ;
        RECT 120.170 141.890 120.430 142.060 ;
        RECT 117.700 141.090 120.430 141.890 ;
        RECT 121.540 142.060 124.270 142.090 ;
        RECT 121.540 141.890 121.710 142.060 ;
        RECT 121.880 141.890 122.150 142.060 ;
        RECT 122.320 141.890 122.560 142.060 ;
        RECT 122.730 141.890 122.990 142.060 ;
        RECT 123.160 141.890 123.430 142.060 ;
        RECT 123.600 141.890 123.840 142.060 ;
        RECT 124.010 141.890 124.270 142.060 ;
        RECT 121.540 141.090 124.270 141.890 ;
        RECT 125.380 142.060 128.110 142.090 ;
        RECT 125.380 141.890 125.550 142.060 ;
        RECT 125.720 141.890 125.990 142.060 ;
        RECT 126.160 141.890 126.400 142.060 ;
        RECT 126.570 141.890 126.830 142.060 ;
        RECT 127.000 141.890 127.270 142.060 ;
        RECT 127.440 141.890 127.680 142.060 ;
        RECT 127.850 141.890 128.110 142.060 ;
        RECT 125.380 141.090 128.110 141.890 ;
        RECT 129.220 142.060 131.950 142.090 ;
        RECT 129.220 141.890 129.390 142.060 ;
        RECT 129.560 141.890 129.830 142.060 ;
        RECT 130.000 141.890 130.240 142.060 ;
        RECT 130.410 141.890 130.670 142.060 ;
        RECT 130.840 141.890 131.110 142.060 ;
        RECT 131.280 141.890 131.520 142.060 ;
        RECT 131.690 141.890 131.950 142.060 ;
        RECT 129.220 141.090 131.950 141.890 ;
        RECT 133.060 142.060 135.790 142.090 ;
        RECT 133.060 141.890 133.230 142.060 ;
        RECT 133.400 141.890 133.670 142.060 ;
        RECT 133.840 141.890 134.080 142.060 ;
        RECT 134.250 141.890 134.510 142.060 ;
        RECT 134.680 141.890 134.950 142.060 ;
        RECT 135.120 141.890 135.360 142.060 ;
        RECT 135.530 141.890 135.790 142.060 ;
        RECT 133.060 141.090 135.790 141.890 ;
        RECT 136.900 142.060 139.630 142.090 ;
        RECT 136.900 141.890 137.070 142.060 ;
        RECT 137.240 141.890 137.510 142.060 ;
        RECT 137.680 141.890 137.920 142.060 ;
        RECT 138.090 141.890 138.350 142.060 ;
        RECT 138.520 141.890 138.790 142.060 ;
        RECT 138.960 141.890 139.200 142.060 ;
        RECT 139.370 141.890 139.630 142.060 ;
        RECT 136.900 141.090 139.630 141.890 ;
        RECT 140.330 142.050 141.940 142.080 ;
        RECT 140.330 141.880 140.380 142.050 ;
        RECT 140.550 141.880 140.820 142.050 ;
        RECT 140.990 141.880 141.260 142.050 ;
        RECT 141.430 141.880 141.670 142.050 ;
        RECT 141.840 141.880 141.940 142.050 ;
        RECT 140.330 141.600 141.940 141.880 ;
        RECT 140.640 141.200 141.940 141.600 ;
        RECT 114.020 140.420 114.350 141.090 ;
        RECT 114.750 139.770 115.080 140.750 ;
        RECT 115.300 140.420 115.630 141.090 ;
        RECT 116.030 139.770 116.360 140.750 ;
        RECT 117.860 140.420 118.190 141.090 ;
        RECT 118.590 139.770 118.920 140.750 ;
        RECT 119.140 140.420 119.470 141.090 ;
        RECT 119.870 139.770 120.200 140.750 ;
        RECT 121.700 140.420 122.030 141.090 ;
        RECT 122.430 139.770 122.760 140.750 ;
        RECT 122.980 140.420 123.310 141.090 ;
        RECT 123.710 139.770 124.040 140.750 ;
        RECT 125.540 140.420 125.870 141.090 ;
        RECT 126.270 139.770 126.600 140.750 ;
        RECT 126.820 140.420 127.150 141.090 ;
        RECT 127.550 139.770 127.880 140.750 ;
        RECT 129.380 140.420 129.710 141.090 ;
        RECT 130.110 139.770 130.440 140.750 ;
        RECT 130.660 140.420 130.990 141.090 ;
        RECT 131.390 139.770 131.720 140.750 ;
        RECT 133.220 140.420 133.550 141.090 ;
        RECT 133.950 139.770 134.280 140.750 ;
        RECT 134.500 140.420 134.830 141.090 ;
        RECT 135.230 139.770 135.560 140.750 ;
        RECT 137.060 140.420 137.390 141.090 ;
        RECT 137.790 139.770 138.120 140.750 ;
        RECT 138.340 140.420 138.670 141.090 ;
        RECT 139.070 139.770 139.400 140.750 ;
        RECT 140.640 140.420 140.970 141.200 ;
        RECT 113.780 138.890 116.520 139.770 ;
        RECT 113.780 138.720 113.990 138.890 ;
        RECT 114.160 138.720 114.430 138.890 ;
        RECT 114.600 138.720 114.840 138.890 ;
        RECT 115.010 138.720 115.270 138.890 ;
        RECT 115.440 138.720 115.710 138.890 ;
        RECT 115.880 138.720 116.120 138.890 ;
        RECT 116.290 138.720 116.520 138.890 ;
        RECT 113.780 138.700 116.520 138.720 ;
        RECT 117.620 138.890 120.360 139.770 ;
        RECT 117.620 138.720 117.830 138.890 ;
        RECT 118.000 138.720 118.270 138.890 ;
        RECT 118.440 138.720 118.680 138.890 ;
        RECT 118.850 138.720 119.110 138.890 ;
        RECT 119.280 138.720 119.550 138.890 ;
        RECT 119.720 138.720 119.960 138.890 ;
        RECT 120.130 138.720 120.360 138.890 ;
        RECT 117.620 138.700 120.360 138.720 ;
        RECT 121.460 138.890 124.200 139.770 ;
        RECT 121.460 138.720 121.670 138.890 ;
        RECT 121.840 138.720 122.110 138.890 ;
        RECT 122.280 138.720 122.520 138.890 ;
        RECT 122.690 138.720 122.950 138.890 ;
        RECT 123.120 138.720 123.390 138.890 ;
        RECT 123.560 138.720 123.800 138.890 ;
        RECT 123.970 138.720 124.200 138.890 ;
        RECT 121.460 138.700 124.200 138.720 ;
        RECT 125.300 138.890 128.040 139.770 ;
        RECT 125.300 138.720 125.510 138.890 ;
        RECT 125.680 138.720 125.950 138.890 ;
        RECT 126.120 138.720 126.360 138.890 ;
        RECT 126.530 138.720 126.790 138.890 ;
        RECT 126.960 138.720 127.230 138.890 ;
        RECT 127.400 138.720 127.640 138.890 ;
        RECT 127.810 138.720 128.040 138.890 ;
        RECT 125.300 138.700 128.040 138.720 ;
        RECT 129.140 138.890 131.880 139.770 ;
        RECT 129.140 138.720 129.350 138.890 ;
        RECT 129.520 138.720 129.790 138.890 ;
        RECT 129.960 138.720 130.200 138.890 ;
        RECT 130.370 138.720 130.630 138.890 ;
        RECT 130.800 138.720 131.070 138.890 ;
        RECT 131.240 138.720 131.480 138.890 ;
        RECT 131.650 138.720 131.880 138.890 ;
        RECT 129.140 138.700 131.880 138.720 ;
        RECT 132.980 138.890 135.720 139.770 ;
        RECT 132.980 138.720 133.190 138.890 ;
        RECT 133.360 138.720 133.630 138.890 ;
        RECT 133.800 138.720 134.040 138.890 ;
        RECT 134.210 138.720 134.470 138.890 ;
        RECT 134.640 138.720 134.910 138.890 ;
        RECT 135.080 138.720 135.320 138.890 ;
        RECT 135.490 138.720 135.720 138.890 ;
        RECT 132.980 138.700 135.720 138.720 ;
        RECT 136.820 138.890 139.560 139.770 ;
        RECT 141.180 139.760 141.510 140.750 ;
        RECT 136.820 138.720 137.030 138.890 ;
        RECT 137.200 138.720 137.470 138.890 ;
        RECT 137.640 138.720 137.880 138.890 ;
        RECT 138.050 138.720 138.310 138.890 ;
        RECT 138.480 138.720 138.750 138.890 ;
        RECT 138.920 138.720 139.160 138.890 ;
        RECT 139.330 138.720 139.560 138.890 ;
        RECT 136.820 138.700 139.560 138.720 ;
        RECT 140.410 138.890 141.860 139.760 ;
        RECT 140.410 138.720 140.660 138.890 ;
        RECT 140.830 138.720 141.020 138.890 ;
        RECT 141.190 138.720 141.460 138.890 ;
        RECT 141.630 138.720 141.860 138.890 ;
        RECT 140.410 138.690 141.860 138.720 ;
        RECT 5.760 138.290 5.920 138.470 ;
        RECT 6.090 138.290 6.400 138.470 ;
        RECT 6.570 138.290 6.880 138.470 ;
        RECT 7.050 138.290 7.360 138.470 ;
        RECT 7.530 138.290 7.840 138.470 ;
        RECT 8.010 138.290 8.320 138.470 ;
        RECT 8.490 138.290 8.800 138.470 ;
        RECT 8.970 138.290 9.280 138.470 ;
        RECT 9.450 138.290 9.760 138.470 ;
        RECT 9.930 138.290 10.240 138.470 ;
        RECT 10.410 138.290 10.720 138.470 ;
        RECT 10.890 138.290 11.200 138.470 ;
        RECT 11.370 138.290 11.680 138.470 ;
        RECT 11.850 138.290 12.160 138.470 ;
        RECT 12.330 138.290 12.640 138.470 ;
        RECT 12.810 138.290 13.120 138.470 ;
        RECT 13.290 138.290 13.600 138.470 ;
        RECT 13.770 138.290 14.080 138.470 ;
        RECT 14.250 138.290 14.560 138.470 ;
        RECT 14.730 138.290 15.040 138.470 ;
        RECT 15.210 138.290 15.520 138.470 ;
        RECT 15.690 138.290 16.000 138.470 ;
        RECT 16.170 138.290 16.480 138.470 ;
        RECT 16.650 138.290 16.960 138.470 ;
        RECT 17.130 138.290 17.440 138.470 ;
        RECT 17.610 138.290 17.920 138.470 ;
        RECT 18.090 138.290 18.400 138.470 ;
        RECT 18.570 138.290 18.880 138.470 ;
        RECT 19.050 138.290 19.360 138.470 ;
        RECT 19.530 138.290 19.840 138.470 ;
        RECT 20.010 138.290 20.320 138.470 ;
        RECT 20.490 138.290 20.800 138.470 ;
        RECT 20.970 138.290 21.280 138.470 ;
        RECT 21.450 138.290 21.760 138.470 ;
        RECT 21.930 138.290 22.240 138.470 ;
        RECT 22.410 138.290 22.720 138.470 ;
        RECT 22.890 138.290 23.200 138.470 ;
        RECT 23.370 138.290 23.680 138.470 ;
        RECT 23.850 138.290 24.160 138.470 ;
        RECT 24.330 138.290 24.640 138.470 ;
        RECT 24.810 138.290 25.120 138.470 ;
        RECT 25.290 138.290 25.600 138.470 ;
        RECT 25.770 138.290 26.080 138.470 ;
        RECT 26.250 138.290 26.560 138.470 ;
        RECT 26.730 138.290 27.040 138.470 ;
        RECT 27.210 138.290 27.520 138.470 ;
        RECT 27.690 138.290 28.000 138.470 ;
        RECT 28.170 138.290 28.480 138.470 ;
        RECT 28.650 138.290 28.960 138.470 ;
        RECT 29.130 138.290 29.440 138.470 ;
        RECT 29.610 138.460 29.920 138.470 ;
        RECT 30.090 138.460 30.240 138.470 ;
        RECT 30.720 138.460 30.880 138.470 ;
        RECT 29.610 138.290 29.760 138.460 ;
        RECT 30.240 138.290 30.400 138.460 ;
        RECT 30.570 138.290 30.880 138.460 ;
        RECT 31.050 138.290 31.360 138.470 ;
        RECT 31.530 138.290 31.840 138.470 ;
        RECT 32.010 138.290 32.320 138.470 ;
        RECT 32.490 138.290 32.800 138.470 ;
        RECT 32.970 138.290 33.280 138.470 ;
        RECT 33.450 138.290 33.760 138.470 ;
        RECT 33.930 138.290 34.240 138.470 ;
        RECT 34.410 138.290 34.720 138.470 ;
        RECT 34.890 138.290 35.200 138.470 ;
        RECT 35.370 138.290 35.680 138.470 ;
        RECT 35.850 138.290 36.160 138.470 ;
        RECT 36.330 138.290 36.640 138.470 ;
        RECT 36.810 138.290 37.120 138.470 ;
        RECT 37.290 138.290 37.600 138.470 ;
        RECT 37.770 138.290 38.080 138.470 ;
        RECT 38.250 138.290 38.560 138.470 ;
        RECT 38.730 138.290 39.040 138.470 ;
        RECT 39.210 138.290 39.520 138.470 ;
        RECT 39.690 138.290 40.000 138.470 ;
        RECT 40.170 138.290 40.480 138.470 ;
        RECT 40.650 138.290 40.960 138.470 ;
        RECT 41.130 138.290 41.440 138.470 ;
        RECT 41.610 138.290 41.920 138.470 ;
        RECT 42.090 138.290 42.400 138.470 ;
        RECT 42.570 138.290 42.880 138.470 ;
        RECT 43.050 138.290 43.360 138.470 ;
        RECT 43.530 138.290 43.840 138.470 ;
        RECT 44.010 138.290 44.320 138.470 ;
        RECT 44.490 138.290 44.800 138.470 ;
        RECT 44.970 138.290 45.280 138.470 ;
        RECT 45.450 138.290 45.760 138.470 ;
        RECT 45.930 138.290 46.240 138.470 ;
        RECT 46.410 138.290 46.720 138.470 ;
        RECT 46.890 138.290 47.200 138.470 ;
        RECT 47.370 138.290 47.680 138.470 ;
        RECT 47.850 138.290 48.160 138.470 ;
        RECT 48.330 138.290 48.640 138.470 ;
        RECT 48.810 138.290 49.120 138.470 ;
        RECT 49.290 138.290 49.600 138.470 ;
        RECT 49.770 138.290 50.080 138.470 ;
        RECT 50.250 138.290 50.560 138.470 ;
        RECT 50.730 138.290 51.040 138.470 ;
        RECT 51.210 138.290 51.520 138.470 ;
        RECT 51.690 138.290 52.000 138.470 ;
        RECT 52.170 138.290 52.480 138.470 ;
        RECT 52.650 138.290 52.960 138.470 ;
        RECT 53.130 138.290 53.440 138.470 ;
        RECT 53.610 138.290 53.920 138.470 ;
        RECT 54.090 138.290 54.400 138.470 ;
        RECT 54.570 138.290 54.880 138.470 ;
        RECT 55.050 138.290 55.360 138.470 ;
        RECT 55.530 138.290 55.840 138.470 ;
        RECT 56.010 138.290 56.320 138.470 ;
        RECT 56.490 138.290 56.800 138.470 ;
        RECT 56.970 138.290 57.280 138.470 ;
        RECT 57.450 138.290 57.760 138.470 ;
        RECT 57.930 138.290 58.240 138.470 ;
        RECT 58.410 138.290 58.720 138.470 ;
        RECT 58.890 138.290 59.200 138.470 ;
        RECT 59.370 138.290 59.680 138.470 ;
        RECT 59.850 138.290 60.160 138.470 ;
        RECT 60.330 138.290 60.640 138.470 ;
        RECT 60.810 138.290 61.120 138.470 ;
        RECT 61.290 138.290 61.600 138.470 ;
        RECT 61.770 138.290 62.080 138.470 ;
        RECT 62.250 138.460 62.400 138.470 ;
        RECT 62.880 138.460 63.040 138.470 ;
        RECT 62.250 138.290 62.560 138.460 ;
        RECT 62.730 138.290 63.040 138.460 ;
        RECT 63.210 138.290 63.520 138.470 ;
        RECT 63.690 138.290 64.000 138.470 ;
        RECT 64.170 138.290 64.480 138.470 ;
        RECT 64.650 138.290 64.960 138.470 ;
        RECT 65.130 138.290 65.440 138.470 ;
        RECT 65.610 138.290 65.920 138.470 ;
        RECT 66.090 138.290 66.400 138.470 ;
        RECT 66.570 138.290 66.880 138.470 ;
        RECT 67.050 138.290 67.360 138.470 ;
        RECT 67.530 138.290 67.840 138.470 ;
        RECT 68.010 138.290 68.320 138.470 ;
        RECT 68.490 138.290 68.800 138.470 ;
        RECT 68.970 138.290 69.280 138.470 ;
        RECT 69.450 138.290 69.760 138.470 ;
        RECT 69.930 138.290 70.240 138.470 ;
        RECT 70.410 138.290 70.720 138.470 ;
        RECT 70.890 138.290 71.200 138.470 ;
        RECT 71.370 138.290 71.680 138.470 ;
        RECT 71.850 138.290 72.160 138.470 ;
        RECT 72.330 138.290 72.640 138.470 ;
        RECT 72.810 138.290 73.120 138.470 ;
        RECT 73.290 138.290 73.600 138.470 ;
        RECT 73.770 138.290 74.080 138.470 ;
        RECT 74.250 138.290 74.560 138.470 ;
        RECT 74.730 138.460 74.880 138.470 ;
        RECT 75.360 138.460 75.520 138.470 ;
        RECT 74.730 138.290 75.040 138.460 ;
        RECT 75.210 138.290 75.520 138.460 ;
        RECT 75.690 138.290 76.000 138.470 ;
        RECT 76.170 138.290 76.480 138.470 ;
        RECT 76.650 138.290 76.960 138.470 ;
        RECT 77.130 138.290 77.440 138.470 ;
        RECT 77.610 138.290 77.920 138.470 ;
        RECT 78.090 138.290 78.400 138.470 ;
        RECT 78.570 138.290 78.880 138.470 ;
        RECT 79.050 138.290 79.360 138.470 ;
        RECT 79.530 138.290 79.840 138.470 ;
        RECT 80.010 138.290 80.320 138.470 ;
        RECT 80.490 138.290 80.800 138.470 ;
        RECT 80.970 138.290 81.280 138.470 ;
        RECT 81.450 138.290 81.760 138.470 ;
        RECT 81.930 138.290 82.240 138.470 ;
        RECT 82.410 138.290 82.720 138.470 ;
        RECT 82.890 138.290 83.200 138.470 ;
        RECT 83.370 138.290 83.680 138.470 ;
        RECT 83.850 138.290 84.160 138.470 ;
        RECT 84.330 138.290 84.640 138.470 ;
        RECT 84.810 138.290 85.120 138.470 ;
        RECT 85.290 138.290 85.600 138.470 ;
        RECT 85.770 138.290 86.080 138.470 ;
        RECT 86.250 138.290 86.560 138.470 ;
        RECT 86.730 138.290 87.040 138.470 ;
        RECT 87.210 138.290 87.520 138.470 ;
        RECT 87.690 138.290 88.000 138.470 ;
        RECT 88.170 138.290 88.480 138.470 ;
        RECT 88.650 138.290 88.960 138.470 ;
        RECT 89.130 138.290 89.440 138.470 ;
        RECT 89.610 138.290 89.920 138.470 ;
        RECT 90.090 138.290 90.400 138.470 ;
        RECT 90.570 138.290 90.880 138.470 ;
        RECT 91.050 138.290 91.360 138.470 ;
        RECT 91.530 138.290 91.840 138.470 ;
        RECT 92.010 138.290 92.320 138.470 ;
        RECT 92.490 138.290 92.800 138.470 ;
        RECT 92.970 138.290 93.280 138.470 ;
        RECT 93.450 138.290 93.760 138.470 ;
        RECT 93.930 138.290 94.240 138.470 ;
        RECT 94.410 138.290 94.720 138.470 ;
        RECT 94.890 138.290 95.200 138.470 ;
        RECT 95.370 138.290 95.680 138.470 ;
        RECT 95.850 138.290 96.160 138.470 ;
        RECT 96.330 138.290 96.640 138.470 ;
        RECT 96.810 138.290 97.120 138.470 ;
        RECT 97.290 138.290 97.600 138.470 ;
        RECT 97.770 138.460 97.920 138.470 ;
        RECT 98.400 138.460 98.560 138.470 ;
        RECT 97.770 138.290 98.080 138.460 ;
        RECT 98.250 138.290 98.560 138.460 ;
        RECT 98.730 138.290 99.040 138.470 ;
        RECT 99.210 138.290 99.520 138.470 ;
        RECT 99.690 138.290 100.000 138.470 ;
        RECT 100.170 138.290 100.480 138.470 ;
        RECT 100.650 138.290 100.960 138.470 ;
        RECT 101.130 138.290 101.440 138.470 ;
        RECT 101.610 138.290 101.920 138.470 ;
        RECT 102.090 138.290 102.400 138.470 ;
        RECT 102.570 138.290 102.880 138.470 ;
        RECT 103.050 138.290 103.360 138.470 ;
        RECT 103.530 138.290 103.840 138.470 ;
        RECT 104.010 138.290 104.320 138.470 ;
        RECT 104.490 138.290 104.800 138.470 ;
        RECT 104.970 138.290 105.280 138.470 ;
        RECT 105.450 138.290 105.760 138.470 ;
        RECT 105.930 138.290 106.240 138.470 ;
        RECT 106.410 138.290 106.720 138.470 ;
        RECT 106.890 138.290 107.200 138.470 ;
        RECT 107.370 138.290 107.680 138.470 ;
        RECT 107.850 138.290 108.160 138.470 ;
        RECT 108.330 138.290 108.640 138.470 ;
        RECT 108.810 138.290 109.120 138.470 ;
        RECT 109.290 138.460 109.440 138.470 ;
        RECT 109.920 138.460 110.080 138.470 ;
        RECT 109.290 138.290 109.600 138.460 ;
        RECT 109.770 138.290 110.080 138.460 ;
        RECT 110.250 138.290 110.560 138.470 ;
        RECT 110.730 138.290 111.040 138.470 ;
        RECT 111.210 138.290 111.520 138.470 ;
        RECT 111.690 138.290 112.000 138.470 ;
        RECT 112.170 138.290 112.480 138.470 ;
        RECT 112.650 138.290 112.960 138.470 ;
        RECT 113.130 138.290 113.440 138.470 ;
        RECT 113.610 138.290 113.920 138.470 ;
        RECT 114.090 138.290 114.400 138.470 ;
        RECT 114.570 138.290 114.880 138.470 ;
        RECT 115.050 138.290 115.360 138.470 ;
        RECT 115.530 138.290 115.840 138.470 ;
        RECT 116.010 138.290 116.320 138.470 ;
        RECT 116.490 138.290 116.800 138.470 ;
        RECT 116.970 138.290 117.280 138.470 ;
        RECT 117.450 138.290 117.760 138.470 ;
        RECT 117.930 138.290 118.240 138.470 ;
        RECT 118.410 138.290 118.720 138.470 ;
        RECT 118.890 138.290 119.200 138.470 ;
        RECT 119.370 138.290 119.680 138.470 ;
        RECT 119.850 138.290 120.160 138.470 ;
        RECT 120.330 138.290 120.640 138.470 ;
        RECT 120.810 138.290 121.120 138.470 ;
        RECT 121.290 138.290 121.600 138.470 ;
        RECT 121.770 138.290 122.080 138.470 ;
        RECT 122.250 138.290 122.560 138.470 ;
        RECT 122.730 138.290 123.040 138.470 ;
        RECT 123.210 138.290 123.520 138.470 ;
        RECT 123.690 138.290 124.000 138.470 ;
        RECT 124.170 138.290 124.480 138.470 ;
        RECT 124.650 138.290 124.960 138.470 ;
        RECT 125.130 138.290 125.440 138.470 ;
        RECT 125.610 138.290 125.920 138.470 ;
        RECT 126.090 138.290 126.400 138.470 ;
        RECT 126.570 138.290 126.880 138.470 ;
        RECT 127.050 138.290 127.360 138.470 ;
        RECT 127.530 138.290 127.840 138.470 ;
        RECT 128.010 138.290 128.320 138.470 ;
        RECT 128.490 138.290 128.800 138.470 ;
        RECT 128.970 138.290 129.280 138.470 ;
        RECT 129.450 138.290 129.760 138.470 ;
        RECT 129.930 138.290 130.240 138.470 ;
        RECT 130.410 138.290 130.720 138.470 ;
        RECT 130.890 138.290 131.200 138.470 ;
        RECT 131.370 138.290 131.680 138.470 ;
        RECT 131.850 138.290 132.160 138.470 ;
        RECT 132.330 138.290 132.640 138.470 ;
        RECT 132.810 138.290 133.120 138.470 ;
        RECT 133.290 138.290 133.600 138.470 ;
        RECT 133.770 138.290 134.080 138.470 ;
        RECT 134.250 138.290 134.560 138.470 ;
        RECT 134.730 138.290 135.040 138.470 ;
        RECT 135.210 138.290 135.520 138.470 ;
        RECT 135.690 138.290 136.000 138.470 ;
        RECT 136.170 138.290 136.480 138.470 ;
        RECT 136.650 138.290 136.960 138.470 ;
        RECT 137.130 138.290 137.440 138.470 ;
        RECT 137.610 138.290 137.920 138.470 ;
        RECT 138.090 138.290 138.400 138.470 ;
        RECT 138.570 138.290 138.880 138.470 ;
        RECT 139.050 138.290 139.360 138.470 ;
        RECT 139.530 138.290 139.840 138.470 ;
        RECT 140.010 138.290 140.320 138.470 ;
        RECT 140.490 138.290 140.800 138.470 ;
        RECT 140.970 138.290 141.280 138.470 ;
        RECT 141.450 138.460 141.600 138.470 ;
        RECT 141.450 138.290 141.760 138.460 ;
        RECT 141.930 138.290 142.080 138.460 ;
        RECT 6.260 138.040 9.000 138.060 ;
        RECT 6.260 137.870 6.470 138.040 ;
        RECT 6.640 137.870 6.910 138.040 ;
        RECT 7.080 137.870 7.320 138.040 ;
        RECT 7.490 137.870 7.750 138.040 ;
        RECT 7.920 137.870 8.190 138.040 ;
        RECT 8.360 137.870 8.600 138.040 ;
        RECT 8.770 137.870 9.000 138.040 ;
        RECT 6.260 136.990 9.000 137.870 ;
        RECT 9.850 138.040 11.300 138.070 ;
        RECT 9.850 137.870 10.100 138.040 ;
        RECT 10.270 137.870 10.460 138.040 ;
        RECT 10.630 137.870 10.900 138.040 ;
        RECT 11.070 137.870 11.300 138.040 ;
        RECT 9.850 137.000 11.300 137.870 ;
        RECT 13.210 137.990 13.770 138.070 ;
        RECT 13.210 137.820 13.220 137.990 ;
        RECT 13.390 137.820 13.580 137.990 ;
        RECT 13.750 137.820 13.770 137.990 ;
        RECT 6.500 135.670 6.830 136.340 ;
        RECT 7.230 136.010 7.560 136.990 ;
        RECT 7.780 135.670 8.110 136.340 ;
        RECT 8.510 136.010 8.840 136.990 ;
        RECT 6.340 134.670 9.070 135.670 ;
        RECT 10.080 135.560 10.410 136.340 ;
        RECT 10.620 136.010 10.950 137.000 ;
        RECT 13.210 136.490 13.770 137.820 ;
        RECT 15.380 138.040 18.120 138.060 ;
        RECT 15.380 137.870 15.590 138.040 ;
        RECT 15.760 137.870 16.030 138.040 ;
        RECT 16.200 137.870 16.440 138.040 ;
        RECT 16.610 137.870 16.870 138.040 ;
        RECT 17.040 137.870 17.310 138.040 ;
        RECT 17.480 137.870 17.720 138.040 ;
        RECT 17.890 137.870 18.120 138.040 ;
        RECT 13.160 135.600 13.490 136.060 ;
        RECT 14.460 135.600 14.710 137.320 ;
        RECT 15.380 136.990 18.120 137.870 ;
        RECT 19.220 138.040 21.960 138.060 ;
        RECT 19.220 137.870 19.430 138.040 ;
        RECT 19.600 137.870 19.870 138.040 ;
        RECT 20.040 137.870 20.280 138.040 ;
        RECT 20.450 137.870 20.710 138.040 ;
        RECT 20.880 137.870 21.150 138.040 ;
        RECT 21.320 137.870 21.560 138.040 ;
        RECT 21.730 137.870 21.960 138.040 ;
        RECT 19.220 136.990 21.960 137.870 ;
        RECT 23.060 138.040 25.800 138.060 ;
        RECT 23.060 137.870 23.270 138.040 ;
        RECT 23.440 137.870 23.710 138.040 ;
        RECT 23.880 137.870 24.120 138.040 ;
        RECT 24.290 137.870 24.550 138.040 ;
        RECT 24.720 137.870 24.990 138.040 ;
        RECT 25.160 137.870 25.400 138.040 ;
        RECT 25.570 137.870 25.800 138.040 ;
        RECT 23.060 136.990 25.800 137.870 ;
        RECT 26.900 138.040 29.640 138.060 ;
        RECT 26.900 137.870 27.110 138.040 ;
        RECT 27.280 137.870 27.550 138.040 ;
        RECT 27.720 137.870 27.960 138.040 ;
        RECT 28.130 137.870 28.390 138.040 ;
        RECT 28.560 137.870 28.830 138.040 ;
        RECT 29.000 137.870 29.240 138.040 ;
        RECT 29.410 137.870 29.640 138.040 ;
        RECT 26.900 136.990 29.640 137.870 ;
        RECT 15.620 135.670 15.950 136.340 ;
        RECT 16.350 136.010 16.680 136.990 ;
        RECT 16.900 135.670 17.230 136.340 ;
        RECT 17.630 136.010 17.960 136.990 ;
        RECT 19.460 135.670 19.790 136.340 ;
        RECT 20.190 136.010 20.520 136.990 ;
        RECT 20.740 135.670 21.070 136.340 ;
        RECT 21.470 136.010 21.800 136.990 ;
        RECT 23.300 135.670 23.630 136.340 ;
        RECT 24.030 136.010 24.360 136.990 ;
        RECT 24.580 135.670 24.910 136.340 ;
        RECT 25.310 136.010 25.640 136.990 ;
        RECT 27.140 135.670 27.470 136.340 ;
        RECT 27.870 136.010 28.200 136.990 ;
        RECT 28.420 135.670 28.750 136.340 ;
        RECT 29.150 136.010 29.480 136.990 ;
      LAYER li1 ;
        RECT 30.840 136.490 31.270 138.070 ;
      LAYER li1 ;
        RECT 31.450 137.990 32.010 138.070 ;
        RECT 31.450 137.820 31.460 137.990 ;
        RECT 31.630 137.820 31.820 137.990 ;
        RECT 31.990 137.820 32.010 137.990 ;
        RECT 31.450 136.490 32.010 137.820 ;
        RECT 33.370 138.040 34.820 138.070 ;
        RECT 33.370 137.870 33.620 138.040 ;
        RECT 33.790 137.870 33.980 138.040 ;
        RECT 34.150 137.870 34.420 138.040 ;
        RECT 34.590 137.870 34.820 138.040 ;
        RECT 10.080 135.160 11.380 135.560 ;
        RECT 13.160 135.430 14.710 135.600 ;
        RECT 9.770 134.680 11.380 135.160 ;
        RECT 13.030 134.680 14.280 135.250 ;
        RECT 14.460 134.810 14.710 135.430 ;
        RECT 15.460 134.670 18.190 135.670 ;
        RECT 19.300 134.670 22.030 135.670 ;
        RECT 23.140 134.670 25.870 135.670 ;
        RECT 26.980 134.670 29.710 135.670 ;
      LAYER li1 ;
        RECT 30.840 134.810 31.090 136.490 ;
      LAYER li1 ;
        RECT 31.400 135.600 31.730 136.060 ;
      LAYER li1 ;
        RECT 32.190 135.780 32.520 137.570 ;
      LAYER li1 ;
        RECT 32.700 135.600 32.950 137.320 ;
        RECT 33.370 137.000 34.820 137.870 ;
        RECT 35.130 137.990 35.720 138.070 ;
        RECT 35.130 137.820 35.160 137.990 ;
        RECT 35.330 137.820 35.520 137.990 ;
        RECT 35.690 137.820 35.720 137.990 ;
        RECT 31.400 135.430 32.950 135.600 ;
        RECT 31.270 134.680 32.520 135.250 ;
        RECT 32.700 134.810 32.950 135.430 ;
        RECT 33.600 135.560 33.930 136.340 ;
        RECT 34.140 136.010 34.470 137.000 ;
        RECT 35.130 136.490 35.720 137.820 ;
      LAYER li1 ;
        RECT 36.000 136.490 36.390 138.070 ;
      LAYER li1 ;
        RECT 36.980 138.040 39.720 138.060 ;
        RECT 36.980 137.870 37.190 138.040 ;
        RECT 37.360 137.870 37.630 138.040 ;
        RECT 37.800 137.870 38.040 138.040 ;
        RECT 38.210 137.870 38.470 138.040 ;
        RECT 38.640 137.870 38.910 138.040 ;
        RECT 39.080 137.870 39.320 138.040 ;
        RECT 39.490 137.870 39.720 138.040 ;
        RECT 36.980 136.990 39.720 137.870 ;
        RECT 40.820 138.040 43.560 138.060 ;
        RECT 40.820 137.870 41.030 138.040 ;
        RECT 41.200 137.870 41.470 138.040 ;
        RECT 41.640 137.870 41.880 138.040 ;
        RECT 42.050 137.870 42.310 138.040 ;
        RECT 42.480 137.870 42.750 138.040 ;
        RECT 42.920 137.870 43.160 138.040 ;
        RECT 43.330 137.870 43.560 138.040 ;
        RECT 40.820 136.990 43.560 137.870 ;
        RECT 44.660 138.040 47.400 138.060 ;
        RECT 44.660 137.870 44.870 138.040 ;
        RECT 45.040 137.870 45.310 138.040 ;
        RECT 45.480 137.870 45.720 138.040 ;
        RECT 45.890 137.870 46.150 138.040 ;
        RECT 46.320 137.870 46.590 138.040 ;
        RECT 46.760 137.870 47.000 138.040 ;
        RECT 47.170 137.870 47.400 138.040 ;
        RECT 44.660 136.990 47.400 137.870 ;
        RECT 48.500 138.040 51.240 138.060 ;
        RECT 48.500 137.870 48.710 138.040 ;
        RECT 48.880 137.870 49.150 138.040 ;
        RECT 49.320 137.870 49.560 138.040 ;
        RECT 49.730 137.870 49.990 138.040 ;
        RECT 50.160 137.870 50.430 138.040 ;
        RECT 50.600 137.870 50.840 138.040 ;
        RECT 51.010 137.870 51.240 138.040 ;
        RECT 48.500 136.990 51.240 137.870 ;
        RECT 52.340 138.040 55.080 138.060 ;
        RECT 52.340 137.870 52.550 138.040 ;
        RECT 52.720 137.870 52.990 138.040 ;
        RECT 53.160 137.870 53.400 138.040 ;
        RECT 53.570 137.870 53.830 138.040 ;
        RECT 54.000 137.870 54.270 138.040 ;
        RECT 54.440 137.870 54.680 138.040 ;
        RECT 54.850 137.870 55.080 138.040 ;
        RECT 52.340 136.990 55.080 137.870 ;
        RECT 56.180 138.040 58.920 138.060 ;
        RECT 56.180 137.870 56.390 138.040 ;
        RECT 56.560 137.870 56.830 138.040 ;
        RECT 57.000 137.870 57.240 138.040 ;
        RECT 57.410 137.870 57.670 138.040 ;
        RECT 57.840 137.870 58.110 138.040 ;
        RECT 58.280 137.870 58.520 138.040 ;
        RECT 58.690 137.870 58.920 138.040 ;
        RECT 56.180 136.990 58.920 137.870 ;
        RECT 59.770 138.040 61.220 138.070 ;
        RECT 59.770 137.870 60.020 138.040 ;
        RECT 60.190 137.870 60.380 138.040 ;
        RECT 60.550 137.870 60.820 138.040 ;
        RECT 60.990 137.870 61.220 138.040 ;
        RECT 59.770 137.000 61.220 137.870 ;
        RECT 62.970 137.990 63.560 138.070 ;
        RECT 62.970 137.820 63.000 137.990 ;
        RECT 63.170 137.820 63.360 137.990 ;
        RECT 63.530 137.820 63.560 137.990 ;
        RECT 33.600 135.160 34.900 135.560 ;
        RECT 33.290 134.680 34.900 135.160 ;
        RECT 35.130 134.680 35.720 135.640 ;
      LAYER li1 ;
        RECT 36.060 134.810 36.390 136.490 ;
      LAYER li1 ;
        RECT 37.220 135.670 37.550 136.340 ;
        RECT 37.950 136.010 38.280 136.990 ;
        RECT 38.500 135.670 38.830 136.340 ;
        RECT 39.230 136.010 39.560 136.990 ;
        RECT 41.060 135.670 41.390 136.340 ;
        RECT 41.790 136.010 42.120 136.990 ;
        RECT 42.340 135.670 42.670 136.340 ;
        RECT 43.070 136.010 43.400 136.990 ;
        RECT 44.900 135.670 45.230 136.340 ;
        RECT 45.630 136.010 45.960 136.990 ;
        RECT 46.180 135.670 46.510 136.340 ;
        RECT 46.910 136.010 47.240 136.990 ;
        RECT 48.740 135.670 49.070 136.340 ;
        RECT 49.470 136.010 49.800 136.990 ;
        RECT 50.020 135.670 50.350 136.340 ;
        RECT 50.750 136.010 51.080 136.990 ;
        RECT 52.580 135.670 52.910 136.340 ;
        RECT 53.310 136.010 53.640 136.990 ;
        RECT 53.860 135.670 54.190 136.340 ;
        RECT 54.590 136.010 54.920 136.990 ;
        RECT 56.420 135.670 56.750 136.340 ;
        RECT 57.150 136.010 57.480 136.990 ;
        RECT 57.700 135.670 58.030 136.340 ;
        RECT 58.430 136.010 58.760 136.990 ;
        RECT 37.060 134.670 39.790 135.670 ;
        RECT 40.900 134.670 43.630 135.670 ;
        RECT 44.740 134.670 47.470 135.670 ;
        RECT 48.580 134.670 51.310 135.670 ;
        RECT 52.420 134.670 55.150 135.670 ;
        RECT 56.260 134.670 58.990 135.670 ;
        RECT 60.000 135.560 60.330 136.340 ;
        RECT 60.540 136.010 60.870 137.000 ;
        RECT 62.970 136.490 63.560 137.820 ;
      LAYER li1 ;
        RECT 63.840 136.490 64.230 138.070 ;
      LAYER li1 ;
        RECT 64.820 138.040 67.560 138.060 ;
        RECT 64.820 137.870 65.030 138.040 ;
        RECT 65.200 137.870 65.470 138.040 ;
        RECT 65.640 137.870 65.880 138.040 ;
        RECT 66.050 137.870 66.310 138.040 ;
        RECT 66.480 137.870 66.750 138.040 ;
        RECT 66.920 137.870 67.160 138.040 ;
        RECT 67.330 137.870 67.560 138.040 ;
        RECT 64.820 136.990 67.560 137.870 ;
        RECT 68.660 138.040 71.400 138.060 ;
        RECT 68.660 137.870 68.870 138.040 ;
        RECT 69.040 137.870 69.310 138.040 ;
        RECT 69.480 137.870 69.720 138.040 ;
        RECT 69.890 137.870 70.150 138.040 ;
        RECT 70.320 137.870 70.590 138.040 ;
        RECT 70.760 137.870 71.000 138.040 ;
        RECT 71.170 137.870 71.400 138.040 ;
        RECT 68.660 136.990 71.400 137.870 ;
        RECT 72.250 138.040 73.700 138.070 ;
        RECT 72.250 137.870 72.500 138.040 ;
        RECT 72.670 137.870 72.860 138.040 ;
        RECT 73.030 137.870 73.300 138.040 ;
        RECT 73.470 137.870 73.700 138.040 ;
        RECT 72.250 137.000 73.700 137.870 ;
        RECT 75.450 137.990 76.710 138.070 ;
        RECT 75.450 137.820 75.460 137.990 ;
        RECT 75.630 137.820 75.820 137.990 ;
        RECT 75.990 137.820 76.180 137.990 ;
        RECT 76.350 137.820 76.540 137.990 ;
        RECT 60.000 135.160 61.300 135.560 ;
        RECT 59.690 134.680 61.300 135.160 ;
        RECT 62.970 134.680 63.560 135.640 ;
      LAYER li1 ;
        RECT 63.900 134.810 64.230 136.490 ;
      LAYER li1 ;
        RECT 65.060 135.670 65.390 136.340 ;
        RECT 65.790 136.010 66.120 136.990 ;
        RECT 66.340 135.670 66.670 136.340 ;
        RECT 67.070 136.010 67.400 136.990 ;
        RECT 68.900 135.670 69.230 136.340 ;
        RECT 69.630 136.010 69.960 136.990 ;
        RECT 70.180 135.670 70.510 136.340 ;
        RECT 70.910 136.010 71.240 136.990 ;
        RECT 64.900 134.670 67.630 135.670 ;
        RECT 68.740 134.670 71.470 135.670 ;
        RECT 72.480 135.560 72.810 136.340 ;
        RECT 73.020 136.010 73.350 137.000 ;
        RECT 75.450 136.590 76.710 137.820 ;
      LAYER li1 ;
        RECT 77.240 137.570 77.410 138.070 ;
        RECT 76.890 136.490 77.410 137.570 ;
      LAYER li1 ;
        RECT 77.670 137.990 78.980 138.070 ;
        RECT 77.670 137.820 77.700 137.990 ;
        RECT 77.870 137.820 78.060 137.990 ;
        RECT 78.230 137.820 78.420 137.990 ;
        RECT 78.590 137.820 78.780 137.990 ;
        RECT 78.950 137.820 78.980 137.990 ;
        RECT 77.670 136.610 78.980 137.820 ;
        RECT 79.700 138.040 82.440 138.060 ;
        RECT 79.700 137.870 79.910 138.040 ;
        RECT 80.080 137.870 80.350 138.040 ;
        RECT 80.520 137.870 80.760 138.040 ;
        RECT 80.930 137.870 81.190 138.040 ;
        RECT 81.360 137.870 81.630 138.040 ;
        RECT 81.800 137.870 82.040 138.040 ;
        RECT 82.210 137.870 82.440 138.040 ;
        RECT 79.700 136.990 82.440 137.870 ;
        RECT 83.540 138.040 86.280 138.060 ;
        RECT 83.540 137.870 83.750 138.040 ;
        RECT 83.920 137.870 84.190 138.040 ;
        RECT 84.360 137.870 84.600 138.040 ;
        RECT 84.770 137.870 85.030 138.040 ;
        RECT 85.200 137.870 85.470 138.040 ;
        RECT 85.640 137.870 85.880 138.040 ;
        RECT 86.050 137.870 86.280 138.040 ;
        RECT 83.540 136.990 86.280 137.870 ;
      LAYER li1 ;
        RECT 76.890 136.410 77.160 136.490 ;
        RECT 76.100 136.240 77.160 136.410 ;
        RECT 75.490 135.850 75.910 136.180 ;
        RECT 76.100 135.670 76.270 136.240 ;
        RECT 77.610 136.120 78.120 136.430 ;
        RECT 78.370 136.120 79.080 136.430 ;
        RECT 76.450 135.850 76.960 136.060 ;
      LAYER li1 ;
        RECT 77.160 135.770 79.030 135.940 ;
        RECT 72.480 135.160 73.780 135.560 ;
        RECT 72.170 134.680 73.780 135.160 ;
        RECT 75.520 134.750 75.850 135.670 ;
      LAYER li1 ;
        RECT 76.100 134.930 76.630 135.670 ;
      LAYER li1 ;
        RECT 77.160 134.750 77.330 135.770 ;
        RECT 75.520 134.580 77.330 134.750 ;
        RECT 77.510 134.680 78.610 135.590 ;
        RECT 78.780 134.840 79.030 135.770 ;
        RECT 79.940 135.670 80.270 136.340 ;
        RECT 80.670 136.010 81.000 136.990 ;
        RECT 81.220 135.670 81.550 136.340 ;
        RECT 81.950 136.010 82.280 136.990 ;
        RECT 83.780 135.670 84.110 136.340 ;
        RECT 84.510 136.010 84.840 136.990 ;
        RECT 85.060 135.670 85.390 136.340 ;
        RECT 85.790 136.010 86.120 136.990 ;
        RECT 79.780 134.670 82.510 135.670 ;
        RECT 83.620 134.670 86.350 135.670 ;
      LAYER li1 ;
        RECT 87.010 134.810 87.260 138.070 ;
      LAYER li1 ;
        RECT 87.440 137.990 90.130 138.070 ;
        RECT 87.610 137.820 87.800 137.990 ;
        RECT 87.970 137.820 88.160 137.990 ;
        RECT 88.330 137.820 88.520 137.990 ;
        RECT 88.690 137.820 88.880 137.990 ;
        RECT 89.050 137.820 89.240 137.990 ;
        RECT 89.410 137.820 89.600 137.990 ;
        RECT 89.770 137.820 89.960 137.990 ;
        RECT 87.440 136.960 90.130 137.820 ;
        RECT 90.310 136.780 90.560 138.070 ;
        RECT 87.470 136.610 90.560 136.780 ;
        RECT 87.470 135.910 87.800 136.610 ;
        RECT 90.310 136.490 90.560 136.610 ;
        RECT 90.740 137.990 92.050 138.050 ;
        RECT 90.740 137.820 90.770 137.990 ;
        RECT 90.940 137.820 91.130 137.990 ;
        RECT 91.300 137.820 91.490 137.990 ;
        RECT 91.660 137.820 91.850 137.990 ;
        RECT 92.020 137.820 92.050 137.990 ;
        RECT 90.740 136.510 92.050 137.820 ;
        RECT 92.660 138.040 95.400 138.060 ;
        RECT 92.660 137.870 92.870 138.040 ;
        RECT 93.040 137.870 93.310 138.040 ;
        RECT 93.480 137.870 93.720 138.040 ;
        RECT 93.890 137.870 94.150 138.040 ;
        RECT 94.320 137.870 94.590 138.040 ;
        RECT 94.760 137.870 95.000 138.040 ;
        RECT 95.170 137.870 95.400 138.040 ;
        RECT 92.660 136.990 95.400 137.870 ;
        RECT 96.250 138.040 97.700 138.070 ;
        RECT 96.250 137.870 96.500 138.040 ;
        RECT 96.670 137.870 96.860 138.040 ;
        RECT 97.030 137.870 97.300 138.040 ;
        RECT 97.470 137.870 97.700 138.040 ;
        RECT 96.250 137.000 97.700 137.870 ;
      LAYER li1 ;
        RECT 88.300 136.090 89.030 136.370 ;
      LAYER li1 ;
        RECT 87.470 135.740 88.680 135.910 ;
        RECT 87.440 134.680 88.330 135.560 ;
        RECT 88.510 135.530 88.680 135.740 ;
      LAYER li1 ;
        RECT 88.860 135.880 89.030 136.090 ;
        RECT 89.210 136.060 89.640 136.430 ;
        RECT 89.840 135.890 90.130 136.430 ;
        RECT 90.370 135.890 91.080 136.220 ;
        RECT 88.860 135.710 89.660 135.880 ;
        RECT 91.430 135.710 91.760 136.330 ;
        RECT 89.490 135.540 91.760 135.710 ;
      LAYER li1 ;
        RECT 92.900 135.670 93.230 136.340 ;
        RECT 93.630 136.010 93.960 136.990 ;
        RECT 94.180 135.670 94.510 136.340 ;
        RECT 94.910 136.010 95.240 136.990 ;
        RECT 88.510 135.360 89.310 135.530 ;
      LAYER li1 ;
        RECT 89.920 135.520 90.590 135.540 ;
      LAYER li1 ;
        RECT 89.140 135.190 89.740 135.360 ;
        RECT 88.630 134.750 88.960 135.180 ;
        RECT 89.410 134.930 89.740 135.190 ;
        RECT 90.230 134.750 90.560 135.340 ;
        RECT 88.630 134.580 90.560 134.750 ;
        RECT 90.770 134.680 92.070 135.360 ;
        RECT 92.740 134.670 95.470 135.670 ;
        RECT 96.480 135.560 96.810 136.340 ;
        RECT 97.020 136.010 97.350 137.000 ;
        RECT 96.480 135.160 97.780 135.560 ;
        RECT 96.170 134.680 97.780 135.160 ;
      LAYER li1 ;
        RECT 98.530 134.810 98.780 138.070 ;
      LAYER li1 ;
        RECT 98.960 137.990 101.650 138.070 ;
        RECT 99.130 137.820 99.320 137.990 ;
        RECT 99.490 137.820 99.680 137.990 ;
        RECT 99.850 137.820 100.040 137.990 ;
        RECT 100.210 137.820 100.400 137.990 ;
        RECT 100.570 137.820 100.760 137.990 ;
        RECT 100.930 137.820 101.120 137.990 ;
        RECT 101.290 137.820 101.480 137.990 ;
        RECT 98.960 136.960 101.650 137.820 ;
        RECT 101.830 136.780 102.080 138.070 ;
        RECT 98.990 136.610 102.080 136.780 ;
        RECT 98.990 135.910 99.320 136.610 ;
        RECT 101.830 136.490 102.080 136.610 ;
        RECT 102.260 137.990 103.570 138.050 ;
        RECT 102.260 137.820 102.290 137.990 ;
        RECT 102.460 137.820 102.650 137.990 ;
        RECT 102.820 137.820 103.010 137.990 ;
        RECT 103.180 137.820 103.370 137.990 ;
        RECT 103.540 137.820 103.570 137.990 ;
        RECT 102.260 136.510 103.570 137.820 ;
        RECT 104.180 138.040 106.920 138.060 ;
        RECT 104.180 137.870 104.390 138.040 ;
        RECT 104.560 137.870 104.830 138.040 ;
        RECT 105.000 137.870 105.240 138.040 ;
        RECT 105.410 137.870 105.670 138.040 ;
        RECT 105.840 137.870 106.110 138.040 ;
        RECT 106.280 137.870 106.520 138.040 ;
        RECT 106.690 137.870 106.920 138.040 ;
        RECT 104.180 136.990 106.920 137.870 ;
        RECT 107.770 138.040 109.220 138.070 ;
        RECT 107.770 137.870 108.020 138.040 ;
        RECT 108.190 137.870 108.380 138.040 ;
        RECT 108.550 137.870 108.820 138.040 ;
        RECT 108.990 137.870 109.220 138.040 ;
        RECT 107.770 137.000 109.220 137.870 ;
      LAYER li1 ;
        RECT 99.820 136.090 100.550 136.370 ;
      LAYER li1 ;
        RECT 98.990 135.740 100.200 135.910 ;
        RECT 98.960 134.680 99.850 135.560 ;
        RECT 100.030 135.530 100.200 135.740 ;
      LAYER li1 ;
        RECT 100.380 135.880 100.550 136.090 ;
        RECT 100.730 136.060 101.160 136.430 ;
        RECT 101.360 135.890 101.650 136.430 ;
        RECT 101.890 135.890 102.600 136.220 ;
        RECT 100.380 135.710 101.180 135.880 ;
        RECT 102.950 135.710 103.280 136.330 ;
        RECT 101.010 135.540 103.280 135.710 ;
      LAYER li1 ;
        RECT 104.420 135.670 104.750 136.340 ;
        RECT 105.150 136.010 105.480 136.990 ;
        RECT 105.700 135.670 106.030 136.340 ;
        RECT 106.430 136.010 106.760 136.990 ;
        RECT 100.030 135.360 100.830 135.530 ;
      LAYER li1 ;
        RECT 101.430 135.520 102.110 135.540 ;
      LAYER li1 ;
        RECT 100.660 135.190 101.260 135.360 ;
        RECT 100.150 134.750 100.480 135.180 ;
        RECT 100.930 134.930 101.260 135.190 ;
        RECT 101.750 134.750 102.080 135.340 ;
        RECT 100.150 134.580 102.080 134.750 ;
        RECT 102.290 134.680 103.590 135.360 ;
        RECT 104.260 134.670 106.990 135.670 ;
        RECT 108.000 135.560 108.330 136.340 ;
        RECT 108.540 136.010 108.870 137.000 ;
      LAYER li1 ;
        RECT 110.040 136.490 110.470 138.070 ;
      LAYER li1 ;
        RECT 110.650 137.990 111.210 138.070 ;
        RECT 110.650 137.820 110.660 137.990 ;
        RECT 110.830 137.820 111.020 137.990 ;
        RECT 111.190 137.820 111.210 137.990 ;
        RECT 110.650 136.490 111.210 137.820 ;
        RECT 112.820 138.040 115.560 138.060 ;
        RECT 112.820 137.870 113.030 138.040 ;
        RECT 113.200 137.870 113.470 138.040 ;
        RECT 113.640 137.870 113.880 138.040 ;
        RECT 114.050 137.870 114.310 138.040 ;
        RECT 114.480 137.870 114.750 138.040 ;
        RECT 114.920 137.870 115.160 138.040 ;
        RECT 115.330 137.870 115.560 138.040 ;
        RECT 108.000 135.160 109.300 135.560 ;
        RECT 107.690 134.680 109.300 135.160 ;
      LAYER li1 ;
        RECT 110.040 134.810 110.290 136.490 ;
      LAYER li1 ;
        RECT 110.600 135.600 110.930 136.060 ;
      LAYER li1 ;
        RECT 111.390 135.780 111.720 137.570 ;
      LAYER li1 ;
        RECT 111.900 135.600 112.150 137.320 ;
        RECT 112.820 136.990 115.560 137.870 ;
        RECT 116.410 138.040 117.860 138.070 ;
        RECT 116.410 137.870 116.660 138.040 ;
        RECT 116.830 137.870 117.020 138.040 ;
        RECT 117.190 137.870 117.460 138.040 ;
        RECT 117.630 137.870 117.860 138.040 ;
        RECT 116.410 137.000 117.860 137.870 ;
        RECT 113.060 135.670 113.390 136.340 ;
        RECT 113.790 136.010 114.120 136.990 ;
        RECT 114.340 135.670 114.670 136.340 ;
        RECT 115.070 136.010 115.400 136.990 ;
        RECT 110.600 135.430 112.150 135.600 ;
        RECT 110.470 134.680 111.720 135.250 ;
        RECT 111.900 134.810 112.150 135.430 ;
        RECT 112.900 134.670 115.630 135.670 ;
        RECT 116.640 135.560 116.970 136.340 ;
        RECT 117.180 136.010 117.510 137.000 ;
      LAYER li1 ;
        RECT 118.200 136.490 118.630 138.070 ;
      LAYER li1 ;
        RECT 118.810 137.990 119.370 138.070 ;
        RECT 118.810 137.820 118.820 137.990 ;
        RECT 118.990 137.820 119.180 137.990 ;
        RECT 119.350 137.820 119.370 137.990 ;
        RECT 118.810 136.490 119.370 137.820 ;
        RECT 120.980 138.040 123.720 138.060 ;
        RECT 120.980 137.870 121.190 138.040 ;
        RECT 121.360 137.870 121.630 138.040 ;
        RECT 121.800 137.870 122.040 138.040 ;
        RECT 122.210 137.870 122.470 138.040 ;
        RECT 122.640 137.870 122.910 138.040 ;
        RECT 123.080 137.870 123.320 138.040 ;
        RECT 123.490 137.870 123.720 138.040 ;
        RECT 116.640 135.160 117.940 135.560 ;
        RECT 116.330 134.680 117.940 135.160 ;
      LAYER li1 ;
        RECT 118.200 134.810 118.450 136.490 ;
      LAYER li1 ;
        RECT 118.760 135.600 119.090 136.060 ;
      LAYER li1 ;
        RECT 119.550 135.780 119.880 137.570 ;
      LAYER li1 ;
        RECT 120.060 135.600 120.310 137.320 ;
        RECT 120.980 136.990 123.720 137.870 ;
        RECT 124.820 138.040 127.560 138.060 ;
        RECT 124.820 137.870 125.030 138.040 ;
        RECT 125.200 137.870 125.470 138.040 ;
        RECT 125.640 137.870 125.880 138.040 ;
        RECT 126.050 137.870 126.310 138.040 ;
        RECT 126.480 137.870 126.750 138.040 ;
        RECT 126.920 137.870 127.160 138.040 ;
        RECT 127.330 137.870 127.560 138.040 ;
        RECT 124.820 136.990 127.560 137.870 ;
        RECT 128.660 138.040 131.400 138.060 ;
        RECT 128.660 137.870 128.870 138.040 ;
        RECT 129.040 137.870 129.310 138.040 ;
        RECT 129.480 137.870 129.720 138.040 ;
        RECT 129.890 137.870 130.150 138.040 ;
        RECT 130.320 137.870 130.590 138.040 ;
        RECT 130.760 137.870 131.000 138.040 ;
        RECT 131.170 137.870 131.400 138.040 ;
        RECT 128.660 136.990 131.400 137.870 ;
        RECT 132.500 138.040 135.240 138.060 ;
        RECT 132.500 137.870 132.710 138.040 ;
        RECT 132.880 137.870 133.150 138.040 ;
        RECT 133.320 137.870 133.560 138.040 ;
        RECT 133.730 137.870 133.990 138.040 ;
        RECT 134.160 137.870 134.430 138.040 ;
        RECT 134.600 137.870 134.840 138.040 ;
        RECT 135.010 137.870 135.240 138.040 ;
        RECT 132.500 136.990 135.240 137.870 ;
        RECT 136.340 138.040 139.080 138.060 ;
        RECT 136.340 137.870 136.550 138.040 ;
        RECT 136.720 137.870 136.990 138.040 ;
        RECT 137.160 137.870 137.400 138.040 ;
        RECT 137.570 137.870 137.830 138.040 ;
        RECT 138.000 137.870 138.270 138.040 ;
        RECT 138.440 137.870 138.680 138.040 ;
        RECT 138.850 137.870 139.080 138.040 ;
        RECT 136.340 136.990 139.080 137.870 ;
        RECT 139.930 138.040 141.380 138.070 ;
        RECT 139.930 137.870 140.180 138.040 ;
        RECT 140.350 137.870 140.540 138.040 ;
        RECT 140.710 137.870 140.980 138.040 ;
        RECT 141.150 137.870 141.380 138.040 ;
        RECT 139.930 137.000 141.380 137.870 ;
        RECT 121.220 135.670 121.550 136.340 ;
        RECT 121.950 136.010 122.280 136.990 ;
        RECT 122.500 135.670 122.830 136.340 ;
        RECT 123.230 136.010 123.560 136.990 ;
        RECT 125.060 135.670 125.390 136.340 ;
        RECT 125.790 136.010 126.120 136.990 ;
        RECT 126.340 135.670 126.670 136.340 ;
        RECT 127.070 136.010 127.400 136.990 ;
        RECT 128.900 135.670 129.230 136.340 ;
        RECT 129.630 136.010 129.960 136.990 ;
        RECT 130.180 135.670 130.510 136.340 ;
        RECT 130.910 136.010 131.240 136.990 ;
        RECT 132.740 135.670 133.070 136.340 ;
        RECT 133.470 136.010 133.800 136.990 ;
        RECT 134.020 135.670 134.350 136.340 ;
        RECT 134.750 136.010 135.080 136.990 ;
        RECT 136.580 135.670 136.910 136.340 ;
        RECT 137.310 136.010 137.640 136.990 ;
        RECT 137.860 135.670 138.190 136.340 ;
        RECT 138.590 136.010 138.920 136.990 ;
        RECT 118.760 135.430 120.310 135.600 ;
        RECT 118.630 134.680 119.880 135.250 ;
        RECT 120.060 134.810 120.310 135.430 ;
        RECT 121.060 134.670 123.790 135.670 ;
        RECT 124.900 134.670 127.630 135.670 ;
        RECT 128.740 134.670 131.470 135.670 ;
        RECT 132.580 134.670 135.310 135.670 ;
        RECT 136.420 134.670 139.150 135.670 ;
        RECT 140.160 135.560 140.490 136.340 ;
        RECT 140.700 136.010 141.030 137.000 ;
        RECT 140.160 135.160 141.460 135.560 ;
        RECT 139.850 134.680 141.460 135.160 ;
        RECT 5.760 134.220 5.920 134.400 ;
        RECT 6.090 134.220 6.400 134.400 ;
        RECT 6.570 134.220 6.880 134.400 ;
        RECT 7.050 134.220 7.360 134.400 ;
        RECT 7.530 134.220 7.840 134.400 ;
        RECT 8.010 134.220 8.320 134.400 ;
        RECT 8.490 134.220 8.800 134.400 ;
        RECT 8.970 134.220 9.280 134.400 ;
        RECT 9.450 134.220 9.760 134.400 ;
        RECT 9.930 134.220 10.240 134.400 ;
        RECT 10.410 134.220 10.720 134.400 ;
        RECT 10.890 134.220 11.200 134.400 ;
        RECT 11.370 134.220 11.680 134.400 ;
        RECT 11.850 134.220 12.160 134.400 ;
        RECT 12.330 134.220 12.640 134.400 ;
        RECT 12.810 134.220 13.120 134.400 ;
        RECT 13.290 134.220 13.600 134.400 ;
        RECT 13.770 134.220 14.080 134.400 ;
        RECT 14.250 134.220 14.560 134.400 ;
        RECT 14.730 134.220 15.040 134.400 ;
        RECT 15.210 134.220 15.520 134.400 ;
        RECT 15.690 134.220 16.000 134.400 ;
        RECT 16.170 134.220 16.480 134.400 ;
        RECT 16.650 134.220 16.960 134.400 ;
        RECT 17.130 134.220 17.440 134.400 ;
        RECT 17.610 134.220 17.920 134.400 ;
        RECT 18.090 134.220 18.400 134.400 ;
        RECT 18.570 134.220 18.880 134.400 ;
        RECT 19.050 134.220 19.360 134.400 ;
        RECT 19.530 134.220 19.840 134.400 ;
        RECT 20.010 134.220 20.320 134.400 ;
        RECT 20.490 134.220 20.800 134.400 ;
        RECT 20.970 134.220 21.280 134.400 ;
        RECT 21.450 134.220 21.760 134.400 ;
        RECT 21.930 134.220 22.240 134.400 ;
        RECT 22.410 134.220 22.720 134.400 ;
        RECT 22.890 134.220 23.200 134.400 ;
        RECT 23.370 134.220 23.680 134.400 ;
        RECT 23.850 134.220 24.160 134.400 ;
        RECT 24.330 134.220 24.640 134.400 ;
        RECT 24.810 134.220 25.120 134.400 ;
        RECT 25.290 134.220 25.600 134.400 ;
        RECT 25.770 134.220 26.080 134.400 ;
        RECT 26.250 134.220 26.560 134.400 ;
        RECT 26.730 134.220 27.040 134.400 ;
        RECT 27.210 134.220 27.520 134.400 ;
        RECT 27.690 134.220 28.000 134.400 ;
        RECT 28.170 134.220 28.480 134.400 ;
        RECT 28.650 134.220 28.960 134.400 ;
        RECT 29.130 134.220 29.440 134.400 ;
        RECT 29.610 134.220 29.920 134.400 ;
        RECT 30.090 134.220 30.240 134.400 ;
        RECT 30.720 134.220 30.880 134.400 ;
        RECT 31.050 134.220 31.360 134.400 ;
        RECT 31.530 134.220 31.840 134.400 ;
        RECT 32.010 134.220 32.320 134.400 ;
        RECT 32.490 134.220 32.800 134.400 ;
        RECT 32.970 134.220 33.280 134.400 ;
        RECT 33.450 134.220 33.760 134.400 ;
        RECT 33.930 134.220 34.240 134.400 ;
        RECT 34.410 134.220 34.720 134.400 ;
        RECT 34.890 134.220 35.200 134.400 ;
        RECT 35.370 134.220 35.680 134.400 ;
        RECT 35.850 134.220 36.160 134.400 ;
        RECT 36.330 134.220 36.640 134.400 ;
        RECT 36.810 134.220 37.120 134.400 ;
        RECT 37.290 134.220 37.600 134.400 ;
        RECT 37.770 134.220 38.080 134.400 ;
        RECT 38.250 134.220 38.560 134.400 ;
        RECT 38.730 134.220 39.040 134.400 ;
        RECT 39.210 134.220 39.520 134.400 ;
        RECT 39.690 134.220 40.000 134.400 ;
        RECT 40.170 134.220 40.480 134.400 ;
        RECT 40.650 134.220 40.960 134.400 ;
        RECT 41.130 134.220 41.440 134.400 ;
        RECT 41.610 134.220 41.920 134.400 ;
        RECT 42.090 134.220 42.400 134.400 ;
        RECT 42.570 134.220 42.880 134.400 ;
        RECT 43.050 134.220 43.360 134.400 ;
        RECT 43.530 134.220 43.840 134.400 ;
        RECT 44.010 134.220 44.320 134.400 ;
        RECT 44.490 134.220 44.800 134.400 ;
        RECT 44.970 134.220 45.280 134.400 ;
        RECT 45.450 134.220 45.760 134.400 ;
        RECT 45.930 134.220 46.240 134.400 ;
        RECT 46.410 134.220 46.720 134.400 ;
        RECT 46.890 134.220 47.200 134.400 ;
        RECT 47.370 134.220 47.680 134.400 ;
        RECT 47.850 134.220 48.160 134.400 ;
        RECT 48.330 134.220 48.640 134.400 ;
        RECT 48.810 134.220 49.120 134.400 ;
        RECT 49.290 134.220 49.600 134.400 ;
        RECT 49.770 134.220 50.080 134.400 ;
        RECT 50.250 134.220 50.560 134.400 ;
        RECT 50.730 134.220 51.040 134.400 ;
        RECT 51.210 134.220 51.520 134.400 ;
        RECT 51.690 134.220 52.000 134.400 ;
        RECT 52.170 134.220 52.480 134.400 ;
        RECT 52.650 134.220 52.960 134.400 ;
        RECT 53.130 134.220 53.440 134.400 ;
        RECT 53.610 134.220 53.920 134.400 ;
        RECT 54.090 134.220 54.400 134.400 ;
        RECT 54.570 134.220 54.880 134.400 ;
        RECT 55.050 134.220 55.360 134.400 ;
        RECT 55.530 134.220 55.840 134.400 ;
        RECT 56.010 134.220 56.320 134.400 ;
        RECT 56.490 134.220 56.800 134.400 ;
        RECT 56.970 134.220 57.280 134.400 ;
        RECT 57.450 134.220 57.760 134.400 ;
        RECT 57.930 134.220 58.240 134.400 ;
        RECT 58.410 134.220 58.720 134.400 ;
        RECT 58.890 134.220 59.200 134.400 ;
        RECT 59.370 134.220 59.680 134.400 ;
        RECT 59.850 134.220 60.160 134.400 ;
        RECT 60.330 134.220 60.640 134.400 ;
        RECT 60.810 134.220 61.120 134.400 ;
        RECT 61.290 134.220 61.600 134.400 ;
        RECT 61.770 134.220 62.080 134.400 ;
        RECT 62.250 134.220 62.400 134.400 ;
        RECT 62.880 134.220 63.040 134.400 ;
        RECT 63.210 134.220 63.520 134.400 ;
        RECT 63.690 134.220 64.000 134.400 ;
        RECT 64.170 134.220 64.480 134.400 ;
        RECT 64.650 134.220 64.960 134.400 ;
        RECT 65.130 134.220 65.440 134.400 ;
        RECT 65.610 134.220 65.920 134.400 ;
        RECT 66.090 134.220 66.400 134.400 ;
        RECT 66.570 134.220 66.880 134.400 ;
        RECT 67.050 134.220 67.360 134.400 ;
        RECT 67.530 134.220 67.840 134.400 ;
        RECT 68.010 134.220 68.320 134.400 ;
        RECT 68.490 134.220 68.800 134.400 ;
        RECT 68.970 134.220 69.280 134.400 ;
        RECT 69.450 134.220 69.760 134.400 ;
        RECT 69.930 134.220 70.240 134.400 ;
        RECT 70.410 134.220 70.720 134.400 ;
        RECT 70.890 134.220 71.200 134.400 ;
        RECT 71.370 134.220 71.680 134.400 ;
        RECT 71.850 134.220 72.160 134.400 ;
        RECT 72.330 134.220 72.640 134.400 ;
        RECT 72.810 134.220 73.120 134.400 ;
        RECT 73.290 134.220 73.600 134.400 ;
        RECT 73.770 134.220 74.080 134.400 ;
        RECT 74.250 134.220 74.560 134.400 ;
        RECT 74.730 134.220 74.880 134.400 ;
        RECT 75.360 134.220 75.520 134.400 ;
        RECT 75.690 134.220 76.000 134.400 ;
        RECT 76.170 134.220 76.480 134.400 ;
        RECT 76.650 134.220 76.960 134.400 ;
        RECT 77.130 134.220 77.440 134.400 ;
        RECT 77.610 134.220 77.920 134.400 ;
        RECT 78.090 134.220 78.400 134.400 ;
        RECT 78.570 134.220 78.880 134.400 ;
        RECT 79.050 134.220 79.360 134.400 ;
        RECT 79.530 134.220 79.840 134.400 ;
        RECT 80.010 134.220 80.320 134.400 ;
        RECT 80.490 134.220 80.800 134.400 ;
        RECT 80.970 134.220 81.280 134.400 ;
        RECT 81.450 134.220 81.760 134.400 ;
        RECT 81.930 134.220 82.240 134.400 ;
        RECT 82.410 134.220 82.720 134.400 ;
        RECT 82.890 134.220 83.200 134.400 ;
        RECT 83.370 134.220 83.680 134.400 ;
        RECT 83.850 134.220 84.160 134.400 ;
        RECT 84.330 134.220 84.640 134.400 ;
        RECT 84.810 134.220 85.120 134.400 ;
        RECT 85.290 134.220 85.600 134.400 ;
        RECT 85.770 134.220 86.080 134.400 ;
        RECT 86.250 134.220 86.560 134.400 ;
        RECT 86.730 134.220 87.040 134.400 ;
        RECT 87.210 134.220 87.520 134.400 ;
        RECT 87.690 134.220 88.000 134.400 ;
        RECT 88.170 134.220 88.480 134.400 ;
        RECT 88.650 134.220 88.960 134.400 ;
        RECT 89.130 134.220 89.440 134.400 ;
        RECT 89.610 134.220 89.920 134.400 ;
        RECT 90.090 134.220 90.400 134.400 ;
        RECT 90.570 134.220 90.880 134.400 ;
        RECT 91.050 134.220 91.360 134.400 ;
        RECT 91.530 134.220 91.840 134.400 ;
        RECT 92.010 134.220 92.320 134.400 ;
        RECT 92.490 134.220 92.800 134.400 ;
        RECT 92.970 134.220 93.280 134.400 ;
        RECT 93.450 134.220 93.760 134.400 ;
        RECT 93.930 134.220 94.240 134.400 ;
        RECT 94.410 134.220 94.720 134.400 ;
        RECT 94.890 134.220 95.200 134.400 ;
        RECT 95.370 134.220 95.680 134.400 ;
        RECT 95.850 134.220 96.160 134.400 ;
        RECT 96.330 134.220 96.640 134.400 ;
        RECT 96.810 134.220 97.120 134.400 ;
        RECT 97.290 134.220 97.600 134.400 ;
        RECT 97.770 134.220 97.920 134.400 ;
        RECT 98.400 134.220 98.560 134.400 ;
        RECT 98.730 134.220 99.040 134.400 ;
        RECT 99.210 134.220 99.520 134.400 ;
        RECT 99.690 134.220 100.000 134.400 ;
        RECT 100.170 134.220 100.480 134.400 ;
        RECT 100.650 134.220 100.960 134.400 ;
        RECT 101.130 134.220 101.440 134.400 ;
        RECT 101.610 134.220 101.920 134.400 ;
        RECT 102.090 134.220 102.400 134.400 ;
        RECT 102.570 134.220 102.880 134.400 ;
        RECT 103.050 134.220 103.360 134.400 ;
        RECT 103.530 134.220 103.840 134.400 ;
        RECT 104.010 134.220 104.320 134.400 ;
        RECT 104.490 134.220 104.800 134.400 ;
        RECT 104.970 134.220 105.280 134.400 ;
        RECT 105.450 134.220 105.760 134.400 ;
        RECT 105.930 134.220 106.240 134.400 ;
        RECT 106.410 134.220 106.720 134.400 ;
        RECT 106.890 134.220 107.200 134.400 ;
        RECT 107.370 134.220 107.680 134.400 ;
        RECT 107.850 134.220 108.160 134.400 ;
        RECT 108.330 134.220 108.640 134.400 ;
        RECT 108.810 134.220 109.120 134.400 ;
        RECT 109.290 134.220 109.440 134.400 ;
        RECT 109.920 134.220 110.080 134.400 ;
        RECT 110.250 134.220 110.560 134.400 ;
        RECT 110.730 134.220 111.040 134.400 ;
        RECT 111.210 134.220 111.520 134.400 ;
        RECT 111.690 134.220 112.000 134.400 ;
        RECT 112.170 134.220 112.480 134.400 ;
        RECT 112.650 134.220 112.960 134.400 ;
        RECT 113.130 134.220 113.440 134.400 ;
        RECT 113.610 134.220 113.920 134.400 ;
        RECT 114.090 134.220 114.400 134.400 ;
        RECT 114.570 134.220 114.880 134.400 ;
        RECT 115.050 134.220 115.360 134.400 ;
        RECT 115.530 134.220 115.840 134.400 ;
        RECT 116.010 134.220 116.320 134.400 ;
        RECT 116.490 134.220 116.800 134.400 ;
        RECT 116.970 134.220 117.280 134.400 ;
        RECT 117.450 134.220 117.760 134.400 ;
        RECT 117.930 134.220 118.240 134.400 ;
        RECT 118.410 134.220 118.720 134.400 ;
        RECT 118.890 134.220 119.200 134.400 ;
        RECT 119.370 134.220 119.680 134.400 ;
        RECT 119.850 134.220 120.160 134.400 ;
        RECT 120.330 134.220 120.640 134.400 ;
        RECT 120.810 134.220 121.120 134.400 ;
        RECT 121.290 134.220 121.600 134.400 ;
        RECT 121.770 134.220 122.080 134.400 ;
        RECT 122.250 134.220 122.560 134.400 ;
        RECT 122.730 134.220 123.040 134.400 ;
        RECT 123.210 134.220 123.520 134.400 ;
        RECT 123.690 134.220 124.000 134.400 ;
        RECT 124.170 134.220 124.480 134.400 ;
        RECT 124.650 134.220 124.960 134.400 ;
        RECT 125.130 134.220 125.440 134.400 ;
        RECT 125.610 134.220 125.920 134.400 ;
        RECT 126.090 134.220 126.400 134.400 ;
        RECT 126.570 134.220 126.880 134.400 ;
        RECT 127.050 134.220 127.360 134.400 ;
        RECT 127.530 134.220 127.840 134.400 ;
        RECT 128.010 134.220 128.320 134.400 ;
        RECT 128.490 134.220 128.800 134.400 ;
        RECT 128.970 134.220 129.280 134.400 ;
        RECT 129.450 134.220 129.760 134.400 ;
        RECT 129.930 134.220 130.240 134.400 ;
        RECT 130.410 134.220 130.720 134.400 ;
        RECT 130.890 134.220 131.200 134.400 ;
        RECT 131.370 134.220 131.680 134.400 ;
        RECT 131.850 134.220 132.160 134.400 ;
        RECT 132.330 134.220 132.640 134.400 ;
        RECT 132.810 134.220 133.120 134.400 ;
        RECT 133.290 134.220 133.600 134.400 ;
        RECT 133.770 134.220 134.080 134.400 ;
        RECT 134.250 134.220 134.560 134.400 ;
        RECT 134.730 134.220 135.040 134.400 ;
        RECT 135.210 134.220 135.520 134.400 ;
        RECT 135.690 134.220 136.000 134.400 ;
        RECT 136.170 134.220 136.480 134.400 ;
        RECT 136.650 134.220 136.960 134.400 ;
        RECT 137.130 134.220 137.440 134.400 ;
        RECT 137.610 134.220 137.920 134.400 ;
        RECT 138.090 134.220 138.400 134.400 ;
        RECT 138.570 134.220 138.880 134.400 ;
        RECT 139.050 134.220 139.360 134.400 ;
        RECT 139.530 134.220 139.840 134.400 ;
        RECT 140.010 134.220 140.320 134.400 ;
        RECT 140.490 134.220 140.800 134.400 ;
        RECT 140.970 134.220 141.280 134.400 ;
        RECT 141.450 134.220 141.600 134.400 ;
        RECT 6.340 133.920 9.070 133.950 ;
        RECT 6.340 133.750 6.510 133.920 ;
        RECT 6.680 133.750 6.950 133.920 ;
        RECT 7.120 133.750 7.360 133.920 ;
        RECT 7.530 133.750 7.790 133.920 ;
        RECT 7.960 133.750 8.230 133.920 ;
        RECT 8.400 133.750 8.640 133.920 ;
        RECT 8.810 133.750 9.070 133.920 ;
        RECT 12.100 133.910 12.750 134.020 ;
        RECT 6.340 132.950 9.070 133.750 ;
      LAYER li1 ;
        RECT 10.850 133.240 11.430 133.880 ;
      LAYER li1 ;
        RECT 12.100 133.740 12.160 133.910 ;
        RECT 12.330 133.740 12.520 133.910 ;
        RECT 12.690 133.740 12.750 133.910 ;
        RECT 12.100 133.680 12.750 133.740 ;
        RECT 12.340 133.240 12.750 133.680 ;
        RECT 13.540 133.920 16.270 133.950 ;
        RECT 13.540 133.750 13.710 133.920 ;
        RECT 13.880 133.750 14.150 133.920 ;
        RECT 14.320 133.750 14.560 133.920 ;
        RECT 14.730 133.750 14.990 133.920 ;
        RECT 15.160 133.750 15.430 133.920 ;
        RECT 15.600 133.750 15.840 133.920 ;
        RECT 16.010 133.750 16.270 133.920 ;
        RECT 6.500 132.280 6.830 132.950 ;
        RECT 7.230 131.630 7.560 132.610 ;
        RECT 7.780 132.280 8.110 132.950 ;
        RECT 8.510 131.630 8.840 132.610 ;
      LAYER li1 ;
        RECT 11.180 132.370 11.430 133.240 ;
      LAYER li1 ;
        RECT 13.540 132.950 16.270 133.750 ;
        RECT 17.380 133.920 20.110 133.950 ;
        RECT 17.380 133.750 17.550 133.920 ;
        RECT 17.720 133.750 17.990 133.920 ;
        RECT 18.160 133.750 18.400 133.920 ;
        RECT 18.570 133.750 18.830 133.920 ;
        RECT 19.000 133.750 19.270 133.920 ;
        RECT 19.440 133.750 19.680 133.920 ;
        RECT 19.850 133.750 20.110 133.920 ;
        RECT 17.380 132.950 20.110 133.750 ;
        RECT 21.220 133.920 23.950 133.950 ;
        RECT 21.220 133.750 21.390 133.920 ;
        RECT 21.560 133.750 21.830 133.920 ;
        RECT 22.000 133.750 22.240 133.920 ;
        RECT 22.410 133.750 22.670 133.920 ;
        RECT 22.840 133.750 23.110 133.920 ;
        RECT 23.280 133.750 23.520 133.920 ;
        RECT 23.690 133.750 23.950 133.920 ;
        RECT 21.220 132.950 23.950 133.750 ;
        RECT 25.060 133.920 27.790 133.950 ;
        RECT 25.060 133.750 25.230 133.920 ;
        RECT 25.400 133.750 25.670 133.920 ;
        RECT 25.840 133.750 26.080 133.920 ;
        RECT 26.250 133.750 26.510 133.920 ;
        RECT 26.680 133.750 26.950 133.920 ;
        RECT 27.120 133.750 27.360 133.920 ;
        RECT 27.530 133.750 27.790 133.920 ;
        RECT 25.060 132.950 27.790 133.750 ;
        RECT 28.490 133.910 30.100 133.940 ;
        RECT 28.490 133.740 28.540 133.910 ;
        RECT 28.710 133.740 28.980 133.910 ;
        RECT 29.150 133.740 29.420 133.910 ;
        RECT 29.590 133.740 29.830 133.910 ;
        RECT 30.000 133.740 30.100 133.910 ;
        RECT 28.490 133.460 30.100 133.740 ;
        RECT 28.800 133.060 30.100 133.460 ;
        RECT 31.840 133.870 33.650 134.040 ;
      LAYER li1 ;
        RECT 11.180 132.120 11.890 132.370 ;
      LAYER li1 ;
        RECT 13.700 132.280 14.030 132.950 ;
        RECT 6.260 130.750 9.000 131.630 ;
        RECT 6.260 130.580 6.470 130.750 ;
        RECT 6.640 130.580 6.910 130.750 ;
        RECT 7.080 130.580 7.320 130.750 ;
        RECT 7.490 130.580 7.750 130.750 ;
        RECT 7.920 130.580 8.190 130.750 ;
        RECT 8.360 130.580 8.600 130.750 ;
        RECT 8.770 130.580 9.000 130.750 ;
        RECT 6.260 130.560 9.000 130.580 ;
        RECT 10.780 130.860 11.180 131.130 ;
        RECT 10.780 130.800 11.430 130.860 ;
        RECT 10.780 130.630 10.840 130.800 ;
        RECT 11.010 130.630 11.200 130.800 ;
        RECT 11.370 130.630 11.430 130.800 ;
      LAYER li1 ;
        RECT 11.640 130.780 11.890 132.120 ;
      LAYER li1 ;
        RECT 14.430 131.630 14.760 132.610 ;
        RECT 14.980 132.280 15.310 132.950 ;
        RECT 15.710 131.630 16.040 132.610 ;
        RECT 17.540 132.280 17.870 132.950 ;
        RECT 18.270 131.630 18.600 132.610 ;
        RECT 18.820 132.280 19.150 132.950 ;
        RECT 19.550 131.630 19.880 132.610 ;
        RECT 21.380 132.280 21.710 132.950 ;
        RECT 22.110 131.630 22.440 132.610 ;
        RECT 22.660 132.280 22.990 132.950 ;
        RECT 23.390 131.630 23.720 132.610 ;
        RECT 25.220 132.280 25.550 132.950 ;
        RECT 25.950 131.630 26.280 132.610 ;
        RECT 26.500 132.280 26.830 132.950 ;
        RECT 27.230 131.630 27.560 132.610 ;
        RECT 28.800 132.280 29.130 133.060 ;
        RECT 31.840 132.950 32.170 133.870 ;
      LAYER li1 ;
        RECT 32.420 133.470 32.950 133.690 ;
        RECT 32.420 133.300 32.960 133.470 ;
        RECT 32.420 132.950 32.950 133.300 ;
      LAYER li1 ;
        RECT 10.780 130.520 11.430 130.630 ;
        RECT 13.460 130.750 16.200 131.630 ;
        RECT 13.460 130.580 13.670 130.750 ;
        RECT 13.840 130.580 14.110 130.750 ;
        RECT 14.280 130.580 14.520 130.750 ;
        RECT 14.690 130.580 14.950 130.750 ;
        RECT 15.120 130.580 15.390 130.750 ;
        RECT 15.560 130.580 15.800 130.750 ;
        RECT 15.970 130.580 16.200 130.750 ;
        RECT 13.460 130.560 16.200 130.580 ;
        RECT 17.300 130.750 20.040 131.630 ;
        RECT 17.300 130.580 17.510 130.750 ;
        RECT 17.680 130.580 17.950 130.750 ;
        RECT 18.120 130.580 18.360 130.750 ;
        RECT 18.530 130.580 18.790 130.750 ;
        RECT 18.960 130.580 19.230 130.750 ;
        RECT 19.400 130.580 19.640 130.750 ;
        RECT 19.810 130.580 20.040 130.750 ;
        RECT 17.300 130.560 20.040 130.580 ;
        RECT 21.140 130.750 23.880 131.630 ;
        RECT 21.140 130.580 21.350 130.750 ;
        RECT 21.520 130.580 21.790 130.750 ;
        RECT 21.960 130.580 22.200 130.750 ;
        RECT 22.370 130.580 22.630 130.750 ;
        RECT 22.800 130.580 23.070 130.750 ;
        RECT 23.240 130.580 23.480 130.750 ;
        RECT 23.650 130.580 23.880 130.750 ;
        RECT 21.140 130.560 23.880 130.580 ;
        RECT 24.980 130.750 27.720 131.630 ;
        RECT 29.340 131.620 29.670 132.610 ;
      LAYER li1 ;
        RECT 31.810 132.440 32.230 132.770 ;
        RECT 32.420 132.380 32.590 132.950 ;
      LAYER li1 ;
        RECT 33.480 132.850 33.650 133.870 ;
        RECT 33.830 133.910 34.930 133.940 ;
        RECT 33.830 133.740 33.880 133.910 ;
        RECT 34.050 133.740 34.240 133.910 ;
        RECT 34.410 133.740 34.600 133.910 ;
        RECT 34.770 133.740 34.930 133.910 ;
        RECT 36.100 133.920 38.830 133.950 ;
        RECT 33.830 133.030 34.930 133.740 ;
        RECT 35.100 132.850 35.350 133.780 ;
        RECT 36.100 133.750 36.270 133.920 ;
        RECT 36.440 133.750 36.710 133.920 ;
        RECT 36.880 133.750 37.120 133.920 ;
        RECT 37.290 133.750 37.550 133.920 ;
        RECT 37.720 133.750 37.990 133.920 ;
        RECT 38.160 133.750 38.400 133.920 ;
        RECT 38.570 133.750 38.830 133.920 ;
        RECT 36.100 132.950 38.830 133.750 ;
        RECT 39.940 133.920 42.670 133.950 ;
        RECT 39.940 133.750 40.110 133.920 ;
        RECT 40.280 133.750 40.550 133.920 ;
        RECT 40.720 133.750 40.960 133.920 ;
        RECT 41.130 133.750 41.390 133.920 ;
        RECT 41.560 133.750 41.830 133.920 ;
        RECT 42.000 133.750 42.240 133.920 ;
        RECT 42.410 133.750 42.670 133.920 ;
        RECT 39.940 132.950 42.670 133.750 ;
        RECT 43.780 133.920 46.510 133.950 ;
        RECT 43.780 133.750 43.950 133.920 ;
        RECT 44.120 133.750 44.390 133.920 ;
        RECT 44.560 133.750 44.800 133.920 ;
        RECT 44.970 133.750 45.230 133.920 ;
        RECT 45.400 133.750 45.670 133.920 ;
        RECT 45.840 133.750 46.080 133.920 ;
        RECT 46.250 133.750 46.510 133.920 ;
        RECT 43.780 132.950 46.510 133.750 ;
        RECT 47.620 133.920 50.350 133.950 ;
        RECT 47.620 133.750 47.790 133.920 ;
        RECT 47.960 133.750 48.230 133.920 ;
        RECT 48.400 133.750 48.640 133.920 ;
        RECT 48.810 133.750 49.070 133.920 ;
        RECT 49.240 133.750 49.510 133.920 ;
        RECT 49.680 133.750 49.920 133.920 ;
        RECT 50.090 133.750 50.350 133.920 ;
        RECT 47.620 132.950 50.350 133.750 ;
        RECT 51.460 133.920 54.190 133.950 ;
        RECT 51.460 133.750 51.630 133.920 ;
        RECT 51.800 133.750 52.070 133.920 ;
        RECT 52.240 133.750 52.480 133.920 ;
        RECT 52.650 133.750 52.910 133.920 ;
        RECT 53.080 133.750 53.350 133.920 ;
        RECT 53.520 133.750 53.760 133.920 ;
        RECT 53.930 133.750 54.190 133.920 ;
        RECT 51.460 132.950 54.190 133.750 ;
        RECT 55.300 133.920 58.030 133.950 ;
        RECT 55.300 133.750 55.470 133.920 ;
        RECT 55.640 133.750 55.910 133.920 ;
        RECT 56.080 133.750 56.320 133.920 ;
        RECT 56.490 133.750 56.750 133.920 ;
        RECT 56.920 133.750 57.190 133.920 ;
        RECT 57.360 133.750 57.600 133.920 ;
        RECT 57.770 133.750 58.030 133.920 ;
        RECT 55.300 132.950 58.030 133.750 ;
        RECT 59.140 133.920 61.870 133.950 ;
        RECT 59.140 133.750 59.310 133.920 ;
        RECT 59.480 133.750 59.750 133.920 ;
        RECT 59.920 133.750 60.160 133.920 ;
        RECT 60.330 133.750 60.590 133.920 ;
        RECT 60.760 133.750 61.030 133.920 ;
        RECT 61.200 133.750 61.440 133.920 ;
        RECT 61.610 133.750 61.870 133.920 ;
        RECT 59.140 132.950 61.870 133.750 ;
        RECT 62.980 133.920 65.710 133.950 ;
        RECT 62.980 133.750 63.150 133.920 ;
        RECT 63.320 133.750 63.590 133.920 ;
        RECT 63.760 133.750 64.000 133.920 ;
        RECT 64.170 133.750 64.430 133.920 ;
        RECT 64.600 133.750 64.870 133.920 ;
        RECT 65.040 133.750 65.280 133.920 ;
        RECT 65.450 133.750 65.710 133.920 ;
        RECT 62.980 132.950 65.710 133.750 ;
        RECT 66.820 133.920 69.550 133.950 ;
        RECT 66.820 133.750 66.990 133.920 ;
        RECT 67.160 133.750 67.430 133.920 ;
        RECT 67.600 133.750 67.840 133.920 ;
        RECT 68.010 133.750 68.270 133.920 ;
        RECT 68.440 133.750 68.710 133.920 ;
        RECT 68.880 133.750 69.120 133.920 ;
        RECT 69.290 133.750 69.550 133.920 ;
        RECT 66.820 132.950 69.550 133.750 ;
        RECT 70.250 133.910 71.860 133.940 ;
        RECT 70.250 133.740 70.300 133.910 ;
        RECT 70.470 133.740 70.740 133.910 ;
        RECT 70.910 133.740 71.180 133.910 ;
        RECT 71.350 133.740 71.590 133.910 ;
        RECT 71.760 133.740 71.860 133.910 ;
        RECT 75.080 133.910 76.070 133.940 ;
        RECT 70.250 133.460 71.860 133.740 ;
        RECT 70.560 133.060 71.860 133.460 ;
        RECT 73.570 133.480 73.820 133.810 ;
        RECT 75.080 133.740 75.130 133.910 ;
        RECT 75.300 133.740 75.490 133.910 ;
        RECT 75.660 133.740 75.850 133.910 ;
        RECT 76.020 133.740 76.070 133.910 ;
        RECT 76.970 133.910 78.580 133.940 ;
        RECT 73.570 133.310 74.330 133.480 ;
      LAYER li1 ;
        RECT 32.770 132.560 33.280 132.770 ;
      LAYER li1 ;
        RECT 33.480 132.680 35.350 132.850 ;
      LAYER li1 ;
        RECT 32.420 132.210 33.480 132.380 ;
        RECT 33.210 132.130 33.480 132.210 ;
        RECT 33.930 132.190 34.440 132.500 ;
        RECT 34.690 132.190 35.400 132.500 ;
      LAYER li1 ;
        RECT 36.260 132.280 36.590 132.950 ;
        RECT 24.980 130.580 25.190 130.750 ;
        RECT 25.360 130.580 25.630 130.750 ;
        RECT 25.800 130.580 26.040 130.750 ;
        RECT 26.210 130.580 26.470 130.750 ;
        RECT 26.640 130.580 26.910 130.750 ;
        RECT 27.080 130.580 27.320 130.750 ;
        RECT 27.490 130.580 27.720 130.750 ;
        RECT 24.980 130.560 27.720 130.580 ;
        RECT 28.570 130.750 30.020 131.620 ;
        RECT 28.570 130.580 28.820 130.750 ;
        RECT 28.990 130.580 29.180 130.750 ;
        RECT 29.350 130.580 29.620 130.750 ;
        RECT 29.790 130.580 30.020 130.750 ;
        RECT 28.570 130.550 30.020 130.580 ;
        RECT 31.770 130.800 33.030 132.030 ;
      LAYER li1 ;
        RECT 33.210 131.050 33.730 132.130 ;
      LAYER li1 ;
        RECT 31.770 130.630 31.780 130.800 ;
        RECT 31.950 130.630 32.140 130.800 ;
        RECT 32.310 130.630 32.500 130.800 ;
        RECT 32.670 130.630 32.860 130.800 ;
        RECT 31.770 130.550 33.030 130.630 ;
      LAYER li1 ;
        RECT 33.560 130.550 33.730 131.050 ;
      LAYER li1 ;
        RECT 33.990 130.800 35.300 132.010 ;
        RECT 36.990 131.630 37.320 132.610 ;
        RECT 37.540 132.280 37.870 132.950 ;
        RECT 38.270 131.630 38.600 132.610 ;
        RECT 40.100 132.280 40.430 132.950 ;
        RECT 40.830 131.630 41.160 132.610 ;
        RECT 41.380 132.280 41.710 132.950 ;
        RECT 42.110 131.630 42.440 132.610 ;
        RECT 43.940 132.280 44.270 132.950 ;
        RECT 44.670 131.630 45.000 132.610 ;
        RECT 45.220 132.280 45.550 132.950 ;
        RECT 45.950 131.630 46.280 132.610 ;
        RECT 47.780 132.280 48.110 132.950 ;
        RECT 48.510 131.630 48.840 132.610 ;
        RECT 49.060 132.280 49.390 132.950 ;
        RECT 49.790 131.630 50.120 132.610 ;
        RECT 51.620 132.280 51.950 132.950 ;
        RECT 52.350 131.630 52.680 132.610 ;
        RECT 52.900 132.280 53.230 132.950 ;
        RECT 53.630 131.630 53.960 132.610 ;
        RECT 55.460 132.280 55.790 132.950 ;
        RECT 56.190 131.630 56.520 132.610 ;
        RECT 56.740 132.280 57.070 132.950 ;
        RECT 57.470 131.630 57.800 132.610 ;
        RECT 59.300 132.280 59.630 132.950 ;
        RECT 60.030 131.630 60.360 132.610 ;
        RECT 60.580 132.280 60.910 132.950 ;
        RECT 61.310 131.630 61.640 132.610 ;
        RECT 63.140 132.280 63.470 132.950 ;
        RECT 63.870 131.630 64.200 132.610 ;
        RECT 64.420 132.280 64.750 132.950 ;
        RECT 65.150 131.630 65.480 132.610 ;
        RECT 66.980 132.280 67.310 132.950 ;
        RECT 67.710 131.630 68.040 132.610 ;
        RECT 68.260 132.280 68.590 132.950 ;
        RECT 68.990 131.630 69.320 132.610 ;
        RECT 70.560 132.280 70.890 133.060 ;
        RECT 33.990 130.630 34.020 130.800 ;
        RECT 34.190 130.630 34.380 130.800 ;
        RECT 34.550 130.630 34.740 130.800 ;
        RECT 34.910 130.630 35.100 130.800 ;
        RECT 35.270 130.630 35.300 130.800 ;
        RECT 33.990 130.550 35.300 130.630 ;
        RECT 36.020 130.750 38.760 131.630 ;
        RECT 36.020 130.580 36.230 130.750 ;
        RECT 36.400 130.580 36.670 130.750 ;
        RECT 36.840 130.580 37.080 130.750 ;
        RECT 37.250 130.580 37.510 130.750 ;
        RECT 37.680 130.580 37.950 130.750 ;
        RECT 38.120 130.580 38.360 130.750 ;
        RECT 38.530 130.580 38.760 130.750 ;
        RECT 36.020 130.560 38.760 130.580 ;
        RECT 39.860 130.750 42.600 131.630 ;
        RECT 39.860 130.580 40.070 130.750 ;
        RECT 40.240 130.580 40.510 130.750 ;
        RECT 40.680 130.580 40.920 130.750 ;
        RECT 41.090 130.580 41.350 130.750 ;
        RECT 41.520 130.580 41.790 130.750 ;
        RECT 41.960 130.580 42.200 130.750 ;
        RECT 42.370 130.580 42.600 130.750 ;
        RECT 39.860 130.560 42.600 130.580 ;
        RECT 43.700 130.750 46.440 131.630 ;
        RECT 43.700 130.580 43.910 130.750 ;
        RECT 44.080 130.580 44.350 130.750 ;
        RECT 44.520 130.580 44.760 130.750 ;
        RECT 44.930 130.580 45.190 130.750 ;
        RECT 45.360 130.580 45.630 130.750 ;
        RECT 45.800 130.580 46.040 130.750 ;
        RECT 46.210 130.580 46.440 130.750 ;
        RECT 43.700 130.560 46.440 130.580 ;
        RECT 47.540 130.750 50.280 131.630 ;
        RECT 47.540 130.580 47.750 130.750 ;
        RECT 47.920 130.580 48.190 130.750 ;
        RECT 48.360 130.580 48.600 130.750 ;
        RECT 48.770 130.580 49.030 130.750 ;
        RECT 49.200 130.580 49.470 130.750 ;
        RECT 49.640 130.580 49.880 130.750 ;
        RECT 50.050 130.580 50.280 130.750 ;
        RECT 47.540 130.560 50.280 130.580 ;
        RECT 51.380 130.750 54.120 131.630 ;
        RECT 51.380 130.580 51.590 130.750 ;
        RECT 51.760 130.580 52.030 130.750 ;
        RECT 52.200 130.580 52.440 130.750 ;
        RECT 52.610 130.580 52.870 130.750 ;
        RECT 53.040 130.580 53.310 130.750 ;
        RECT 53.480 130.580 53.720 130.750 ;
        RECT 53.890 130.580 54.120 130.750 ;
        RECT 51.380 130.560 54.120 130.580 ;
        RECT 55.220 130.750 57.960 131.630 ;
        RECT 55.220 130.580 55.430 130.750 ;
        RECT 55.600 130.580 55.870 130.750 ;
        RECT 56.040 130.580 56.280 130.750 ;
        RECT 56.450 130.580 56.710 130.750 ;
        RECT 56.880 130.580 57.150 130.750 ;
        RECT 57.320 130.580 57.560 130.750 ;
        RECT 57.730 130.580 57.960 130.750 ;
        RECT 55.220 130.560 57.960 130.580 ;
        RECT 59.060 130.750 61.800 131.630 ;
        RECT 59.060 130.580 59.270 130.750 ;
        RECT 59.440 130.580 59.710 130.750 ;
        RECT 59.880 130.580 60.120 130.750 ;
        RECT 60.290 130.580 60.550 130.750 ;
        RECT 60.720 130.580 60.990 130.750 ;
        RECT 61.160 130.580 61.400 130.750 ;
        RECT 61.570 130.580 61.800 130.750 ;
        RECT 59.060 130.560 61.800 130.580 ;
        RECT 62.900 130.750 65.640 131.630 ;
        RECT 62.900 130.580 63.110 130.750 ;
        RECT 63.280 130.580 63.550 130.750 ;
        RECT 63.720 130.580 63.960 130.750 ;
        RECT 64.130 130.580 64.390 130.750 ;
        RECT 64.560 130.580 64.830 130.750 ;
        RECT 65.000 130.580 65.240 130.750 ;
        RECT 65.410 130.580 65.640 130.750 ;
        RECT 62.900 130.560 65.640 130.580 ;
        RECT 66.740 130.750 69.480 131.630 ;
        RECT 71.100 131.620 71.430 132.610 ;
        RECT 74.160 132.400 74.330 133.310 ;
      LAYER li1 ;
        RECT 74.510 132.580 74.900 133.500 ;
      LAYER li1 ;
        RECT 75.080 132.980 76.070 133.740 ;
        RECT 75.890 132.400 76.220 132.580 ;
        RECT 74.160 132.230 76.220 132.400 ;
        RECT 66.740 130.580 66.950 130.750 ;
        RECT 67.120 130.580 67.390 130.750 ;
        RECT 67.560 130.580 67.800 130.750 ;
        RECT 67.970 130.580 68.230 130.750 ;
        RECT 68.400 130.580 68.670 130.750 ;
        RECT 68.840 130.580 69.080 130.750 ;
        RECT 69.250 130.580 69.480 130.750 ;
        RECT 66.740 130.560 69.480 130.580 ;
        RECT 70.330 130.750 71.780 131.620 ;
        RECT 70.330 130.580 70.580 130.750 ;
        RECT 70.750 130.580 70.940 130.750 ;
        RECT 71.110 130.580 71.380 130.750 ;
        RECT 71.550 130.580 71.780 130.750 ;
        RECT 73.530 130.800 74.460 132.050 ;
        RECT 74.640 131.630 74.810 132.230 ;
        RECT 74.990 130.800 76.240 132.050 ;
        RECT 73.530 130.630 73.550 130.800 ;
        RECT 73.720 130.630 73.910 130.800 ;
        RECT 74.080 130.630 74.270 130.800 ;
        RECT 74.440 130.630 74.460 130.800 ;
        RECT 75.160 130.630 75.350 130.800 ;
        RECT 75.520 130.630 75.710 130.800 ;
        RECT 75.880 130.630 76.070 130.800 ;
        RECT 73.530 130.600 74.460 130.630 ;
        RECT 70.330 130.550 71.780 130.580 ;
        RECT 74.990 130.550 76.240 130.630 ;
      LAYER li1 ;
        RECT 76.420 130.550 76.700 133.810 ;
      LAYER li1 ;
        RECT 76.970 133.740 77.020 133.910 ;
        RECT 77.190 133.740 77.460 133.910 ;
        RECT 77.630 133.740 77.900 133.910 ;
        RECT 78.070 133.740 78.310 133.910 ;
        RECT 78.480 133.740 78.580 133.910 ;
        RECT 76.970 133.460 78.580 133.740 ;
        RECT 77.280 133.060 78.580 133.460 ;
        RECT 78.810 133.910 79.400 133.940 ;
        RECT 78.810 133.740 78.840 133.910 ;
        RECT 79.010 133.740 79.200 133.910 ;
        RECT 79.370 133.740 79.400 133.910 ;
        RECT 80.080 133.910 81.030 133.940 ;
        RECT 77.280 132.280 77.610 133.060 ;
        RECT 78.810 132.980 79.400 133.740 ;
      LAYER li1 ;
        RECT 79.650 132.880 79.900 133.810 ;
      LAYER li1 ;
        RECT 80.080 133.740 80.110 133.910 ;
        RECT 80.280 133.740 80.470 133.910 ;
        RECT 80.640 133.740 80.830 133.910 ;
        RECT 81.000 133.740 81.030 133.910 ;
        RECT 82.250 133.910 83.860 133.940 ;
        RECT 85.520 133.910 86.410 133.940 ;
        RECT 80.080 133.060 81.030 133.740 ;
      LAYER li1 ;
        RECT 81.210 132.880 81.480 133.810 ;
      LAYER li1 ;
        RECT 82.250 133.740 82.300 133.910 ;
        RECT 82.470 133.740 82.740 133.910 ;
        RECT 82.910 133.740 83.180 133.910 ;
        RECT 83.350 133.740 83.590 133.910 ;
        RECT 83.760 133.740 83.860 133.910 ;
        RECT 82.250 133.460 83.860 133.740 ;
        RECT 77.820 131.620 78.150 132.610 ;
      LAYER li1 ;
        RECT 78.850 132.190 79.150 132.780 ;
        RECT 79.650 132.710 81.480 132.880 ;
        RECT 79.330 132.190 80.520 132.530 ;
      LAYER li1 ;
        RECT 77.050 130.750 78.500 131.620 ;
        RECT 77.050 130.580 77.300 130.750 ;
        RECT 77.470 130.580 77.660 130.750 ;
        RECT 77.830 130.580 78.100 130.750 ;
        RECT 78.270 130.580 78.500 130.750 ;
        RECT 77.050 130.550 78.500 130.580 ;
        RECT 78.810 130.800 80.480 132.010 ;
      LAYER li1 ;
        RECT 80.700 131.050 81.030 132.530 ;
      LAYER li1 ;
        RECT 78.810 130.630 78.840 130.800 ;
        RECT 79.010 130.630 79.200 130.800 ;
        RECT 79.370 130.630 79.560 130.800 ;
        RECT 79.730 130.630 79.920 130.800 ;
        RECT 80.090 130.630 80.280 130.800 ;
        RECT 80.450 130.630 80.480 130.800 ;
        RECT 78.810 130.550 80.480 130.630 ;
      LAYER li1 ;
        RECT 81.210 130.550 81.480 132.710 ;
      LAYER li1 ;
        RECT 82.560 133.060 83.860 133.460 ;
        RECT 82.560 132.280 82.890 133.060 ;
        RECT 83.100 131.620 83.430 132.610 ;
        RECT 82.330 130.750 83.780 131.620 ;
        RECT 82.330 130.580 82.580 130.750 ;
        RECT 82.750 130.580 82.940 130.750 ;
        RECT 83.110 130.580 83.380 130.750 ;
        RECT 83.550 130.580 83.780 130.750 ;
        RECT 82.330 130.550 83.780 130.580 ;
      LAYER li1 ;
        RECT 85.090 130.550 85.340 133.810 ;
      LAYER li1 ;
        RECT 85.690 133.740 85.880 133.910 ;
        RECT 86.050 133.740 86.240 133.910 ;
        RECT 86.710 133.870 88.640 134.040 ;
        RECT 85.520 133.060 86.410 133.740 ;
        RECT 86.710 133.440 87.040 133.870 ;
        RECT 87.490 133.430 87.820 133.690 ;
        RECT 87.220 133.260 87.820 133.430 ;
        RECT 88.310 133.280 88.640 133.870 ;
        RECT 88.850 133.910 90.150 133.940 ;
        RECT 88.850 133.740 88.880 133.910 ;
        RECT 89.050 133.740 89.240 133.910 ;
        RECT 89.410 133.740 89.600 133.910 ;
        RECT 89.770 133.740 89.960 133.910 ;
        RECT 90.130 133.740 90.150 133.910 ;
        RECT 88.850 133.260 90.150 133.740 ;
        RECT 90.820 133.920 93.550 133.950 ;
        RECT 90.820 133.750 90.990 133.920 ;
        RECT 91.160 133.750 91.430 133.920 ;
        RECT 91.600 133.750 91.840 133.920 ;
        RECT 92.010 133.750 92.270 133.920 ;
        RECT 92.440 133.750 92.710 133.920 ;
        RECT 92.880 133.750 93.120 133.920 ;
        RECT 93.290 133.750 93.550 133.920 ;
        RECT 86.590 133.090 87.390 133.260 ;
        RECT 86.590 132.880 86.760 133.090 ;
      LAYER li1 ;
        RECT 88.000 133.080 88.670 133.100 ;
        RECT 87.570 132.910 89.840 133.080 ;
      LAYER li1 ;
        RECT 90.820 132.950 93.550 133.750 ;
        RECT 94.660 133.920 97.390 133.950 ;
        RECT 94.660 133.750 94.830 133.920 ;
        RECT 95.000 133.750 95.270 133.920 ;
        RECT 95.440 133.750 95.680 133.920 ;
        RECT 95.850 133.750 96.110 133.920 ;
        RECT 96.280 133.750 96.550 133.920 ;
        RECT 96.720 133.750 96.960 133.920 ;
        RECT 97.130 133.750 97.390 133.920 ;
        RECT 98.480 133.910 99.370 133.940 ;
        RECT 94.660 132.950 97.390 133.750 ;
        RECT 85.550 132.710 86.760 132.880 ;
      LAYER li1 ;
        RECT 86.940 132.740 87.740 132.910 ;
      LAYER li1 ;
        RECT 85.550 132.010 85.880 132.710 ;
      LAYER li1 ;
        RECT 86.940 132.530 87.110 132.740 ;
        RECT 89.510 132.730 89.840 132.910 ;
        RECT 86.380 132.250 87.110 132.530 ;
        RECT 87.290 132.190 87.720 132.560 ;
        RECT 87.920 132.190 88.210 132.730 ;
        RECT 88.450 132.400 89.160 132.730 ;
        RECT 89.430 132.560 89.840 132.730 ;
        RECT 89.510 132.290 89.840 132.560 ;
      LAYER li1 ;
        RECT 90.980 132.280 91.310 132.950 ;
        RECT 88.390 132.010 88.640 132.130 ;
        RECT 85.550 131.840 88.640 132.010 ;
        RECT 85.520 130.800 88.210 131.660 ;
        RECT 85.690 130.630 85.880 130.800 ;
        RECT 86.050 130.630 86.240 130.800 ;
        RECT 86.410 130.630 86.600 130.800 ;
        RECT 86.770 130.630 86.960 130.800 ;
        RECT 87.130 130.630 87.320 130.800 ;
        RECT 87.490 130.630 87.680 130.800 ;
        RECT 87.850 130.630 88.040 130.800 ;
        RECT 85.520 130.550 88.210 130.630 ;
        RECT 88.390 130.550 88.640 131.840 ;
        RECT 88.820 130.800 90.130 132.110 ;
        RECT 91.710 131.630 92.040 132.610 ;
        RECT 92.260 132.280 92.590 132.950 ;
        RECT 92.990 131.630 93.320 132.610 ;
        RECT 94.820 132.280 95.150 132.950 ;
        RECT 95.550 131.630 95.880 132.610 ;
        RECT 96.100 132.280 96.430 132.950 ;
        RECT 96.830 131.630 97.160 132.610 ;
        RECT 88.820 130.630 88.850 130.800 ;
        RECT 89.020 130.630 89.210 130.800 ;
        RECT 89.380 130.630 89.570 130.800 ;
        RECT 89.740 130.630 89.930 130.800 ;
        RECT 90.100 130.630 90.130 130.800 ;
        RECT 88.820 130.570 90.130 130.630 ;
        RECT 90.740 130.750 93.480 131.630 ;
        RECT 90.740 130.580 90.950 130.750 ;
        RECT 91.120 130.580 91.390 130.750 ;
        RECT 91.560 130.580 91.800 130.750 ;
        RECT 91.970 130.580 92.230 130.750 ;
        RECT 92.400 130.580 92.670 130.750 ;
        RECT 92.840 130.580 93.080 130.750 ;
        RECT 93.250 130.580 93.480 130.750 ;
        RECT 90.740 130.560 93.480 130.580 ;
        RECT 94.580 130.750 97.320 131.630 ;
        RECT 94.580 130.580 94.790 130.750 ;
        RECT 94.960 130.580 95.230 130.750 ;
        RECT 95.400 130.580 95.640 130.750 ;
        RECT 95.810 130.580 96.070 130.750 ;
        RECT 96.240 130.580 96.510 130.750 ;
        RECT 96.680 130.580 96.920 130.750 ;
        RECT 97.090 130.580 97.320 130.750 ;
        RECT 94.580 130.560 97.320 130.580 ;
      LAYER li1 ;
        RECT 98.050 130.550 98.300 133.810 ;
      LAYER li1 ;
        RECT 98.650 133.740 98.840 133.910 ;
        RECT 99.010 133.740 99.200 133.910 ;
        RECT 99.670 133.870 101.600 134.040 ;
        RECT 98.480 133.060 99.370 133.740 ;
        RECT 99.670 133.440 100.000 133.870 ;
        RECT 100.450 133.430 100.780 133.690 ;
        RECT 100.180 133.260 100.780 133.430 ;
        RECT 101.270 133.280 101.600 133.870 ;
        RECT 101.810 133.910 103.110 133.940 ;
        RECT 101.810 133.740 101.840 133.910 ;
        RECT 102.010 133.740 102.200 133.910 ;
        RECT 102.370 133.740 102.560 133.910 ;
        RECT 102.730 133.740 102.920 133.910 ;
        RECT 103.090 133.740 103.110 133.910 ;
        RECT 101.810 133.260 103.110 133.740 ;
        RECT 103.370 133.910 104.980 133.940 ;
        RECT 105.760 133.910 106.650 133.940 ;
        RECT 108.650 133.910 110.260 133.940 ;
        RECT 103.370 133.740 103.420 133.910 ;
        RECT 103.590 133.740 103.860 133.910 ;
        RECT 104.030 133.740 104.300 133.910 ;
        RECT 104.470 133.740 104.710 133.910 ;
        RECT 104.880 133.740 104.980 133.910 ;
        RECT 103.370 133.460 104.980 133.740 ;
        RECT 99.550 133.090 100.350 133.260 ;
        RECT 99.550 132.880 99.720 133.090 ;
      LAYER li1 ;
        RECT 100.960 133.080 101.630 133.100 ;
        RECT 100.530 132.910 102.800 133.080 ;
      LAYER li1 ;
        RECT 98.510 132.710 99.720 132.880 ;
      LAYER li1 ;
        RECT 99.900 132.740 100.700 132.910 ;
      LAYER li1 ;
        RECT 98.510 132.010 98.840 132.710 ;
      LAYER li1 ;
        RECT 99.900 132.530 100.070 132.740 ;
        RECT 102.470 132.730 102.800 132.910 ;
        RECT 99.340 132.250 100.070 132.530 ;
        RECT 100.250 132.190 100.680 132.560 ;
        RECT 100.880 132.190 101.170 132.730 ;
        RECT 101.410 132.400 102.120 132.730 ;
        RECT 102.390 132.560 102.800 132.730 ;
        RECT 102.470 132.290 102.800 132.560 ;
      LAYER li1 ;
        RECT 103.680 133.060 104.980 133.460 ;
        RECT 105.250 133.200 105.580 133.810 ;
        RECT 105.930 133.740 106.120 133.910 ;
        RECT 106.290 133.740 106.480 133.910 ;
        RECT 105.760 133.380 106.650 133.740 ;
        RECT 106.830 133.200 107.160 133.810 ;
        RECT 103.680 132.280 104.010 133.060 ;
        RECT 105.250 133.030 107.160 133.200 ;
        RECT 105.250 132.980 105.580 133.030 ;
      LAYER li1 ;
        RECT 107.610 132.850 107.940 133.810 ;
      LAYER li1 ;
        RECT 108.650 133.740 108.700 133.910 ;
        RECT 108.870 133.740 109.140 133.910 ;
        RECT 109.310 133.740 109.580 133.910 ;
        RECT 109.750 133.740 109.990 133.910 ;
        RECT 110.160 133.740 110.260 133.910 ;
        RECT 111.440 133.910 112.390 133.940 ;
        RECT 108.650 133.460 110.260 133.740 ;
        RECT 101.350 132.010 101.600 132.130 ;
        RECT 98.510 131.840 101.600 132.010 ;
        RECT 98.480 130.800 101.170 131.660 ;
        RECT 98.650 130.630 98.840 130.800 ;
        RECT 99.010 130.630 99.200 130.800 ;
        RECT 99.370 130.630 99.560 130.800 ;
        RECT 99.730 130.630 99.920 130.800 ;
        RECT 100.090 130.630 100.280 130.800 ;
        RECT 100.450 130.630 100.640 130.800 ;
        RECT 100.810 130.630 101.000 130.800 ;
        RECT 98.480 130.550 101.170 130.630 ;
        RECT 101.350 130.550 101.600 131.840 ;
        RECT 101.780 130.800 103.090 132.110 ;
        RECT 104.220 131.620 104.550 132.610 ;
      LAYER li1 ;
        RECT 105.250 132.470 105.980 132.800 ;
        RECT 106.190 132.550 106.920 132.800 ;
        RECT 107.100 132.680 107.940 132.850 ;
      LAYER li1 ;
        RECT 108.960 133.060 110.260 133.460 ;
      LAYER li1 ;
        RECT 107.100 132.370 107.270 132.680 ;
        RECT 106.690 132.200 107.270 132.370 ;
      LAYER li1 ;
        RECT 101.780 130.630 101.810 130.800 ;
        RECT 101.980 130.630 102.170 130.800 ;
        RECT 102.340 130.630 102.530 130.800 ;
        RECT 102.700 130.630 102.890 130.800 ;
        RECT 103.060 130.630 103.090 130.800 ;
        RECT 101.780 130.570 103.090 130.630 ;
        RECT 103.450 130.750 104.900 131.620 ;
        RECT 103.450 130.580 103.700 130.750 ;
        RECT 103.870 130.580 104.060 130.750 ;
        RECT 104.230 130.580 104.500 130.750 ;
        RECT 104.670 130.580 104.900 130.750 ;
        RECT 103.450 130.550 104.900 130.580 ;
        RECT 105.210 130.800 106.160 132.130 ;
        RECT 105.210 130.630 105.240 130.800 ;
        RECT 105.410 130.630 105.600 130.800 ;
        RECT 105.770 130.630 105.960 130.800 ;
        RECT 106.130 130.630 106.160 130.800 ;
        RECT 105.210 130.550 106.160 130.630 ;
      LAYER li1 ;
        RECT 106.690 130.550 107.160 132.200 ;
        RECT 107.450 132.190 108.360 132.500 ;
      LAYER li1 ;
        RECT 108.960 132.280 109.290 133.060 ;
        RECT 107.340 130.800 108.290 132.010 ;
        RECT 109.500 131.620 109.830 132.610 ;
        RECT 110.990 131.950 111.260 133.810 ;
        RECT 111.440 133.740 111.470 133.910 ;
        RECT 111.640 133.740 111.830 133.910 ;
        RECT 112.000 133.740 112.190 133.910 ;
        RECT 112.360 133.740 112.390 133.910 ;
        RECT 113.080 133.910 113.670 133.940 ;
        RECT 111.440 133.310 112.390 133.740 ;
        RECT 112.570 133.310 112.900 133.810 ;
      LAYER li1 ;
        RECT 111.440 132.160 111.770 133.130 ;
      LAYER li1 ;
        RECT 112.120 131.950 112.450 132.450 ;
        RECT 110.990 131.780 112.450 131.950 ;
        RECT 107.340 130.630 107.370 130.800 ;
        RECT 107.540 130.630 107.730 130.800 ;
        RECT 107.900 130.630 108.090 130.800 ;
        RECT 108.260 130.630 108.290 130.800 ;
        RECT 107.340 130.550 108.290 130.630 ;
        RECT 108.730 130.750 110.180 131.620 ;
        RECT 110.990 130.850 111.320 131.780 ;
        RECT 108.730 130.580 108.980 130.750 ;
        RECT 109.150 130.580 109.340 130.750 ;
        RECT 109.510 130.580 109.780 130.750 ;
        RECT 109.950 130.580 110.180 130.750 ;
        RECT 111.510 130.800 112.100 131.580 ;
        RECT 111.510 130.630 111.540 130.800 ;
        RECT 111.710 130.630 111.900 130.800 ;
        RECT 112.070 130.630 112.100 130.800 ;
        RECT 111.510 130.600 112.100 130.630 ;
        RECT 112.280 130.670 112.450 131.780 ;
        RECT 112.630 132.390 112.900 133.310 ;
        RECT 113.080 133.740 113.110 133.910 ;
        RECT 113.280 133.740 113.470 133.910 ;
        RECT 113.640 133.740 113.670 133.910 ;
        RECT 118.040 133.910 118.990 133.940 ;
        RECT 113.080 133.060 113.670 133.740 ;
      LAYER li1 ;
        RECT 113.950 133.680 116.890 133.850 ;
        RECT 113.950 133.470 114.120 133.680 ;
        RECT 113.910 133.300 114.120 133.470 ;
        RECT 113.950 132.690 114.120 133.300 ;
      LAYER li1 ;
        RECT 112.630 132.160 113.160 132.390 ;
        RECT 112.630 130.850 112.880 132.160 ;
      LAYER li1 ;
        RECT 113.580 131.820 114.120 132.690 ;
        RECT 114.300 132.200 114.630 133.500 ;
      LAYER li1 ;
        RECT 114.810 132.980 115.080 133.480 ;
        RECT 115.530 133.230 115.860 133.480 ;
        RECT 115.530 133.060 116.540 133.230 ;
        RECT 114.810 131.990 114.980 132.980 ;
        RECT 115.860 132.390 116.190 132.880 ;
        RECT 114.760 131.820 114.980 131.990 ;
        RECT 115.160 132.160 116.190 132.390 ;
        RECT 116.370 132.830 116.540 133.060 ;
      LAYER li1 ;
        RECT 116.720 133.180 116.890 133.680 ;
      LAYER li1 ;
        RECT 118.040 133.740 118.070 133.910 ;
        RECT 118.240 133.740 118.430 133.910 ;
        RECT 118.600 133.740 118.790 133.910 ;
        RECT 118.960 133.740 118.990 133.910 ;
        RECT 118.040 133.360 118.990 133.740 ;
      LAYER li1 ;
        RECT 119.170 133.870 121.830 134.040 ;
        RECT 119.170 133.180 119.340 133.870 ;
        RECT 116.720 133.010 119.340 133.180 ;
      LAYER li1 ;
        RECT 116.370 132.660 118.990 132.830 ;
        RECT 114.760 131.640 114.930 131.820 ;
        RECT 115.160 131.640 115.330 132.160 ;
        RECT 116.370 131.980 116.540 132.660 ;
      LAYER li1 ;
        RECT 119.170 132.480 119.340 133.010 ;
      LAYER li1 ;
        RECT 113.120 131.470 114.930 131.640 ;
        RECT 113.120 130.850 113.370 131.470 ;
        RECT 113.550 131.120 114.580 131.290 ;
        RECT 113.550 130.670 113.720 131.120 ;
        RECT 108.730 130.550 110.180 130.580 ;
        RECT 112.280 130.500 113.720 130.670 ;
        RECT 113.900 130.800 114.230 130.940 ;
        RECT 113.900 130.630 113.930 130.800 ;
        RECT 114.100 130.630 114.230 130.800 ;
        RECT 113.900 130.600 114.230 130.630 ;
        RECT 114.410 130.670 114.580 131.120 ;
        RECT 114.760 130.850 114.930 131.470 ;
        RECT 115.110 131.310 115.330 131.640 ;
        RECT 115.510 131.810 116.540 131.980 ;
        RECT 116.720 132.130 117.050 132.480 ;
      LAYER li1 ;
        RECT 117.490 132.310 119.340 132.480 ;
      LAYER li1 ;
        RECT 119.520 132.980 119.850 133.690 ;
        RECT 120.310 133.520 121.480 133.690 ;
        RECT 120.310 132.980 120.640 133.520 ;
        RECT 119.520 132.130 119.780 132.980 ;
        RECT 120.850 132.720 121.130 133.220 ;
        RECT 116.720 131.960 119.780 132.130 ;
        RECT 115.510 131.110 115.680 131.810 ;
        RECT 116.370 131.780 116.540 131.810 ;
        RECT 115.860 131.430 116.190 131.630 ;
        RECT 116.370 131.610 118.140 131.780 ;
        RECT 115.860 131.310 117.630 131.430 ;
        RECT 115.980 131.260 117.630 131.310 ;
        RECT 115.460 130.850 115.790 131.110 ;
        RECT 115.980 130.670 116.150 131.260 ;
        RECT 114.410 130.500 116.150 130.670 ;
        RECT 116.330 130.800 117.280 131.080 ;
        RECT 116.330 130.630 116.360 130.800 ;
        RECT 116.530 130.630 116.720 130.800 ;
        RECT 116.890 130.630 117.080 130.800 ;
        RECT 117.250 130.630 117.280 130.800 ;
        RECT 116.330 130.600 117.280 130.630 ;
        RECT 117.460 130.670 117.630 131.260 ;
        RECT 117.810 130.850 118.140 131.610 ;
        RECT 119.450 131.380 119.780 131.960 ;
        RECT 119.960 132.550 121.130 132.720 ;
        RECT 119.960 131.200 120.130 132.550 ;
        RECT 120.510 131.870 120.840 132.370 ;
        RECT 121.310 132.120 121.480 133.520 ;
      LAYER li1 ;
        RECT 121.660 133.210 121.830 133.870 ;
      LAYER li1 ;
        RECT 122.010 133.910 122.960 133.940 ;
        RECT 122.010 133.740 122.040 133.910 ;
        RECT 122.210 133.740 122.400 133.910 ;
        RECT 122.570 133.740 122.760 133.910 ;
        RECT 122.930 133.740 122.960 133.910 ;
        RECT 124.620 133.910 125.570 133.940 ;
        RECT 122.010 133.390 122.960 133.740 ;
        RECT 123.500 133.310 123.830 133.810 ;
        RECT 124.620 133.740 124.650 133.910 ;
        RECT 124.820 133.740 125.010 133.910 ;
        RECT 125.180 133.740 125.370 133.910 ;
        RECT 125.540 133.740 125.570 133.910 ;
      LAYER li1 ;
        RECT 121.660 133.040 122.670 133.210 ;
      LAYER li1 ;
        RECT 121.690 132.470 122.020 132.860 ;
      LAYER li1 ;
        RECT 122.340 132.650 122.670 133.040 ;
      LAYER li1 ;
        RECT 123.500 132.470 123.730 133.310 ;
        RECT 124.110 132.810 124.440 133.310 ;
        RECT 124.620 132.810 125.570 133.740 ;
        RECT 126.820 133.920 129.550 133.950 ;
        RECT 126.820 133.750 126.990 133.920 ;
        RECT 127.160 133.750 127.430 133.920 ;
        RECT 127.600 133.750 127.840 133.920 ;
        RECT 128.010 133.750 128.270 133.920 ;
        RECT 128.440 133.750 128.710 133.920 ;
        RECT 128.880 133.750 129.120 133.920 ;
        RECT 129.290 133.750 129.550 133.920 ;
        RECT 121.690 132.300 123.730 132.470 ;
        RECT 121.020 131.950 123.380 132.120 ;
        RECT 121.020 131.630 121.190 131.950 ;
        RECT 123.560 131.770 123.730 132.300 ;
        RECT 118.320 131.030 120.130 131.200 ;
        RECT 120.310 131.460 121.190 131.630 ;
        RECT 118.320 130.670 118.490 131.030 ;
        RECT 117.460 130.500 118.490 130.670 ;
        RECT 118.670 130.800 119.620 130.850 ;
        RECT 118.670 130.630 118.700 130.800 ;
        RECT 118.870 130.630 119.060 130.800 ;
        RECT 119.230 130.630 119.420 130.800 ;
        RECT 119.590 130.630 119.620 130.800 ;
        RECT 118.670 130.550 119.620 130.630 ;
        RECT 120.310 130.550 120.560 131.460 ;
        RECT 121.370 130.800 122.320 131.630 ;
        RECT 122.720 131.600 123.730 131.770 ;
        RECT 124.230 132.630 124.440 132.810 ;
        RECT 124.230 132.300 125.600 132.630 ;
        RECT 122.720 131.130 122.970 131.600 ;
        RECT 123.150 130.800 124.050 131.420 ;
        RECT 124.230 131.300 124.480 132.300 ;
        RECT 121.370 130.630 121.400 130.800 ;
        RECT 121.570 130.630 121.760 130.800 ;
        RECT 121.930 130.630 122.120 130.800 ;
        RECT 122.290 130.630 122.320 130.800 ;
        RECT 123.320 130.630 123.510 130.800 ;
        RECT 123.680 130.630 123.870 130.800 ;
        RECT 124.040 130.630 124.050 130.800 ;
        RECT 121.370 130.600 122.320 130.630 ;
        RECT 123.150 130.600 124.050 130.630 ;
        RECT 124.660 130.800 125.600 132.110 ;
        RECT 124.660 130.630 124.680 130.800 ;
        RECT 124.850 130.630 125.040 130.800 ;
        RECT 125.210 130.630 125.400 130.800 ;
        RECT 125.570 130.630 125.600 130.800 ;
        RECT 124.660 130.570 125.600 130.630 ;
      LAYER li1 ;
        RECT 125.780 130.570 126.120 133.640 ;
      LAYER li1 ;
        RECT 126.820 132.950 129.550 133.750 ;
        RECT 130.660 133.920 133.390 133.950 ;
        RECT 130.660 133.750 130.830 133.920 ;
        RECT 131.000 133.750 131.270 133.920 ;
        RECT 131.440 133.750 131.680 133.920 ;
        RECT 131.850 133.750 132.110 133.920 ;
        RECT 132.280 133.750 132.550 133.920 ;
        RECT 132.720 133.750 132.960 133.920 ;
        RECT 133.130 133.750 133.390 133.920 ;
        RECT 130.660 132.950 133.390 133.750 ;
        RECT 134.500 133.920 137.230 133.950 ;
        RECT 134.500 133.750 134.670 133.920 ;
        RECT 134.840 133.750 135.110 133.920 ;
        RECT 135.280 133.750 135.520 133.920 ;
        RECT 135.690 133.750 135.950 133.920 ;
        RECT 136.120 133.750 136.390 133.920 ;
        RECT 136.560 133.750 136.800 133.920 ;
        RECT 136.970 133.750 137.230 133.920 ;
        RECT 134.500 132.950 137.230 133.750 ;
        RECT 138.340 133.920 141.070 133.950 ;
        RECT 138.340 133.750 138.510 133.920 ;
        RECT 138.680 133.750 138.950 133.920 ;
        RECT 139.120 133.750 139.360 133.920 ;
        RECT 139.530 133.750 139.790 133.920 ;
        RECT 139.960 133.750 140.230 133.920 ;
        RECT 140.400 133.750 140.640 133.920 ;
        RECT 140.810 133.750 141.070 133.920 ;
        RECT 138.340 132.950 141.070 133.750 ;
        RECT 126.980 132.280 127.310 132.950 ;
        RECT 127.710 131.630 128.040 132.610 ;
        RECT 128.260 132.280 128.590 132.950 ;
        RECT 128.990 131.630 129.320 132.610 ;
        RECT 130.820 132.280 131.150 132.950 ;
        RECT 131.550 131.630 131.880 132.610 ;
        RECT 132.100 132.280 132.430 132.950 ;
        RECT 132.830 131.630 133.160 132.610 ;
        RECT 134.660 132.280 134.990 132.950 ;
        RECT 135.390 131.630 135.720 132.610 ;
        RECT 135.940 132.280 136.270 132.950 ;
        RECT 136.670 131.630 137.000 132.610 ;
        RECT 138.500 132.280 138.830 132.950 ;
        RECT 139.230 131.630 139.560 132.610 ;
        RECT 139.780 132.280 140.110 132.950 ;
        RECT 140.510 131.630 140.840 132.610 ;
        RECT 126.740 130.750 129.480 131.630 ;
        RECT 126.740 130.580 126.950 130.750 ;
        RECT 127.120 130.580 127.390 130.750 ;
        RECT 127.560 130.580 127.800 130.750 ;
        RECT 127.970 130.580 128.230 130.750 ;
        RECT 128.400 130.580 128.670 130.750 ;
        RECT 128.840 130.580 129.080 130.750 ;
        RECT 129.250 130.580 129.480 130.750 ;
        RECT 126.740 130.560 129.480 130.580 ;
        RECT 130.580 130.750 133.320 131.630 ;
        RECT 130.580 130.580 130.790 130.750 ;
        RECT 130.960 130.580 131.230 130.750 ;
        RECT 131.400 130.580 131.640 130.750 ;
        RECT 131.810 130.580 132.070 130.750 ;
        RECT 132.240 130.580 132.510 130.750 ;
        RECT 132.680 130.580 132.920 130.750 ;
        RECT 133.090 130.580 133.320 130.750 ;
        RECT 130.580 130.560 133.320 130.580 ;
        RECT 134.420 130.750 137.160 131.630 ;
        RECT 134.420 130.580 134.630 130.750 ;
        RECT 134.800 130.580 135.070 130.750 ;
        RECT 135.240 130.580 135.480 130.750 ;
        RECT 135.650 130.580 135.910 130.750 ;
        RECT 136.080 130.580 136.350 130.750 ;
        RECT 136.520 130.580 136.760 130.750 ;
        RECT 136.930 130.580 137.160 130.750 ;
        RECT 134.420 130.560 137.160 130.580 ;
        RECT 138.260 130.750 141.000 131.630 ;
        RECT 138.260 130.580 138.470 130.750 ;
        RECT 138.640 130.580 138.910 130.750 ;
        RECT 139.080 130.580 139.320 130.750 ;
        RECT 139.490 130.580 139.750 130.750 ;
        RECT 139.920 130.580 140.190 130.750 ;
        RECT 140.360 130.580 140.600 130.750 ;
        RECT 140.770 130.580 141.000 130.750 ;
        RECT 138.260 130.560 141.000 130.580 ;
        RECT 5.760 130.150 5.920 130.330 ;
        RECT 6.090 130.150 6.400 130.330 ;
        RECT 6.570 130.150 6.880 130.330 ;
        RECT 7.050 130.150 7.360 130.330 ;
        RECT 7.530 130.150 7.840 130.330 ;
        RECT 8.010 130.150 8.320 130.330 ;
        RECT 8.490 130.150 8.800 130.330 ;
        RECT 8.970 130.150 9.280 130.330 ;
        RECT 9.450 130.150 9.760 130.330 ;
        RECT 9.930 130.150 10.240 130.330 ;
        RECT 10.410 130.150 10.720 130.330 ;
        RECT 10.890 130.150 11.200 130.330 ;
        RECT 11.370 130.150 11.680 130.330 ;
        RECT 11.850 130.150 12.160 130.330 ;
        RECT 12.330 130.150 12.640 130.330 ;
        RECT 12.810 130.150 13.120 130.330 ;
        RECT 13.290 130.150 13.600 130.330 ;
        RECT 13.770 130.150 14.080 130.330 ;
        RECT 14.250 130.150 14.560 130.330 ;
        RECT 14.730 130.150 15.040 130.330 ;
        RECT 15.210 130.150 15.520 130.330 ;
        RECT 15.690 130.150 16.000 130.330 ;
        RECT 16.170 130.150 16.480 130.330 ;
        RECT 16.650 130.150 16.960 130.330 ;
        RECT 17.130 130.150 17.440 130.330 ;
        RECT 17.610 130.150 17.920 130.330 ;
        RECT 18.090 130.150 18.400 130.330 ;
        RECT 18.570 130.150 18.880 130.330 ;
        RECT 19.050 130.150 19.360 130.330 ;
        RECT 19.530 130.150 19.840 130.330 ;
        RECT 20.010 130.150 20.320 130.330 ;
        RECT 20.490 130.150 20.800 130.330 ;
        RECT 20.970 130.150 21.280 130.330 ;
        RECT 21.450 130.150 21.760 130.330 ;
        RECT 21.930 130.150 22.240 130.330 ;
        RECT 22.410 130.150 22.720 130.330 ;
        RECT 22.890 130.150 23.200 130.330 ;
        RECT 23.370 130.150 23.680 130.330 ;
        RECT 23.850 130.150 24.160 130.330 ;
        RECT 24.330 130.150 24.640 130.330 ;
        RECT 24.810 130.150 25.120 130.330 ;
        RECT 25.290 130.150 25.600 130.330 ;
        RECT 25.770 130.150 26.080 130.330 ;
        RECT 26.250 130.150 26.560 130.330 ;
        RECT 26.730 130.150 27.040 130.330 ;
        RECT 27.210 130.150 27.520 130.330 ;
        RECT 27.690 130.150 28.000 130.330 ;
        RECT 28.170 130.150 28.480 130.330 ;
        RECT 28.650 130.150 28.960 130.330 ;
        RECT 29.130 130.150 29.440 130.330 ;
        RECT 29.610 130.150 29.920 130.330 ;
        RECT 30.090 130.150 30.400 130.330 ;
        RECT 30.570 130.150 30.880 130.330 ;
        RECT 31.050 130.320 31.360 130.330 ;
        RECT 31.530 130.320 31.840 130.330 ;
        RECT 31.050 130.150 31.200 130.320 ;
        RECT 31.680 130.150 31.840 130.320 ;
        RECT 32.010 130.150 32.320 130.330 ;
        RECT 32.490 130.150 32.800 130.330 ;
        RECT 32.970 130.150 33.280 130.330 ;
        RECT 33.450 130.150 33.760 130.330 ;
        RECT 33.930 130.320 34.080 130.330 ;
        RECT 34.560 130.320 34.720 130.330 ;
        RECT 33.930 130.150 34.240 130.320 ;
        RECT 34.410 130.150 34.720 130.320 ;
        RECT 34.890 130.150 35.200 130.330 ;
        RECT 35.370 130.150 35.680 130.330 ;
        RECT 35.850 130.150 36.160 130.330 ;
        RECT 36.330 130.150 36.640 130.330 ;
        RECT 36.810 130.150 37.120 130.330 ;
        RECT 37.290 130.150 37.600 130.330 ;
        RECT 37.770 130.150 38.080 130.330 ;
        RECT 38.250 130.150 38.560 130.330 ;
        RECT 38.730 130.150 39.040 130.330 ;
        RECT 39.210 130.150 39.520 130.330 ;
        RECT 39.690 130.150 40.000 130.330 ;
        RECT 40.170 130.150 40.480 130.330 ;
        RECT 40.650 130.150 40.960 130.330 ;
        RECT 41.130 130.150 41.440 130.330 ;
        RECT 41.610 130.150 41.920 130.330 ;
        RECT 42.090 130.150 42.400 130.330 ;
        RECT 42.570 130.150 42.880 130.330 ;
        RECT 43.050 130.150 43.360 130.330 ;
        RECT 43.530 130.320 43.680 130.330 ;
        RECT 44.160 130.320 44.320 130.330 ;
        RECT 43.530 130.150 43.840 130.320 ;
        RECT 44.010 130.150 44.320 130.320 ;
        RECT 44.490 130.150 44.800 130.330 ;
        RECT 44.970 130.150 45.280 130.330 ;
        RECT 45.450 130.150 45.760 130.330 ;
        RECT 45.930 130.150 46.240 130.330 ;
        RECT 46.410 130.150 46.720 130.330 ;
        RECT 46.890 130.150 47.200 130.330 ;
        RECT 47.370 130.150 47.680 130.330 ;
        RECT 47.850 130.150 48.160 130.330 ;
        RECT 48.330 130.150 48.640 130.330 ;
        RECT 48.810 130.150 49.120 130.330 ;
        RECT 49.290 130.150 49.600 130.330 ;
        RECT 49.770 130.150 50.080 130.330 ;
        RECT 50.250 130.150 50.560 130.330 ;
        RECT 50.730 130.150 51.040 130.330 ;
        RECT 51.210 130.150 51.520 130.330 ;
        RECT 51.690 130.150 52.000 130.330 ;
        RECT 52.170 130.150 52.480 130.330 ;
        RECT 52.650 130.150 52.960 130.330 ;
        RECT 53.130 130.150 53.440 130.330 ;
        RECT 53.610 130.150 53.920 130.330 ;
        RECT 54.090 130.150 54.400 130.330 ;
        RECT 54.570 130.150 54.880 130.330 ;
        RECT 55.050 130.150 55.360 130.330 ;
        RECT 55.530 130.150 55.840 130.330 ;
        RECT 56.010 130.150 56.320 130.330 ;
        RECT 56.490 130.150 56.800 130.330 ;
        RECT 56.970 130.150 57.280 130.330 ;
        RECT 57.450 130.150 57.760 130.330 ;
        RECT 57.930 130.150 58.240 130.330 ;
        RECT 58.410 130.150 58.720 130.330 ;
        RECT 58.890 130.150 59.200 130.330 ;
        RECT 59.370 130.150 59.680 130.330 ;
        RECT 59.850 130.150 60.160 130.330 ;
        RECT 60.330 130.150 60.640 130.330 ;
        RECT 60.810 130.150 61.120 130.330 ;
        RECT 61.290 130.150 61.600 130.330 ;
        RECT 61.770 130.150 62.080 130.330 ;
        RECT 62.250 130.150 62.560 130.330 ;
        RECT 62.730 130.150 63.040 130.330 ;
        RECT 63.210 130.150 63.520 130.330 ;
        RECT 63.690 130.150 64.000 130.330 ;
        RECT 64.170 130.150 64.480 130.330 ;
        RECT 64.650 130.150 64.960 130.330 ;
        RECT 65.130 130.150 65.440 130.330 ;
        RECT 65.610 130.150 65.920 130.330 ;
        RECT 66.090 130.150 66.400 130.330 ;
        RECT 66.570 130.150 66.880 130.330 ;
        RECT 67.050 130.150 67.360 130.330 ;
        RECT 67.530 130.150 67.840 130.330 ;
        RECT 68.010 130.150 68.320 130.330 ;
        RECT 68.490 130.150 68.800 130.330 ;
        RECT 68.970 130.150 69.280 130.330 ;
        RECT 69.450 130.150 69.760 130.330 ;
        RECT 69.930 130.150 70.240 130.330 ;
        RECT 70.410 130.150 70.720 130.330 ;
        RECT 70.890 130.150 71.200 130.330 ;
        RECT 71.370 130.150 71.680 130.330 ;
        RECT 71.850 130.150 72.160 130.330 ;
        RECT 72.330 130.150 72.640 130.330 ;
        RECT 72.810 130.320 73.120 130.330 ;
        RECT 73.290 130.320 73.600 130.330 ;
        RECT 72.810 130.150 72.960 130.320 ;
        RECT 73.440 130.150 73.600 130.320 ;
        RECT 73.770 130.320 73.920 130.330 ;
        RECT 74.400 130.320 74.560 130.330 ;
        RECT 73.770 130.150 74.080 130.320 ;
        RECT 74.250 130.150 74.560 130.320 ;
        RECT 74.730 130.150 75.040 130.330 ;
        RECT 75.210 130.150 75.520 130.330 ;
        RECT 75.690 130.150 76.000 130.330 ;
        RECT 76.170 130.150 76.480 130.330 ;
        RECT 76.650 130.150 76.960 130.330 ;
        RECT 77.130 130.150 77.440 130.330 ;
        RECT 77.610 130.150 77.920 130.330 ;
        RECT 78.090 130.150 78.400 130.330 ;
        RECT 78.570 130.150 78.880 130.330 ;
        RECT 79.050 130.150 79.360 130.330 ;
        RECT 79.530 130.150 79.840 130.330 ;
        RECT 80.010 130.150 80.320 130.330 ;
        RECT 80.490 130.150 80.800 130.330 ;
        RECT 80.970 130.150 81.280 130.330 ;
        RECT 81.450 130.150 81.760 130.330 ;
        RECT 81.930 130.150 82.240 130.330 ;
        RECT 82.410 130.150 82.720 130.330 ;
        RECT 82.890 130.150 83.200 130.330 ;
        RECT 83.370 130.150 83.680 130.330 ;
        RECT 83.850 130.150 84.160 130.330 ;
        RECT 84.330 130.150 84.640 130.330 ;
        RECT 84.810 130.150 85.120 130.330 ;
        RECT 85.290 130.150 85.600 130.330 ;
        RECT 85.770 130.150 86.080 130.330 ;
        RECT 86.250 130.150 86.560 130.330 ;
        RECT 86.730 130.150 87.040 130.330 ;
        RECT 87.210 130.150 87.520 130.330 ;
        RECT 87.690 130.150 88.000 130.330 ;
        RECT 88.170 130.150 88.480 130.330 ;
        RECT 88.650 130.150 88.960 130.330 ;
        RECT 89.130 130.150 89.440 130.330 ;
        RECT 89.610 130.150 89.920 130.330 ;
        RECT 90.090 130.150 90.400 130.330 ;
        RECT 90.570 130.150 90.880 130.330 ;
        RECT 91.050 130.150 91.360 130.330 ;
        RECT 91.530 130.150 91.840 130.330 ;
        RECT 92.010 130.150 92.320 130.330 ;
        RECT 92.490 130.150 92.800 130.330 ;
        RECT 92.970 130.150 93.280 130.330 ;
        RECT 93.450 130.150 93.760 130.330 ;
        RECT 93.930 130.150 94.240 130.330 ;
        RECT 94.410 130.150 94.720 130.330 ;
        RECT 94.890 130.150 95.200 130.330 ;
        RECT 95.370 130.150 95.680 130.330 ;
        RECT 95.850 130.150 96.160 130.330 ;
        RECT 96.330 130.150 96.640 130.330 ;
        RECT 96.810 130.150 97.120 130.330 ;
        RECT 97.290 130.150 97.600 130.330 ;
        RECT 97.770 130.150 98.080 130.330 ;
        RECT 98.250 130.150 98.560 130.330 ;
        RECT 98.730 130.150 99.040 130.330 ;
        RECT 99.210 130.150 99.520 130.330 ;
        RECT 99.690 130.150 100.000 130.330 ;
        RECT 100.170 130.150 100.480 130.330 ;
        RECT 100.650 130.150 100.960 130.330 ;
        RECT 101.130 130.150 101.440 130.330 ;
        RECT 101.610 130.150 101.920 130.330 ;
        RECT 102.090 130.150 102.400 130.330 ;
        RECT 102.570 130.150 102.880 130.330 ;
        RECT 103.050 130.150 103.360 130.330 ;
        RECT 103.530 130.150 103.840 130.330 ;
        RECT 104.010 130.150 104.320 130.330 ;
        RECT 104.490 130.150 104.800 130.330 ;
        RECT 104.970 130.150 105.280 130.330 ;
        RECT 105.450 130.150 105.760 130.330 ;
        RECT 105.930 130.150 106.240 130.330 ;
        RECT 106.410 130.150 106.720 130.330 ;
        RECT 106.890 130.150 107.200 130.330 ;
        RECT 107.370 130.150 107.680 130.330 ;
        RECT 107.850 130.150 108.160 130.330 ;
        RECT 108.330 130.150 108.640 130.330 ;
        RECT 108.810 130.150 109.120 130.330 ;
        RECT 109.290 130.150 109.600 130.330 ;
        RECT 109.770 130.150 110.080 130.330 ;
        RECT 110.250 130.150 110.400 130.330 ;
        RECT 110.880 130.150 111.040 130.330 ;
        RECT 111.210 130.150 111.520 130.330 ;
        RECT 111.690 130.150 112.000 130.330 ;
        RECT 112.170 130.150 112.480 130.330 ;
        RECT 112.650 130.150 112.960 130.330 ;
        RECT 113.130 130.150 113.440 130.330 ;
        RECT 113.610 130.150 113.920 130.330 ;
        RECT 114.090 130.150 114.400 130.330 ;
        RECT 114.570 130.150 114.880 130.330 ;
        RECT 115.050 130.150 115.360 130.330 ;
        RECT 115.530 130.150 115.840 130.330 ;
        RECT 116.010 130.150 116.320 130.330 ;
        RECT 116.490 130.150 116.800 130.330 ;
        RECT 116.970 130.150 117.280 130.330 ;
        RECT 117.450 130.150 117.760 130.330 ;
        RECT 117.930 130.320 118.080 130.330 ;
        RECT 118.560 130.320 118.720 130.330 ;
        RECT 117.930 130.150 118.240 130.320 ;
        RECT 118.410 130.150 118.720 130.320 ;
        RECT 118.890 130.150 119.200 130.330 ;
        RECT 119.370 130.150 119.680 130.330 ;
        RECT 119.850 130.150 120.160 130.330 ;
        RECT 120.330 130.150 120.640 130.330 ;
        RECT 120.810 130.150 121.120 130.330 ;
        RECT 121.290 130.150 121.600 130.330 ;
        RECT 121.770 130.150 122.080 130.330 ;
        RECT 122.250 130.150 122.560 130.330 ;
        RECT 122.730 130.150 123.040 130.330 ;
        RECT 123.210 130.150 123.520 130.330 ;
        RECT 123.690 130.150 124.000 130.330 ;
        RECT 124.170 130.150 124.480 130.330 ;
        RECT 124.650 130.150 124.960 130.330 ;
        RECT 125.130 130.150 125.440 130.330 ;
        RECT 125.610 130.150 125.920 130.330 ;
        RECT 126.090 130.150 126.400 130.330 ;
        RECT 126.570 130.150 126.880 130.330 ;
        RECT 127.050 130.150 127.360 130.330 ;
        RECT 127.530 130.150 127.840 130.330 ;
        RECT 128.010 130.150 128.320 130.330 ;
        RECT 128.490 130.150 128.800 130.330 ;
        RECT 128.970 130.150 129.280 130.330 ;
        RECT 129.450 130.150 129.760 130.330 ;
        RECT 129.930 130.150 130.240 130.330 ;
        RECT 130.410 130.150 130.720 130.330 ;
        RECT 130.890 130.150 131.200 130.330 ;
        RECT 131.370 130.150 131.680 130.330 ;
        RECT 131.850 130.150 132.160 130.330 ;
        RECT 132.330 130.150 132.640 130.330 ;
        RECT 132.810 130.150 133.120 130.330 ;
        RECT 133.290 130.150 133.600 130.330 ;
        RECT 133.770 130.150 134.080 130.330 ;
        RECT 134.250 130.150 134.560 130.330 ;
        RECT 134.730 130.150 135.040 130.330 ;
        RECT 135.210 130.150 135.520 130.330 ;
        RECT 135.690 130.150 136.000 130.330 ;
        RECT 136.170 130.150 136.480 130.330 ;
        RECT 136.650 130.150 136.960 130.330 ;
        RECT 137.130 130.150 137.440 130.330 ;
        RECT 137.610 130.150 137.920 130.330 ;
        RECT 138.090 130.150 138.400 130.330 ;
        RECT 138.570 130.150 138.880 130.330 ;
        RECT 139.050 130.150 139.360 130.330 ;
        RECT 139.530 130.150 139.840 130.330 ;
        RECT 140.010 130.150 140.320 130.330 ;
        RECT 140.490 130.150 140.800 130.330 ;
        RECT 140.970 130.150 141.280 130.330 ;
        RECT 141.450 130.320 141.760 130.330 ;
        RECT 141.930 130.320 142.080 130.330 ;
        RECT 141.450 130.150 141.600 130.320 ;
        RECT 6.260 129.900 9.000 129.920 ;
        RECT 6.260 129.730 6.470 129.900 ;
        RECT 6.640 129.730 6.910 129.900 ;
        RECT 7.080 129.730 7.320 129.900 ;
        RECT 7.490 129.730 7.750 129.900 ;
        RECT 7.920 129.730 8.190 129.900 ;
        RECT 8.360 129.730 8.600 129.900 ;
        RECT 8.770 129.730 9.000 129.900 ;
        RECT 6.260 128.850 9.000 129.730 ;
        RECT 10.100 129.900 12.840 129.920 ;
        RECT 10.100 129.730 10.310 129.900 ;
        RECT 10.480 129.730 10.750 129.900 ;
        RECT 10.920 129.730 11.160 129.900 ;
        RECT 11.330 129.730 11.590 129.900 ;
        RECT 11.760 129.730 12.030 129.900 ;
        RECT 12.200 129.730 12.440 129.900 ;
        RECT 12.610 129.730 12.840 129.900 ;
        RECT 10.100 128.850 12.840 129.730 ;
        RECT 13.690 129.900 15.140 129.930 ;
        RECT 13.690 129.730 13.940 129.900 ;
        RECT 14.110 129.730 14.300 129.900 ;
        RECT 14.470 129.730 14.740 129.900 ;
        RECT 14.910 129.730 15.140 129.900 ;
        RECT 13.690 128.860 15.140 129.730 ;
        RECT 6.500 127.530 6.830 128.200 ;
        RECT 7.230 127.870 7.560 128.850 ;
        RECT 7.780 127.530 8.110 128.200 ;
        RECT 8.510 127.870 8.840 128.850 ;
        RECT 10.340 127.530 10.670 128.200 ;
        RECT 11.070 127.870 11.400 128.850 ;
        RECT 11.620 127.530 11.950 128.200 ;
        RECT 12.350 127.870 12.680 128.850 ;
        RECT 6.340 126.530 9.070 127.530 ;
        RECT 10.180 126.530 12.910 127.530 ;
        RECT 13.920 127.420 14.250 128.200 ;
        RECT 14.460 127.870 14.790 128.860 ;
      LAYER li1 ;
        RECT 15.480 128.350 15.910 129.930 ;
      LAYER li1 ;
        RECT 16.090 129.850 16.650 129.930 ;
        RECT 16.090 129.680 16.100 129.850 ;
        RECT 16.270 129.680 16.460 129.850 ;
        RECT 16.630 129.680 16.650 129.850 ;
        RECT 16.090 128.350 16.650 129.680 ;
        RECT 18.260 129.900 21.000 129.920 ;
        RECT 18.260 129.730 18.470 129.900 ;
        RECT 18.640 129.730 18.910 129.900 ;
        RECT 19.080 129.730 19.320 129.900 ;
        RECT 19.490 129.730 19.750 129.900 ;
        RECT 19.920 129.730 20.190 129.900 ;
        RECT 20.360 129.730 20.600 129.900 ;
        RECT 20.770 129.730 21.000 129.900 ;
        RECT 13.920 127.020 15.220 127.420 ;
        RECT 13.610 126.540 15.220 127.020 ;
      LAYER li1 ;
        RECT 15.480 126.670 15.730 128.350 ;
      LAYER li1 ;
        RECT 16.040 127.460 16.370 127.920 ;
      LAYER li1 ;
        RECT 16.830 127.640 17.160 129.430 ;
      LAYER li1 ;
        RECT 17.340 127.460 17.590 129.180 ;
        RECT 18.260 128.850 21.000 129.730 ;
        RECT 22.100 129.900 24.840 129.920 ;
        RECT 22.100 129.730 22.310 129.900 ;
        RECT 22.480 129.730 22.750 129.900 ;
        RECT 22.920 129.730 23.160 129.900 ;
        RECT 23.330 129.730 23.590 129.900 ;
        RECT 23.760 129.730 24.030 129.900 ;
        RECT 24.200 129.730 24.440 129.900 ;
        RECT 24.610 129.730 24.840 129.900 ;
        RECT 22.100 128.850 24.840 129.730 ;
        RECT 25.940 129.900 28.680 129.920 ;
        RECT 25.940 129.730 26.150 129.900 ;
        RECT 26.320 129.730 26.590 129.900 ;
        RECT 26.760 129.730 27.000 129.900 ;
        RECT 27.170 129.730 27.430 129.900 ;
        RECT 27.600 129.730 27.870 129.900 ;
        RECT 28.040 129.730 28.280 129.900 ;
        RECT 28.450 129.730 28.680 129.900 ;
        RECT 25.940 128.850 28.680 129.730 ;
        RECT 29.780 129.900 32.520 129.920 ;
        RECT 29.780 129.730 29.990 129.900 ;
        RECT 30.160 129.730 30.430 129.900 ;
        RECT 30.600 129.730 30.840 129.900 ;
        RECT 31.010 129.730 31.270 129.900 ;
        RECT 31.440 129.730 31.710 129.900 ;
        RECT 31.880 129.730 32.120 129.900 ;
        RECT 32.290 129.730 32.520 129.900 ;
        RECT 29.780 128.850 32.520 129.730 ;
        RECT 18.500 127.530 18.830 128.200 ;
        RECT 19.230 127.870 19.560 128.850 ;
        RECT 19.780 127.530 20.110 128.200 ;
        RECT 20.510 127.870 20.840 128.850 ;
        RECT 22.340 127.530 22.670 128.200 ;
        RECT 23.070 127.870 23.400 128.850 ;
        RECT 23.620 127.530 23.950 128.200 ;
        RECT 24.350 127.870 24.680 128.850 ;
        RECT 26.180 127.530 26.510 128.200 ;
        RECT 26.910 127.870 27.240 128.850 ;
        RECT 27.460 127.530 27.790 128.200 ;
        RECT 28.190 127.870 28.520 128.850 ;
        RECT 30.020 127.530 30.350 128.200 ;
        RECT 30.750 127.870 31.080 128.850 ;
        RECT 31.300 127.530 31.630 128.200 ;
        RECT 32.030 127.870 32.360 128.850 ;
        RECT 16.040 127.290 17.590 127.460 ;
        RECT 15.910 126.540 17.160 127.110 ;
        RECT 17.340 126.670 17.590 127.290 ;
        RECT 18.340 126.530 21.070 127.530 ;
        RECT 22.180 126.530 24.910 127.530 ;
        RECT 26.020 126.530 28.750 127.530 ;
        RECT 29.860 126.530 32.590 127.530 ;
      LAYER li1 ;
        RECT 34.670 126.670 34.940 129.930 ;
      LAYER li1 ;
        RECT 35.120 129.850 36.020 129.930 ;
        RECT 35.120 129.680 35.130 129.850 ;
        RECT 35.300 129.680 35.490 129.850 ;
        RECT 35.660 129.680 35.850 129.850 ;
        RECT 36.200 129.810 38.090 129.980 ;
        RECT 35.120 128.350 36.020 129.680 ;
        RECT 36.200 128.350 36.370 129.810 ;
      LAYER li1 ;
        RECT 36.550 127.950 36.880 129.430 ;
      LAYER li1 ;
        RECT 35.150 127.770 35.480 127.930 ;
        RECT 37.060 127.770 37.390 129.630 ;
        RECT 37.840 128.270 38.090 129.810 ;
        RECT 38.270 129.850 39.220 129.930 ;
        RECT 38.270 129.680 38.300 129.850 ;
        RECT 38.470 129.680 38.660 129.850 ;
        RECT 38.830 129.680 39.020 129.850 ;
        RECT 39.190 129.680 39.220 129.850 ;
        RECT 38.270 128.450 39.220 129.680 ;
        RECT 39.400 128.270 39.730 129.910 ;
        RECT 40.340 129.900 43.080 129.920 ;
        RECT 40.340 129.730 40.550 129.900 ;
        RECT 40.720 129.730 40.990 129.900 ;
        RECT 41.160 129.730 41.400 129.900 ;
        RECT 41.570 129.730 41.830 129.900 ;
        RECT 42.000 129.730 42.270 129.900 ;
        RECT 42.440 129.730 42.680 129.900 ;
        RECT 42.850 129.730 43.080 129.900 ;
        RECT 40.340 128.850 43.080 129.730 ;
        RECT 44.250 129.850 45.510 129.930 ;
        RECT 44.250 129.680 44.260 129.850 ;
        RECT 44.430 129.680 44.620 129.850 ;
        RECT 44.790 129.680 44.980 129.850 ;
        RECT 45.150 129.680 45.340 129.850 ;
        RECT 37.840 128.100 39.730 128.270 ;
        RECT 35.150 127.600 37.420 127.770 ;
        RECT 35.110 126.540 36.820 127.420 ;
        RECT 37.250 126.800 37.420 127.600 ;
      LAYER li1 ;
        RECT 37.600 127.180 37.770 127.920 ;
        RECT 39.390 127.680 39.720 127.920 ;
      LAYER li1 ;
        RECT 40.580 127.530 40.910 128.200 ;
        RECT 41.310 127.870 41.640 128.850 ;
        RECT 41.860 127.530 42.190 128.200 ;
        RECT 42.590 127.870 42.920 128.850 ;
        RECT 44.250 128.450 45.510 129.680 ;
      LAYER li1 ;
        RECT 46.040 129.430 46.210 129.930 ;
        RECT 45.690 128.350 46.210 129.430 ;
      LAYER li1 ;
        RECT 46.470 129.850 47.780 129.930 ;
        RECT 46.470 129.680 46.500 129.850 ;
        RECT 46.670 129.680 46.860 129.850 ;
        RECT 47.030 129.680 47.220 129.850 ;
        RECT 47.390 129.680 47.580 129.850 ;
        RECT 47.750 129.680 47.780 129.850 ;
        RECT 46.470 128.470 47.780 129.680 ;
        RECT 48.250 129.900 49.700 129.930 ;
        RECT 48.250 129.730 48.500 129.900 ;
        RECT 48.670 129.730 48.860 129.900 ;
        RECT 49.030 129.730 49.300 129.900 ;
        RECT 49.470 129.730 49.700 129.900 ;
        RECT 48.250 128.860 49.700 129.730 ;
      LAYER li1 ;
        RECT 45.690 128.270 45.960 128.350 ;
        RECT 44.900 128.100 45.960 128.270 ;
        RECT 44.290 127.710 44.710 128.040 ;
        RECT 44.900 127.530 45.070 128.100 ;
        RECT 46.410 127.980 46.920 128.290 ;
        RECT 47.170 127.980 47.880 128.290 ;
        RECT 45.250 127.710 45.760 127.920 ;
      LAYER li1 ;
        RECT 45.960 127.630 47.830 127.800 ;
      LAYER li1 ;
        RECT 37.590 127.010 37.770 127.180 ;
        RECT 37.600 126.980 37.770 127.010 ;
      LAYER li1 ;
        RECT 37.950 126.800 38.200 127.500 ;
        RECT 37.250 126.630 38.200 126.800 ;
        RECT 38.380 126.540 39.690 127.500 ;
        RECT 40.420 126.530 43.150 127.530 ;
        RECT 44.320 126.610 44.650 127.530 ;
      LAYER li1 ;
        RECT 44.900 126.790 45.430 127.530 ;
      LAYER li1 ;
        RECT 45.960 126.610 46.130 127.630 ;
        RECT 44.320 126.440 46.130 126.610 ;
        RECT 46.310 126.540 47.410 127.450 ;
        RECT 47.580 126.700 47.830 127.630 ;
        RECT 48.480 127.420 48.810 128.200 ;
        RECT 49.020 127.870 49.350 128.860 ;
        RECT 50.040 127.640 50.290 129.910 ;
        RECT 50.470 129.850 51.420 129.930 ;
        RECT 50.470 129.680 50.500 129.850 ;
        RECT 50.670 129.680 50.860 129.850 ;
        RECT 51.030 129.680 51.220 129.850 ;
        RECT 51.390 129.680 51.420 129.850 ;
        RECT 50.470 129.100 51.420 129.680 ;
        RECT 51.600 129.120 51.930 129.910 ;
        RECT 51.610 128.620 51.930 129.120 ;
        RECT 52.160 129.850 52.410 129.880 ;
        RECT 52.160 129.680 52.190 129.850 ;
        RECT 52.360 129.680 52.410 129.850 ;
        RECT 52.160 128.800 52.410 129.680 ;
        RECT 52.590 128.620 52.760 129.930 ;
        RECT 55.530 129.850 55.860 129.880 ;
        RECT 51.610 128.450 52.760 128.620 ;
        RECT 52.940 129.460 54.930 129.790 ;
        RECT 51.100 127.640 51.430 128.070 ;
        RECT 50.040 127.470 51.430 127.640 ;
        RECT 48.480 127.020 49.780 127.420 ;
        RECT 48.170 126.540 49.780 127.020 ;
        RECT 50.040 126.790 50.300 127.470 ;
        RECT 50.490 126.540 51.080 127.290 ;
        RECT 51.260 126.610 51.430 127.470 ;
        RECT 51.610 126.790 51.860 128.450 ;
      LAYER li1 ;
        RECT 52.430 127.700 52.760 128.270 ;
      LAYER li1 ;
        RECT 52.940 127.520 53.110 129.460 ;
        RECT 52.040 127.350 53.110 127.520 ;
        RECT 52.040 126.610 52.210 127.350 ;
        RECT 53.290 127.170 53.460 129.280 ;
        RECT 53.640 127.260 53.810 129.460 ;
        RECT 53.990 128.780 54.320 129.280 ;
        RECT 53.990 127.310 54.160 128.780 ;
        RECT 54.760 128.500 54.930 129.460 ;
        RECT 55.110 128.850 55.350 129.730 ;
        RECT 55.530 129.680 55.560 129.850 ;
        RECT 55.730 129.680 55.860 129.850 ;
        RECT 55.530 129.030 55.860 129.680 ;
        RECT 57.000 129.850 57.950 129.880 ;
        RECT 57.000 129.680 57.030 129.850 ;
        RECT 57.200 129.680 57.390 129.850 ;
        RECT 57.560 129.680 57.750 129.850 ;
        RECT 57.920 129.680 57.950 129.850 ;
        RECT 56.490 129.020 56.820 129.280 ;
        RECT 56.040 128.850 56.820 129.020 ;
        RECT 57.000 128.850 57.950 129.680 ;
        RECT 58.620 129.770 59.750 129.980 ;
        RECT 59.930 129.850 60.880 129.880 ;
        RECT 58.620 129.020 58.790 129.770 ;
        RECT 59.930 129.680 59.960 129.850 ;
        RECT 60.130 129.680 60.320 129.850 ;
        RECT 60.490 129.680 60.680 129.850 ;
        RECT 60.850 129.680 60.880 129.850 ;
        RECT 58.970 129.200 59.580 129.590 ;
        RECT 58.620 128.850 59.230 129.020 ;
        RECT 55.110 128.680 56.210 128.850 ;
        RECT 56.390 128.500 58.880 128.670 ;
        RECT 54.340 128.150 54.580 128.340 ;
        RECT 54.760 128.330 56.560 128.500 ;
        RECT 56.740 128.150 58.370 128.320 ;
        RECT 58.550 128.260 58.880 128.500 ;
        RECT 54.340 127.980 56.910 128.150 ;
        RECT 58.200 128.050 58.370 128.150 ;
        RECT 59.060 128.050 59.230 128.850 ;
        RECT 54.340 127.670 54.580 127.980 ;
        RECT 55.060 127.490 55.790 127.800 ;
      LAYER li1 ;
        RECT 57.090 127.730 58.020 127.970 ;
      LAYER li1 ;
        RECT 51.260 126.440 52.210 126.610 ;
        RECT 52.390 126.540 52.930 127.170 ;
        RECT 53.110 126.670 53.460 127.170 ;
        RECT 53.990 127.140 56.240 127.310 ;
        RECT 53.990 126.670 54.240 127.140 ;
        RECT 54.780 126.540 55.730 126.960 ;
        RECT 55.910 126.440 56.240 127.140 ;
        RECT 56.720 126.540 57.670 127.550 ;
      LAYER li1 ;
        RECT 57.850 127.180 58.020 127.730 ;
      LAYER li1 ;
        RECT 58.200 127.880 59.230 128.050 ;
        RECT 59.410 128.660 59.580 129.200 ;
        RECT 59.930 128.840 60.880 129.680 ;
        RECT 61.220 129.430 61.470 129.930 ;
        RECT 61.650 129.850 62.600 129.910 ;
        RECT 65.050 129.900 66.500 129.930 ;
        RECT 61.650 129.680 61.680 129.850 ;
        RECT 61.850 129.680 62.040 129.850 ;
        RECT 62.210 129.680 62.400 129.850 ;
        RECT 62.570 129.680 62.600 129.850 ;
        RECT 61.650 129.530 62.600 129.680 ;
        RECT 63.220 129.850 64.160 129.880 ;
        RECT 63.220 129.680 63.240 129.850 ;
        RECT 63.410 129.680 63.600 129.850 ;
        RECT 63.770 129.680 63.960 129.850 ;
        RECT 64.130 129.680 64.160 129.850 ;
        RECT 61.300 129.350 61.470 129.430 ;
        RECT 61.300 129.180 62.480 129.350 ;
        RECT 61.330 128.850 61.660 129.000 ;
        RECT 61.330 128.660 62.130 128.850 ;
        RECT 59.410 128.490 62.130 128.660 ;
        RECT 58.200 127.720 58.710 127.880 ;
        RECT 59.410 127.650 59.580 128.490 ;
        RECT 60.230 128.000 60.560 128.310 ;
        RECT 61.800 128.180 62.130 128.490 ;
        RECT 62.310 128.000 62.480 129.180 ;
        RECT 60.230 127.830 62.480 128.000 ;
        RECT 62.790 128.570 63.040 129.540 ;
        RECT 63.220 128.750 64.160 129.680 ;
        RECT 65.050 129.730 65.300 129.900 ;
        RECT 65.470 129.730 65.660 129.900 ;
        RECT 65.830 129.730 66.100 129.900 ;
        RECT 66.270 129.730 66.500 129.900 ;
        RECT 65.050 128.860 66.500 129.730 ;
        RECT 67.770 129.850 68.360 129.930 ;
        RECT 67.770 129.680 67.800 129.850 ;
        RECT 67.970 129.680 68.160 129.850 ;
        RECT 68.330 129.680 68.360 129.850 ;
        RECT 62.790 128.400 64.160 128.570 ;
        RECT 60.230 127.720 60.560 127.830 ;
        RECT 58.950 127.360 59.580 127.650 ;
      LAYER li1 ;
        RECT 60.810 127.180 61.080 127.210 ;
        RECT 57.850 127.010 61.080 127.180 ;
        RECT 58.210 126.730 61.080 127.010 ;
      LAYER li1 ;
        RECT 61.260 126.540 61.850 127.650 ;
        RECT 62.040 127.150 62.370 127.830 ;
        RECT 62.790 127.650 63.000 128.400 ;
        RECT 63.830 127.900 64.160 128.400 ;
        RECT 62.670 127.150 63.000 127.650 ;
        RECT 63.180 126.540 64.130 127.650 ;
        RECT 65.280 127.420 65.610 128.200 ;
        RECT 65.820 127.870 66.150 128.860 ;
        RECT 67.770 128.350 68.360 129.680 ;
      LAYER li1 ;
        RECT 68.640 128.350 69.030 129.930 ;
      LAYER li1 ;
        RECT 69.620 129.900 72.360 129.920 ;
        RECT 69.620 129.730 69.830 129.900 ;
        RECT 70.000 129.730 70.270 129.900 ;
        RECT 70.440 129.730 70.680 129.900 ;
        RECT 70.850 129.730 71.110 129.900 ;
        RECT 71.280 129.730 71.550 129.900 ;
        RECT 71.720 129.730 71.960 129.900 ;
        RECT 72.130 129.730 72.360 129.900 ;
        RECT 69.620 128.850 72.360 129.730 ;
        RECT 65.280 127.020 66.580 127.420 ;
        RECT 64.970 126.540 66.580 127.020 ;
        RECT 67.770 126.540 68.360 127.500 ;
      LAYER li1 ;
        RECT 68.700 126.670 69.030 128.350 ;
      LAYER li1 ;
        RECT 69.860 127.530 70.190 128.200 ;
        RECT 70.590 127.870 70.920 128.850 ;
        RECT 71.140 127.530 71.470 128.200 ;
        RECT 71.870 127.870 72.200 128.850 ;
        RECT 69.700 126.530 72.430 127.530 ;
      LAYER li1 ;
        RECT 74.510 127.500 74.760 129.910 ;
      LAYER li1 ;
        RECT 74.940 129.850 75.840 129.930 ;
        RECT 74.940 129.680 74.950 129.850 ;
        RECT 75.120 129.680 75.310 129.850 ;
        RECT 75.480 129.680 75.670 129.850 ;
        RECT 74.940 128.450 75.840 129.680 ;
        RECT 76.020 128.270 76.270 129.930 ;
        RECT 76.720 128.620 77.050 129.930 ;
        RECT 77.230 129.850 78.180 129.930 ;
        RECT 77.230 129.680 77.260 129.850 ;
        RECT 77.430 129.680 77.620 129.850 ;
        RECT 77.790 129.680 77.980 129.850 ;
        RECT 78.150 129.680 78.180 129.850 ;
        RECT 77.230 128.800 78.180 129.680 ;
        RECT 78.360 128.620 78.610 129.910 ;
        RECT 78.970 129.900 80.420 129.930 ;
        RECT 78.970 129.730 79.220 129.900 ;
        RECT 79.390 129.730 79.580 129.900 ;
        RECT 79.750 129.730 80.020 129.900 ;
        RECT 80.190 129.730 80.420 129.900 ;
        RECT 78.970 128.860 80.420 129.730 ;
        RECT 80.730 129.850 82.400 129.930 ;
        RECT 80.730 129.680 80.760 129.850 ;
        RECT 80.930 129.680 81.120 129.850 ;
        RECT 81.290 129.680 81.480 129.850 ;
        RECT 81.650 129.680 81.840 129.850 ;
        RECT 82.010 129.680 82.200 129.850 ;
        RECT 82.370 129.680 82.400 129.850 ;
        RECT 76.720 128.450 78.610 128.620 ;
        RECT 78.360 128.370 78.610 128.450 ;
        RECT 74.970 128.100 77.030 128.270 ;
        RECT 74.970 127.900 75.300 128.100 ;
      LAYER li1 ;
        RECT 75.490 127.680 76.680 127.920 ;
      LAYER li1 ;
        RECT 76.860 127.500 77.030 128.100 ;
      LAYER li1 ;
        RECT 78.300 127.680 78.600 128.010 ;
        RECT 74.510 126.670 74.860 127.500 ;
      LAYER li1 ;
        RECT 75.040 126.540 76.650 127.500 ;
        RECT 76.830 126.670 77.080 127.500 ;
        RECT 77.260 126.540 78.570 127.500 ;
        RECT 79.200 127.420 79.530 128.200 ;
        RECT 79.740 127.870 80.070 128.860 ;
        RECT 80.730 128.470 82.400 129.680 ;
      LAYER li1 ;
        RECT 80.770 127.700 81.070 128.290 ;
        RECT 81.250 127.950 82.440 128.290 ;
        RECT 82.620 127.950 82.950 129.430 ;
        RECT 83.130 127.770 83.400 129.930 ;
      LAYER li1 ;
        RECT 84.500 129.900 87.240 129.920 ;
        RECT 84.500 129.730 84.710 129.900 ;
        RECT 84.880 129.730 85.150 129.900 ;
        RECT 85.320 129.730 85.560 129.900 ;
        RECT 85.730 129.730 85.990 129.900 ;
        RECT 86.160 129.730 86.430 129.900 ;
        RECT 86.600 129.730 86.840 129.900 ;
        RECT 87.010 129.730 87.240 129.900 ;
        RECT 84.500 128.850 87.240 129.730 ;
        RECT 88.340 129.900 91.080 129.920 ;
        RECT 88.340 129.730 88.550 129.900 ;
        RECT 88.720 129.730 88.990 129.900 ;
        RECT 89.160 129.730 89.400 129.900 ;
        RECT 89.570 129.730 89.830 129.900 ;
        RECT 90.000 129.730 90.270 129.900 ;
        RECT 90.440 129.730 90.680 129.900 ;
        RECT 90.850 129.730 91.080 129.900 ;
        RECT 88.340 128.850 91.080 129.730 ;
        RECT 92.180 129.900 94.920 129.920 ;
        RECT 92.180 129.730 92.390 129.900 ;
        RECT 92.560 129.730 92.830 129.900 ;
        RECT 93.000 129.730 93.240 129.900 ;
        RECT 93.410 129.730 93.670 129.900 ;
        RECT 93.840 129.730 94.110 129.900 ;
        RECT 94.280 129.730 94.520 129.900 ;
        RECT 94.690 129.730 94.920 129.900 ;
        RECT 92.180 128.850 94.920 129.730 ;
        RECT 95.770 129.900 97.220 129.930 ;
        RECT 95.770 129.730 96.020 129.900 ;
        RECT 96.190 129.730 96.380 129.900 ;
        RECT 96.550 129.730 96.820 129.900 ;
        RECT 96.990 129.730 97.220 129.900 ;
        RECT 95.770 128.860 97.220 129.730 ;
      LAYER li1 ;
        RECT 81.570 127.600 83.400 127.770 ;
      LAYER li1 ;
        RECT 79.200 127.020 80.500 127.420 ;
        RECT 78.890 126.540 80.500 127.020 ;
        RECT 80.730 126.540 81.320 127.500 ;
      LAYER li1 ;
        RECT 81.570 126.670 81.820 127.600 ;
      LAYER li1 ;
        RECT 82.000 126.540 82.950 127.420 ;
      LAYER li1 ;
        RECT 83.130 126.670 83.400 127.600 ;
      LAYER li1 ;
        RECT 84.740 127.530 85.070 128.200 ;
        RECT 85.470 127.870 85.800 128.850 ;
        RECT 86.020 127.530 86.350 128.200 ;
        RECT 86.750 127.870 87.080 128.850 ;
        RECT 88.580 127.530 88.910 128.200 ;
        RECT 89.310 127.870 89.640 128.850 ;
        RECT 89.860 127.530 90.190 128.200 ;
        RECT 90.590 127.870 90.920 128.850 ;
        RECT 92.420 127.530 92.750 128.200 ;
        RECT 93.150 127.870 93.480 128.850 ;
        RECT 93.700 127.530 94.030 128.200 ;
        RECT 94.430 127.870 94.760 128.850 ;
        RECT 84.580 126.530 87.310 127.530 ;
        RECT 88.420 126.530 91.150 127.530 ;
        RECT 92.260 126.530 94.990 127.530 ;
        RECT 96.000 127.420 96.330 128.200 ;
        RECT 96.540 127.870 96.870 128.860 ;
        RECT 96.000 127.020 97.300 127.420 ;
        RECT 95.690 126.540 97.300 127.020 ;
      LAYER li1 ;
        RECT 97.570 126.670 97.820 129.930 ;
      LAYER li1 ;
        RECT 98.000 129.850 100.690 129.930 ;
        RECT 98.170 129.680 98.360 129.850 ;
        RECT 98.530 129.680 98.720 129.850 ;
        RECT 98.890 129.680 99.080 129.850 ;
        RECT 99.250 129.680 99.440 129.850 ;
        RECT 99.610 129.680 99.800 129.850 ;
        RECT 99.970 129.680 100.160 129.850 ;
        RECT 100.330 129.680 100.520 129.850 ;
        RECT 98.000 128.820 100.690 129.680 ;
        RECT 100.870 128.640 101.120 129.930 ;
        RECT 98.030 128.470 101.120 128.640 ;
        RECT 98.030 127.770 98.360 128.470 ;
        RECT 100.870 128.350 101.120 128.470 ;
        RECT 101.300 129.850 102.610 129.910 ;
        RECT 101.300 129.680 101.330 129.850 ;
        RECT 101.500 129.680 101.690 129.850 ;
        RECT 101.860 129.680 102.050 129.850 ;
        RECT 102.220 129.680 102.410 129.850 ;
        RECT 102.580 129.680 102.610 129.850 ;
        RECT 101.300 128.370 102.610 129.680 ;
        RECT 103.220 129.900 105.960 129.920 ;
        RECT 103.220 129.730 103.430 129.900 ;
        RECT 103.600 129.730 103.870 129.900 ;
        RECT 104.040 129.730 104.280 129.900 ;
        RECT 104.450 129.730 104.710 129.900 ;
        RECT 104.880 129.730 105.150 129.900 ;
        RECT 105.320 129.730 105.560 129.900 ;
        RECT 105.730 129.730 105.960 129.900 ;
        RECT 103.220 128.850 105.960 129.730 ;
        RECT 107.060 129.900 109.800 129.920 ;
        RECT 107.060 129.730 107.270 129.900 ;
        RECT 107.440 129.730 107.710 129.900 ;
        RECT 107.880 129.730 108.120 129.900 ;
        RECT 108.290 129.730 108.550 129.900 ;
        RECT 108.720 129.730 108.990 129.900 ;
        RECT 109.160 129.730 109.400 129.900 ;
        RECT 109.570 129.730 109.800 129.900 ;
        RECT 107.060 128.850 109.800 129.730 ;
      LAYER li1 ;
        RECT 99.030 128.230 99.200 128.290 ;
        RECT 98.860 127.950 99.590 128.230 ;
      LAYER li1 ;
        RECT 98.030 127.600 99.240 127.770 ;
        RECT 98.000 126.540 98.890 127.420 ;
        RECT 99.070 127.390 99.240 127.600 ;
      LAYER li1 ;
        RECT 99.420 127.740 99.590 127.950 ;
        RECT 99.770 127.920 100.200 128.290 ;
        RECT 100.400 127.750 100.690 128.290 ;
        RECT 100.930 127.750 101.640 128.080 ;
        RECT 99.420 127.570 100.220 127.740 ;
        RECT 101.990 127.570 102.320 128.190 ;
        RECT 100.050 127.400 102.320 127.570 ;
      LAYER li1 ;
        RECT 103.460 127.530 103.790 128.200 ;
        RECT 104.190 127.870 104.520 128.850 ;
        RECT 104.740 127.530 105.070 128.200 ;
        RECT 105.470 127.870 105.800 128.850 ;
        RECT 107.300 127.530 107.630 128.200 ;
        RECT 108.030 127.870 108.360 128.850 ;
        RECT 108.580 127.530 108.910 128.200 ;
        RECT 109.310 127.870 109.640 128.850 ;
      LAYER li1 ;
        RECT 111.000 128.350 111.430 129.930 ;
      LAYER li1 ;
        RECT 111.610 129.850 112.170 129.930 ;
        RECT 111.610 129.680 111.620 129.850 ;
        RECT 111.790 129.680 111.980 129.850 ;
        RECT 112.150 129.680 112.170 129.850 ;
        RECT 111.610 128.350 112.170 129.680 ;
        RECT 113.780 129.900 116.520 129.920 ;
        RECT 113.780 129.730 113.990 129.900 ;
        RECT 114.160 129.730 114.430 129.900 ;
        RECT 114.600 129.730 114.840 129.900 ;
        RECT 115.010 129.730 115.270 129.900 ;
        RECT 115.440 129.730 115.710 129.900 ;
        RECT 115.880 129.730 116.120 129.900 ;
        RECT 116.290 129.730 116.520 129.900 ;
        RECT 99.070 127.220 99.870 127.390 ;
      LAYER li1 ;
        RECT 100.480 127.380 101.150 127.400 ;
      LAYER li1 ;
        RECT 99.700 127.050 100.300 127.220 ;
        RECT 99.190 126.610 99.520 127.040 ;
        RECT 99.970 126.790 100.300 127.050 ;
        RECT 100.790 126.610 101.120 127.200 ;
        RECT 99.190 126.440 101.120 126.610 ;
        RECT 101.330 126.540 102.630 127.220 ;
        RECT 103.300 126.530 106.030 127.530 ;
        RECT 107.140 126.530 109.870 127.530 ;
      LAYER li1 ;
        RECT 111.000 126.670 111.250 128.350 ;
      LAYER li1 ;
        RECT 111.560 127.460 111.890 127.920 ;
      LAYER li1 ;
        RECT 112.350 127.640 112.680 129.430 ;
      LAYER li1 ;
        RECT 112.860 127.460 113.110 129.180 ;
        RECT 113.780 128.850 116.520 129.730 ;
        RECT 114.020 127.530 114.350 128.200 ;
        RECT 114.750 127.870 115.080 128.850 ;
        RECT 115.300 127.530 115.630 128.200 ;
        RECT 116.030 127.870 116.360 128.850 ;
      LAYER li1 ;
        RECT 118.680 128.350 119.110 129.930 ;
      LAYER li1 ;
        RECT 119.290 129.850 119.850 129.930 ;
        RECT 119.290 129.680 119.300 129.850 ;
        RECT 119.470 129.680 119.660 129.850 ;
        RECT 119.830 129.680 119.850 129.850 ;
        RECT 119.290 128.350 119.850 129.680 ;
        RECT 121.460 129.900 124.200 129.920 ;
        RECT 121.460 129.730 121.670 129.900 ;
        RECT 121.840 129.730 122.110 129.900 ;
        RECT 122.280 129.730 122.520 129.900 ;
        RECT 122.690 129.730 122.950 129.900 ;
        RECT 123.120 129.730 123.390 129.900 ;
        RECT 123.560 129.730 123.800 129.900 ;
        RECT 123.970 129.730 124.200 129.900 ;
        RECT 111.560 127.290 113.110 127.460 ;
        RECT 111.430 126.540 112.680 127.110 ;
        RECT 112.860 126.670 113.110 127.290 ;
        RECT 113.860 126.530 116.590 127.530 ;
      LAYER li1 ;
        RECT 118.680 126.670 118.930 128.350 ;
      LAYER li1 ;
        RECT 119.240 127.460 119.570 127.920 ;
      LAYER li1 ;
        RECT 120.030 127.640 120.360 129.430 ;
      LAYER li1 ;
        RECT 120.540 127.460 120.790 129.180 ;
        RECT 121.460 128.850 124.200 129.730 ;
        RECT 125.300 129.900 128.040 129.920 ;
        RECT 125.300 129.730 125.510 129.900 ;
        RECT 125.680 129.730 125.950 129.900 ;
        RECT 126.120 129.730 126.360 129.900 ;
        RECT 126.530 129.730 126.790 129.900 ;
        RECT 126.960 129.730 127.230 129.900 ;
        RECT 127.400 129.730 127.640 129.900 ;
        RECT 127.810 129.730 128.040 129.900 ;
        RECT 125.300 128.850 128.040 129.730 ;
        RECT 129.140 129.900 131.880 129.920 ;
        RECT 129.140 129.730 129.350 129.900 ;
        RECT 129.520 129.730 129.790 129.900 ;
        RECT 129.960 129.730 130.200 129.900 ;
        RECT 130.370 129.730 130.630 129.900 ;
        RECT 130.800 129.730 131.070 129.900 ;
        RECT 131.240 129.730 131.480 129.900 ;
        RECT 131.650 129.730 131.880 129.900 ;
        RECT 129.140 128.850 131.880 129.730 ;
        RECT 132.980 129.900 135.720 129.920 ;
        RECT 132.980 129.730 133.190 129.900 ;
        RECT 133.360 129.730 133.630 129.900 ;
        RECT 133.800 129.730 134.040 129.900 ;
        RECT 134.210 129.730 134.470 129.900 ;
        RECT 134.640 129.730 134.910 129.900 ;
        RECT 135.080 129.730 135.320 129.900 ;
        RECT 135.490 129.730 135.720 129.900 ;
        RECT 132.980 128.850 135.720 129.730 ;
        RECT 136.820 129.900 139.560 129.920 ;
        RECT 136.820 129.730 137.030 129.900 ;
        RECT 137.200 129.730 137.470 129.900 ;
        RECT 137.640 129.730 137.880 129.900 ;
        RECT 138.050 129.730 138.310 129.900 ;
        RECT 138.480 129.730 138.750 129.900 ;
        RECT 138.920 129.730 139.160 129.900 ;
        RECT 139.330 129.730 139.560 129.900 ;
        RECT 136.820 128.850 139.560 129.730 ;
        RECT 140.410 129.900 141.860 129.930 ;
        RECT 140.410 129.730 140.660 129.900 ;
        RECT 140.830 129.730 141.020 129.900 ;
        RECT 141.190 129.730 141.460 129.900 ;
        RECT 141.630 129.730 141.860 129.900 ;
        RECT 140.410 128.860 141.860 129.730 ;
        RECT 121.700 127.530 122.030 128.200 ;
        RECT 122.430 127.870 122.760 128.850 ;
        RECT 122.980 127.530 123.310 128.200 ;
        RECT 123.710 127.870 124.040 128.850 ;
        RECT 125.540 127.530 125.870 128.200 ;
        RECT 126.270 127.870 126.600 128.850 ;
        RECT 126.820 127.530 127.150 128.200 ;
        RECT 127.550 127.870 127.880 128.850 ;
        RECT 129.380 127.530 129.710 128.200 ;
        RECT 130.110 127.870 130.440 128.850 ;
        RECT 130.660 127.530 130.990 128.200 ;
        RECT 131.390 127.870 131.720 128.850 ;
        RECT 133.220 127.530 133.550 128.200 ;
        RECT 133.950 127.870 134.280 128.850 ;
        RECT 134.500 127.530 134.830 128.200 ;
        RECT 135.230 127.870 135.560 128.850 ;
        RECT 137.060 127.530 137.390 128.200 ;
        RECT 137.790 127.870 138.120 128.850 ;
        RECT 138.340 127.530 138.670 128.200 ;
        RECT 139.070 127.870 139.400 128.850 ;
        RECT 119.240 127.290 120.790 127.460 ;
        RECT 119.110 126.540 120.360 127.110 ;
        RECT 120.540 126.670 120.790 127.290 ;
        RECT 121.540 126.530 124.270 127.530 ;
        RECT 125.380 126.530 128.110 127.530 ;
        RECT 129.220 126.530 131.950 127.530 ;
        RECT 133.060 126.530 135.790 127.530 ;
        RECT 136.900 126.530 139.630 127.530 ;
        RECT 140.640 127.420 140.970 128.200 ;
        RECT 141.180 127.870 141.510 128.860 ;
        RECT 140.640 127.020 141.940 127.420 ;
        RECT 140.330 126.540 141.940 127.020 ;
        RECT 5.760 126.080 5.920 126.260 ;
        RECT 6.090 126.080 6.400 126.260 ;
        RECT 6.570 126.080 6.880 126.260 ;
        RECT 7.050 126.080 7.360 126.260 ;
        RECT 7.530 126.080 7.840 126.260 ;
        RECT 8.010 126.080 8.320 126.260 ;
        RECT 8.490 126.080 8.800 126.260 ;
        RECT 8.970 126.080 9.280 126.260 ;
        RECT 9.450 126.080 9.760 126.260 ;
        RECT 9.930 126.080 10.240 126.260 ;
        RECT 10.410 126.080 10.720 126.260 ;
        RECT 10.890 126.080 11.200 126.260 ;
        RECT 11.370 126.080 11.680 126.260 ;
        RECT 11.850 126.080 12.160 126.260 ;
        RECT 12.330 126.080 12.640 126.260 ;
        RECT 12.810 126.080 13.120 126.260 ;
        RECT 13.290 126.080 13.600 126.260 ;
        RECT 13.770 126.080 14.080 126.260 ;
        RECT 14.250 126.080 14.560 126.260 ;
        RECT 14.730 126.080 15.040 126.260 ;
        RECT 15.210 126.080 15.520 126.260 ;
        RECT 15.690 126.080 16.000 126.260 ;
        RECT 16.170 126.080 16.480 126.260 ;
        RECT 16.650 126.080 16.960 126.260 ;
        RECT 17.130 126.080 17.440 126.260 ;
        RECT 17.610 126.080 17.920 126.260 ;
        RECT 18.090 126.080 18.400 126.260 ;
        RECT 18.570 126.080 18.880 126.260 ;
        RECT 19.050 126.080 19.360 126.260 ;
        RECT 19.530 126.080 19.840 126.260 ;
        RECT 20.010 126.080 20.320 126.260 ;
        RECT 20.490 126.080 20.800 126.260 ;
        RECT 20.970 126.080 21.280 126.260 ;
        RECT 21.450 126.080 21.760 126.260 ;
        RECT 21.930 126.080 22.240 126.260 ;
        RECT 22.410 126.080 22.720 126.260 ;
        RECT 22.890 126.080 23.200 126.260 ;
        RECT 23.370 126.080 23.680 126.260 ;
        RECT 23.850 126.080 24.160 126.260 ;
        RECT 24.330 126.080 24.640 126.260 ;
        RECT 24.810 126.080 25.120 126.260 ;
        RECT 25.290 126.080 25.600 126.260 ;
        RECT 25.770 126.080 26.080 126.260 ;
        RECT 26.250 126.080 26.560 126.260 ;
        RECT 26.730 126.080 27.040 126.260 ;
        RECT 27.210 126.080 27.520 126.260 ;
        RECT 27.690 126.080 28.000 126.260 ;
        RECT 28.170 126.080 28.480 126.260 ;
        RECT 28.650 126.080 28.960 126.260 ;
        RECT 29.130 126.080 29.440 126.260 ;
        RECT 29.610 126.080 29.920 126.260 ;
        RECT 30.090 126.080 30.400 126.260 ;
        RECT 30.570 126.080 30.880 126.260 ;
        RECT 31.050 126.080 31.360 126.260 ;
        RECT 31.530 126.080 31.840 126.260 ;
        RECT 32.010 126.080 32.320 126.260 ;
        RECT 32.490 126.080 32.800 126.260 ;
        RECT 32.970 126.080 33.280 126.260 ;
        RECT 33.450 126.080 33.760 126.260 ;
        RECT 33.930 126.080 34.080 126.260 ;
        RECT 34.560 126.080 34.720 126.260 ;
        RECT 34.890 126.080 35.200 126.260 ;
        RECT 35.370 126.080 35.680 126.260 ;
        RECT 35.850 126.080 36.160 126.260 ;
        RECT 36.330 126.080 36.640 126.260 ;
        RECT 36.810 126.080 37.120 126.260 ;
        RECT 37.290 126.080 37.600 126.260 ;
        RECT 37.770 126.080 38.080 126.260 ;
        RECT 38.250 126.080 38.560 126.260 ;
        RECT 38.730 126.080 39.040 126.260 ;
        RECT 39.210 126.080 39.520 126.260 ;
        RECT 39.690 126.080 40.000 126.260 ;
        RECT 40.170 126.080 40.480 126.260 ;
        RECT 40.650 126.080 40.960 126.260 ;
        RECT 41.130 126.080 41.440 126.260 ;
        RECT 41.610 126.080 41.920 126.260 ;
        RECT 42.090 126.080 42.400 126.260 ;
        RECT 42.570 126.080 42.880 126.260 ;
        RECT 43.050 126.080 43.360 126.260 ;
        RECT 43.530 126.080 43.680 126.260 ;
        RECT 44.160 126.080 44.320 126.260 ;
        RECT 44.490 126.080 44.800 126.260 ;
        RECT 44.970 126.080 45.280 126.260 ;
        RECT 45.450 126.080 45.760 126.260 ;
        RECT 45.930 126.080 46.240 126.260 ;
        RECT 46.410 126.080 46.720 126.260 ;
        RECT 46.890 126.080 47.200 126.260 ;
        RECT 47.370 126.080 47.680 126.260 ;
        RECT 47.850 126.080 48.160 126.260 ;
        RECT 48.330 126.080 48.640 126.260 ;
        RECT 48.810 126.080 49.120 126.260 ;
        RECT 49.290 126.080 49.600 126.260 ;
        RECT 49.770 126.080 50.080 126.260 ;
        RECT 50.250 126.080 50.560 126.260 ;
        RECT 50.730 126.080 51.040 126.260 ;
        RECT 51.210 126.080 51.520 126.260 ;
        RECT 51.690 126.080 52.000 126.260 ;
        RECT 52.170 126.080 52.480 126.260 ;
        RECT 52.650 126.080 52.960 126.260 ;
        RECT 53.130 126.080 53.440 126.260 ;
        RECT 53.610 126.080 53.920 126.260 ;
        RECT 54.090 126.080 54.400 126.260 ;
        RECT 54.570 126.080 54.880 126.260 ;
        RECT 55.050 126.080 55.360 126.260 ;
        RECT 55.530 126.080 55.840 126.260 ;
        RECT 56.010 126.080 56.320 126.260 ;
        RECT 56.490 126.080 56.800 126.260 ;
        RECT 56.970 126.080 57.280 126.260 ;
        RECT 57.450 126.080 57.760 126.260 ;
        RECT 57.930 126.080 58.240 126.260 ;
        RECT 58.410 126.080 58.720 126.260 ;
        RECT 58.890 126.080 59.200 126.260 ;
        RECT 59.370 126.080 59.680 126.260 ;
        RECT 59.850 126.080 60.160 126.260 ;
        RECT 60.330 126.080 60.640 126.260 ;
        RECT 60.810 126.080 61.120 126.260 ;
        RECT 61.290 126.080 61.600 126.260 ;
        RECT 61.770 126.080 62.080 126.260 ;
        RECT 62.250 126.080 62.560 126.260 ;
        RECT 62.730 126.080 63.040 126.260 ;
        RECT 63.210 126.080 63.520 126.260 ;
        RECT 63.690 126.080 64.000 126.260 ;
        RECT 64.170 126.080 64.480 126.260 ;
        RECT 64.650 126.080 64.960 126.260 ;
        RECT 65.130 126.080 65.440 126.260 ;
        RECT 65.610 126.080 65.920 126.260 ;
        RECT 66.090 126.080 66.400 126.260 ;
        RECT 66.570 126.080 66.880 126.260 ;
        RECT 67.050 126.080 67.360 126.260 ;
        RECT 67.530 126.080 67.840 126.260 ;
        RECT 68.010 126.080 68.320 126.260 ;
        RECT 68.490 126.080 68.800 126.260 ;
        RECT 68.970 126.080 69.280 126.260 ;
        RECT 69.450 126.080 69.760 126.260 ;
        RECT 69.930 126.080 70.240 126.260 ;
        RECT 70.410 126.080 70.720 126.260 ;
        RECT 70.890 126.080 71.200 126.260 ;
        RECT 71.370 126.080 71.680 126.260 ;
        RECT 71.850 126.080 72.160 126.260 ;
        RECT 72.330 126.080 72.640 126.260 ;
        RECT 72.810 126.080 73.120 126.260 ;
        RECT 73.290 126.080 73.600 126.260 ;
        RECT 73.770 126.080 73.920 126.260 ;
        RECT 74.400 126.080 74.560 126.260 ;
        RECT 74.730 126.080 75.040 126.260 ;
        RECT 75.210 126.080 75.520 126.260 ;
        RECT 75.690 126.080 76.000 126.260 ;
        RECT 76.170 126.080 76.480 126.260 ;
        RECT 76.650 126.080 76.960 126.260 ;
        RECT 77.130 126.080 77.440 126.260 ;
        RECT 77.610 126.080 77.920 126.260 ;
        RECT 78.090 126.080 78.400 126.260 ;
        RECT 78.570 126.080 78.880 126.260 ;
        RECT 79.050 126.080 79.360 126.260 ;
        RECT 79.530 126.080 79.840 126.260 ;
        RECT 80.010 126.080 80.320 126.260 ;
        RECT 80.490 126.080 80.800 126.260 ;
        RECT 80.970 126.080 81.280 126.260 ;
        RECT 81.450 126.080 81.760 126.260 ;
        RECT 81.930 126.080 82.240 126.260 ;
        RECT 82.410 126.080 82.720 126.260 ;
        RECT 82.890 126.080 83.200 126.260 ;
        RECT 83.370 126.080 83.680 126.260 ;
        RECT 83.850 126.080 84.160 126.260 ;
        RECT 84.330 126.080 84.640 126.260 ;
        RECT 84.810 126.080 85.120 126.260 ;
        RECT 85.290 126.080 85.600 126.260 ;
        RECT 85.770 126.080 86.080 126.260 ;
        RECT 86.250 126.080 86.560 126.260 ;
        RECT 86.730 126.080 87.040 126.260 ;
        RECT 87.210 126.080 87.520 126.260 ;
        RECT 87.690 126.080 88.000 126.260 ;
        RECT 88.170 126.080 88.480 126.260 ;
        RECT 88.650 126.080 88.960 126.260 ;
        RECT 89.130 126.080 89.440 126.260 ;
        RECT 89.610 126.080 89.920 126.260 ;
        RECT 90.090 126.080 90.400 126.260 ;
        RECT 90.570 126.080 90.880 126.260 ;
        RECT 91.050 126.080 91.360 126.260 ;
        RECT 91.530 126.080 91.840 126.260 ;
        RECT 92.010 126.080 92.320 126.260 ;
        RECT 92.490 126.080 92.800 126.260 ;
        RECT 92.970 126.080 93.280 126.260 ;
        RECT 93.450 126.080 93.760 126.260 ;
        RECT 93.930 126.080 94.240 126.260 ;
        RECT 94.410 126.080 94.720 126.260 ;
        RECT 94.890 126.080 95.200 126.260 ;
        RECT 95.370 126.080 95.680 126.260 ;
        RECT 95.850 126.080 96.160 126.260 ;
        RECT 96.330 126.080 96.640 126.260 ;
        RECT 96.810 126.080 97.120 126.260 ;
        RECT 97.290 126.080 97.600 126.260 ;
        RECT 97.770 126.080 98.080 126.260 ;
        RECT 98.250 126.080 98.560 126.260 ;
        RECT 98.730 126.080 99.040 126.260 ;
        RECT 99.210 126.080 99.520 126.260 ;
        RECT 99.690 126.080 100.000 126.260 ;
        RECT 100.170 126.080 100.480 126.260 ;
        RECT 100.650 126.080 100.960 126.260 ;
        RECT 101.130 126.080 101.440 126.260 ;
        RECT 101.610 126.080 101.920 126.260 ;
        RECT 102.090 126.080 102.400 126.260 ;
        RECT 102.570 126.080 102.880 126.260 ;
        RECT 103.050 126.080 103.360 126.260 ;
        RECT 103.530 126.080 103.840 126.260 ;
        RECT 104.010 126.080 104.320 126.260 ;
        RECT 104.490 126.080 104.800 126.260 ;
        RECT 104.970 126.080 105.280 126.260 ;
        RECT 105.450 126.080 105.760 126.260 ;
        RECT 105.930 126.080 106.240 126.260 ;
        RECT 106.410 126.080 106.720 126.260 ;
        RECT 106.890 126.080 107.200 126.260 ;
        RECT 107.370 126.080 107.680 126.260 ;
        RECT 107.850 126.080 108.160 126.260 ;
        RECT 108.330 126.080 108.640 126.260 ;
        RECT 108.810 126.080 109.120 126.260 ;
        RECT 109.290 126.080 109.600 126.260 ;
        RECT 109.770 126.080 110.080 126.260 ;
        RECT 110.250 126.080 110.400 126.260 ;
        RECT 110.880 126.080 111.040 126.260 ;
        RECT 111.210 126.080 111.520 126.260 ;
        RECT 111.690 126.080 112.000 126.260 ;
        RECT 112.170 126.080 112.480 126.260 ;
        RECT 112.650 126.080 112.960 126.260 ;
        RECT 113.130 126.080 113.440 126.260 ;
        RECT 113.610 126.080 113.920 126.260 ;
        RECT 114.090 126.080 114.400 126.260 ;
        RECT 114.570 126.080 114.880 126.260 ;
        RECT 115.050 126.080 115.360 126.260 ;
        RECT 115.530 126.080 115.840 126.260 ;
        RECT 116.010 126.080 116.320 126.260 ;
        RECT 116.490 126.080 116.800 126.260 ;
        RECT 116.970 126.080 117.280 126.260 ;
        RECT 117.450 126.080 117.760 126.260 ;
        RECT 117.930 126.080 118.080 126.260 ;
        RECT 118.560 126.080 118.720 126.260 ;
        RECT 118.890 126.080 119.200 126.260 ;
        RECT 119.370 126.080 119.680 126.260 ;
        RECT 119.850 126.080 120.160 126.260 ;
        RECT 120.330 126.080 120.640 126.260 ;
        RECT 120.810 126.080 121.120 126.260 ;
        RECT 121.290 126.080 121.600 126.260 ;
        RECT 121.770 126.080 122.080 126.260 ;
        RECT 122.250 126.080 122.560 126.260 ;
        RECT 122.730 126.080 123.040 126.260 ;
        RECT 123.210 126.080 123.520 126.260 ;
        RECT 123.690 126.080 124.000 126.260 ;
        RECT 124.170 126.080 124.480 126.260 ;
        RECT 124.650 126.080 124.960 126.260 ;
        RECT 125.130 126.080 125.440 126.260 ;
        RECT 125.610 126.080 125.920 126.260 ;
        RECT 126.090 126.080 126.400 126.260 ;
        RECT 126.570 126.080 126.880 126.260 ;
        RECT 127.050 126.080 127.360 126.260 ;
        RECT 127.530 126.080 127.840 126.260 ;
        RECT 128.010 126.080 128.320 126.260 ;
        RECT 128.490 126.080 128.800 126.260 ;
        RECT 128.970 126.080 129.280 126.260 ;
        RECT 129.450 126.080 129.760 126.260 ;
        RECT 129.930 126.080 130.240 126.260 ;
        RECT 130.410 126.080 130.720 126.260 ;
        RECT 130.890 126.080 131.200 126.260 ;
        RECT 131.370 126.080 131.680 126.260 ;
        RECT 131.850 126.080 132.160 126.260 ;
        RECT 132.330 126.080 132.640 126.260 ;
        RECT 132.810 126.080 133.120 126.260 ;
        RECT 133.290 126.080 133.600 126.260 ;
        RECT 133.770 126.080 134.080 126.260 ;
        RECT 134.250 126.080 134.560 126.260 ;
        RECT 134.730 126.080 135.040 126.260 ;
        RECT 135.210 126.080 135.520 126.260 ;
        RECT 135.690 126.080 136.000 126.260 ;
        RECT 136.170 126.080 136.480 126.260 ;
        RECT 136.650 126.080 136.960 126.260 ;
        RECT 137.130 126.080 137.440 126.260 ;
        RECT 137.610 126.080 137.920 126.260 ;
        RECT 138.090 126.080 138.400 126.260 ;
        RECT 138.570 126.080 138.880 126.260 ;
        RECT 139.050 126.080 139.360 126.260 ;
        RECT 139.530 126.080 139.840 126.260 ;
        RECT 140.010 126.080 140.320 126.260 ;
        RECT 140.490 126.080 140.800 126.260 ;
        RECT 140.970 126.080 141.280 126.260 ;
        RECT 141.450 126.080 141.760 126.260 ;
        RECT 141.930 126.080 142.080 126.260 ;
        RECT 5.930 125.770 7.540 125.800 ;
        RECT 5.930 125.600 5.980 125.770 ;
        RECT 6.150 125.600 6.420 125.770 ;
        RECT 6.590 125.600 6.860 125.770 ;
        RECT 7.030 125.600 7.270 125.770 ;
        RECT 7.440 125.600 7.540 125.770 ;
        RECT 8.720 125.770 9.670 125.800 ;
        RECT 5.930 125.320 7.540 125.600 ;
        RECT 6.240 124.920 7.540 125.320 ;
        RECT 6.240 124.140 6.570 124.920 ;
        RECT 6.780 123.480 7.110 124.470 ;
        RECT 8.270 123.810 8.540 125.670 ;
        RECT 8.720 125.600 8.750 125.770 ;
        RECT 8.920 125.600 9.110 125.770 ;
        RECT 9.280 125.600 9.470 125.770 ;
        RECT 9.640 125.600 9.670 125.770 ;
        RECT 10.360 125.770 10.950 125.800 ;
        RECT 8.720 125.170 9.670 125.600 ;
        RECT 9.850 125.170 10.180 125.670 ;
        RECT 9.400 123.810 9.730 124.310 ;
        RECT 8.270 123.640 9.730 123.810 ;
        RECT 6.010 122.610 7.460 123.480 ;
        RECT 8.270 122.710 8.600 123.640 ;
        RECT 6.010 122.440 6.260 122.610 ;
        RECT 6.430 122.440 6.620 122.610 ;
        RECT 6.790 122.440 7.060 122.610 ;
        RECT 7.230 122.440 7.460 122.610 ;
        RECT 8.790 122.660 9.380 123.440 ;
        RECT 8.790 122.490 8.820 122.660 ;
        RECT 8.990 122.490 9.180 122.660 ;
        RECT 9.350 122.490 9.380 122.660 ;
        RECT 8.790 122.460 9.380 122.490 ;
        RECT 9.560 122.530 9.730 123.640 ;
        RECT 9.910 124.250 10.180 125.170 ;
        RECT 10.360 125.600 10.390 125.770 ;
        RECT 10.560 125.600 10.750 125.770 ;
        RECT 10.920 125.600 10.950 125.770 ;
        RECT 15.320 125.770 16.270 125.800 ;
        RECT 10.360 124.920 10.950 125.600 ;
      LAYER li1 ;
        RECT 11.230 125.540 14.170 125.710 ;
        RECT 11.230 125.330 11.400 125.540 ;
        RECT 11.190 125.160 11.400 125.330 ;
        RECT 11.230 124.550 11.400 125.160 ;
      LAYER li1 ;
        RECT 9.910 124.020 10.440 124.250 ;
        RECT 9.910 122.710 10.160 124.020 ;
      LAYER li1 ;
        RECT 10.860 123.680 11.400 124.550 ;
        RECT 11.580 124.060 11.910 125.360 ;
      LAYER li1 ;
        RECT 12.090 124.840 12.360 125.340 ;
        RECT 12.810 125.090 13.140 125.340 ;
        RECT 12.810 124.920 13.820 125.090 ;
        RECT 12.090 123.850 12.260 124.840 ;
        RECT 13.140 124.250 13.470 124.740 ;
        RECT 12.040 123.680 12.260 123.850 ;
        RECT 12.440 124.020 13.470 124.250 ;
        RECT 13.650 124.690 13.820 124.920 ;
      LAYER li1 ;
        RECT 14.000 125.040 14.170 125.540 ;
      LAYER li1 ;
        RECT 15.320 125.600 15.350 125.770 ;
        RECT 15.520 125.600 15.710 125.770 ;
        RECT 15.880 125.600 16.070 125.770 ;
        RECT 16.240 125.600 16.270 125.770 ;
        RECT 15.320 125.220 16.270 125.600 ;
      LAYER li1 ;
        RECT 16.450 125.730 19.110 125.900 ;
        RECT 16.450 125.040 16.620 125.730 ;
        RECT 14.000 124.870 16.620 125.040 ;
      LAYER li1 ;
        RECT 13.650 124.520 16.270 124.690 ;
        RECT 12.040 123.500 12.210 123.680 ;
        RECT 12.440 123.500 12.610 124.020 ;
        RECT 13.650 123.840 13.820 124.520 ;
      LAYER li1 ;
        RECT 16.450 124.340 16.620 124.870 ;
      LAYER li1 ;
        RECT 10.400 123.330 12.210 123.500 ;
        RECT 10.400 122.710 10.650 123.330 ;
        RECT 10.830 122.980 11.860 123.150 ;
        RECT 10.830 122.530 11.000 122.980 ;
        RECT 6.010 122.410 7.460 122.440 ;
        RECT 9.560 122.360 11.000 122.530 ;
        RECT 11.180 122.660 11.510 122.800 ;
        RECT 11.180 122.490 11.210 122.660 ;
        RECT 11.380 122.490 11.510 122.660 ;
        RECT 11.180 122.460 11.510 122.490 ;
        RECT 11.690 122.530 11.860 122.980 ;
        RECT 12.040 122.710 12.210 123.330 ;
        RECT 12.390 123.170 12.610 123.500 ;
        RECT 12.790 123.670 13.820 123.840 ;
        RECT 14.000 123.990 14.330 124.340 ;
      LAYER li1 ;
        RECT 14.770 124.170 16.620 124.340 ;
      LAYER li1 ;
        RECT 16.800 124.840 17.130 125.550 ;
        RECT 17.590 125.380 18.760 125.550 ;
        RECT 17.590 124.840 17.920 125.380 ;
        RECT 16.800 123.990 17.060 124.840 ;
        RECT 18.130 124.580 18.410 125.080 ;
        RECT 14.000 123.820 17.060 123.990 ;
        RECT 12.790 122.970 12.960 123.670 ;
        RECT 13.650 123.640 13.820 123.670 ;
        RECT 13.140 123.290 13.470 123.490 ;
        RECT 13.650 123.470 15.420 123.640 ;
        RECT 13.140 123.170 14.910 123.290 ;
        RECT 13.260 123.120 14.910 123.170 ;
        RECT 12.740 122.710 13.070 122.970 ;
        RECT 13.260 122.530 13.430 123.120 ;
        RECT 11.690 122.360 13.430 122.530 ;
        RECT 13.610 122.660 14.560 122.940 ;
        RECT 13.610 122.490 13.640 122.660 ;
        RECT 13.810 122.490 14.000 122.660 ;
        RECT 14.170 122.490 14.360 122.660 ;
        RECT 14.530 122.490 14.560 122.660 ;
        RECT 13.610 122.460 14.560 122.490 ;
        RECT 14.740 122.530 14.910 123.120 ;
        RECT 15.090 122.710 15.420 123.470 ;
        RECT 16.730 123.240 17.060 123.820 ;
        RECT 17.240 124.410 18.410 124.580 ;
        RECT 17.240 123.060 17.410 124.410 ;
        RECT 17.790 123.730 18.120 124.230 ;
        RECT 18.590 123.980 18.760 125.380 ;
      LAYER li1 ;
        RECT 18.940 125.070 19.110 125.730 ;
      LAYER li1 ;
        RECT 19.290 125.770 20.240 125.800 ;
        RECT 19.290 125.600 19.320 125.770 ;
        RECT 19.490 125.600 19.680 125.770 ;
        RECT 19.850 125.600 20.040 125.770 ;
        RECT 20.210 125.600 20.240 125.770 ;
        RECT 21.900 125.770 22.850 125.800 ;
        RECT 19.290 125.250 20.240 125.600 ;
        RECT 20.780 125.170 21.110 125.670 ;
        RECT 21.900 125.600 21.930 125.770 ;
        RECT 22.100 125.600 22.290 125.770 ;
        RECT 22.460 125.600 22.650 125.770 ;
        RECT 22.820 125.600 22.850 125.770 ;
      LAYER li1 ;
        RECT 18.940 124.900 19.950 125.070 ;
      LAYER li1 ;
        RECT 18.970 124.330 19.300 124.720 ;
      LAYER li1 ;
        RECT 19.620 124.510 19.950 124.900 ;
      LAYER li1 ;
        RECT 20.780 124.330 21.010 125.170 ;
        RECT 21.390 124.670 21.720 125.170 ;
        RECT 21.900 124.670 22.850 125.600 ;
        RECT 23.690 125.770 25.300 125.800 ;
        RECT 23.690 125.600 23.740 125.770 ;
        RECT 23.910 125.600 24.180 125.770 ;
        RECT 24.350 125.600 24.620 125.770 ;
        RECT 24.790 125.600 25.030 125.770 ;
        RECT 25.200 125.600 25.300 125.770 ;
        RECT 26.960 125.770 27.910 125.800 ;
        RECT 18.970 124.160 21.010 124.330 ;
        RECT 18.300 123.810 20.660 123.980 ;
        RECT 18.300 123.490 18.470 123.810 ;
        RECT 20.840 123.630 21.010 124.160 ;
        RECT 15.600 122.890 17.410 123.060 ;
        RECT 17.590 123.320 18.470 123.490 ;
        RECT 15.600 122.530 15.770 122.890 ;
        RECT 14.740 122.360 15.770 122.530 ;
        RECT 15.950 122.660 16.900 122.710 ;
        RECT 15.950 122.490 15.980 122.660 ;
        RECT 16.150 122.490 16.340 122.660 ;
        RECT 16.510 122.490 16.700 122.660 ;
        RECT 16.870 122.490 16.900 122.660 ;
        RECT 15.950 122.410 16.900 122.490 ;
        RECT 17.590 122.410 17.840 123.320 ;
        RECT 18.650 122.660 19.600 123.490 ;
        RECT 20.000 123.460 21.010 123.630 ;
        RECT 21.510 124.490 21.720 124.670 ;
        RECT 21.510 124.160 22.880 124.490 ;
        RECT 20.000 122.990 20.250 123.460 ;
        RECT 20.430 122.660 21.330 123.280 ;
        RECT 21.510 123.160 21.760 124.160 ;
        RECT 18.650 122.490 18.680 122.660 ;
        RECT 18.850 122.490 19.040 122.660 ;
        RECT 19.210 122.490 19.400 122.660 ;
        RECT 19.570 122.490 19.600 122.660 ;
        RECT 20.600 122.490 20.790 122.660 ;
        RECT 20.960 122.490 21.150 122.660 ;
        RECT 21.320 122.490 21.330 122.660 ;
        RECT 18.650 122.460 19.600 122.490 ;
        RECT 20.430 122.460 21.330 122.490 ;
        RECT 21.940 122.660 22.880 123.970 ;
        RECT 21.940 122.490 21.960 122.660 ;
        RECT 22.130 122.490 22.320 122.660 ;
        RECT 22.490 122.490 22.680 122.660 ;
        RECT 22.850 122.490 22.880 122.660 ;
        RECT 21.940 122.430 22.880 122.490 ;
      LAYER li1 ;
        RECT 23.060 122.430 23.400 125.500 ;
      LAYER li1 ;
        RECT 23.690 125.320 25.300 125.600 ;
        RECT 24.000 124.920 25.300 125.320 ;
        RECT 24.000 124.140 24.330 124.920 ;
        RECT 24.540 123.480 24.870 124.470 ;
        RECT 26.510 123.810 26.780 125.670 ;
        RECT 26.960 125.600 26.990 125.770 ;
        RECT 27.160 125.600 27.350 125.770 ;
        RECT 27.520 125.600 27.710 125.770 ;
        RECT 27.880 125.600 27.910 125.770 ;
        RECT 28.600 125.770 29.190 125.800 ;
        RECT 26.960 125.170 27.910 125.600 ;
        RECT 28.090 125.170 28.420 125.670 ;
        RECT 27.640 123.810 27.970 124.310 ;
        RECT 26.510 123.640 27.970 123.810 ;
        RECT 23.770 122.610 25.220 123.480 ;
        RECT 26.510 122.710 26.840 123.640 ;
        RECT 23.770 122.440 24.020 122.610 ;
        RECT 24.190 122.440 24.380 122.610 ;
        RECT 24.550 122.440 24.820 122.610 ;
        RECT 24.990 122.440 25.220 122.610 ;
        RECT 27.030 122.660 27.620 123.440 ;
        RECT 27.030 122.490 27.060 122.660 ;
        RECT 27.230 122.490 27.420 122.660 ;
        RECT 27.590 122.490 27.620 122.660 ;
        RECT 27.030 122.460 27.620 122.490 ;
        RECT 27.800 122.530 27.970 123.640 ;
        RECT 28.150 124.250 28.420 125.170 ;
        RECT 28.600 125.600 28.630 125.770 ;
        RECT 28.800 125.600 28.990 125.770 ;
        RECT 29.160 125.600 29.190 125.770 ;
        RECT 33.560 125.770 34.510 125.800 ;
        RECT 28.600 124.920 29.190 125.600 ;
      LAYER li1 ;
        RECT 29.470 125.540 32.410 125.710 ;
        RECT 29.470 124.550 29.640 125.540 ;
      LAYER li1 ;
        RECT 28.150 124.020 28.680 124.250 ;
        RECT 28.150 122.710 28.400 124.020 ;
      LAYER li1 ;
        RECT 29.100 123.680 29.640 124.550 ;
        RECT 29.820 124.060 30.150 125.360 ;
      LAYER li1 ;
        RECT 30.330 124.840 30.600 125.340 ;
        RECT 31.050 125.090 31.380 125.340 ;
        RECT 31.050 124.920 32.060 125.090 ;
        RECT 30.330 123.850 30.500 124.840 ;
        RECT 31.380 124.250 31.710 124.740 ;
        RECT 30.280 123.680 30.500 123.850 ;
        RECT 30.680 124.020 31.710 124.250 ;
        RECT 31.890 124.690 32.060 124.920 ;
      LAYER li1 ;
        RECT 32.240 125.040 32.410 125.540 ;
      LAYER li1 ;
        RECT 33.560 125.600 33.590 125.770 ;
        RECT 33.760 125.600 33.950 125.770 ;
        RECT 34.120 125.600 34.310 125.770 ;
        RECT 34.480 125.600 34.510 125.770 ;
        RECT 33.560 125.220 34.510 125.600 ;
      LAYER li1 ;
        RECT 34.690 125.730 37.350 125.900 ;
        RECT 34.690 125.040 34.860 125.730 ;
        RECT 32.240 124.870 34.860 125.040 ;
      LAYER li1 ;
        RECT 31.890 124.520 34.510 124.690 ;
        RECT 30.280 123.500 30.450 123.680 ;
        RECT 30.680 123.500 30.850 124.020 ;
        RECT 31.890 123.840 32.060 124.520 ;
      LAYER li1 ;
        RECT 34.690 124.340 34.860 124.870 ;
      LAYER li1 ;
        RECT 28.640 123.330 30.450 123.500 ;
        RECT 28.640 122.710 28.890 123.330 ;
        RECT 29.070 122.980 30.100 123.150 ;
        RECT 29.070 122.530 29.240 122.980 ;
        RECT 23.770 122.410 25.220 122.440 ;
        RECT 27.800 122.360 29.240 122.530 ;
        RECT 29.420 122.660 29.750 122.800 ;
        RECT 29.420 122.490 29.450 122.660 ;
        RECT 29.620 122.490 29.750 122.660 ;
        RECT 29.420 122.460 29.750 122.490 ;
        RECT 29.930 122.530 30.100 122.980 ;
        RECT 30.280 122.710 30.450 123.330 ;
        RECT 30.630 123.170 30.850 123.500 ;
        RECT 31.030 123.670 32.060 123.840 ;
        RECT 32.240 123.990 32.570 124.340 ;
      LAYER li1 ;
        RECT 33.010 124.170 34.860 124.340 ;
      LAYER li1 ;
        RECT 35.040 124.840 35.370 125.550 ;
        RECT 35.830 125.380 37.000 125.550 ;
        RECT 35.830 124.840 36.160 125.380 ;
        RECT 35.040 123.990 35.300 124.840 ;
        RECT 36.370 124.580 36.650 125.080 ;
        RECT 32.240 123.820 35.300 123.990 ;
        RECT 31.030 122.970 31.200 123.670 ;
        RECT 31.890 123.640 32.060 123.670 ;
        RECT 31.380 123.290 31.710 123.490 ;
        RECT 31.890 123.470 33.660 123.640 ;
        RECT 31.380 123.170 33.150 123.290 ;
        RECT 31.500 123.120 33.150 123.170 ;
        RECT 30.980 122.710 31.310 122.970 ;
        RECT 31.500 122.530 31.670 123.120 ;
        RECT 29.930 122.360 31.670 122.530 ;
        RECT 31.850 122.660 32.800 122.940 ;
        RECT 31.850 122.490 31.880 122.660 ;
        RECT 32.050 122.490 32.240 122.660 ;
        RECT 32.410 122.490 32.600 122.660 ;
        RECT 32.770 122.490 32.800 122.660 ;
        RECT 31.850 122.460 32.800 122.490 ;
        RECT 32.980 122.530 33.150 123.120 ;
        RECT 33.330 122.710 33.660 123.470 ;
        RECT 34.970 123.240 35.300 123.820 ;
        RECT 35.480 124.410 36.650 124.580 ;
        RECT 35.480 123.060 35.650 124.410 ;
        RECT 36.030 123.730 36.360 124.230 ;
        RECT 36.830 123.980 37.000 125.380 ;
      LAYER li1 ;
        RECT 37.180 125.070 37.350 125.730 ;
      LAYER li1 ;
        RECT 37.530 125.770 38.480 125.800 ;
        RECT 37.530 125.600 37.560 125.770 ;
        RECT 37.730 125.600 37.920 125.770 ;
        RECT 38.090 125.600 38.280 125.770 ;
        RECT 38.450 125.600 38.480 125.770 ;
        RECT 40.140 125.770 41.090 125.800 ;
        RECT 37.530 125.250 38.480 125.600 ;
        RECT 39.020 125.170 39.350 125.670 ;
        RECT 40.140 125.600 40.170 125.770 ;
        RECT 40.340 125.600 40.530 125.770 ;
        RECT 40.700 125.600 40.890 125.770 ;
        RECT 41.060 125.600 41.090 125.770 ;
      LAYER li1 ;
        RECT 37.180 124.960 38.190 125.070 ;
        RECT 37.180 124.900 38.240 124.960 ;
        RECT 37.860 124.790 38.240 124.900 ;
      LAYER li1 ;
        RECT 37.210 124.330 37.540 124.720 ;
      LAYER li1 ;
        RECT 37.860 124.510 38.190 124.790 ;
      LAYER li1 ;
        RECT 39.020 124.330 39.250 125.170 ;
        RECT 39.630 124.670 39.960 125.170 ;
        RECT 40.140 124.670 41.090 125.600 ;
        RECT 41.930 125.770 43.540 125.800 ;
        RECT 41.930 125.600 41.980 125.770 ;
        RECT 42.150 125.600 42.420 125.770 ;
        RECT 42.590 125.600 42.860 125.770 ;
        RECT 43.030 125.600 43.270 125.770 ;
        RECT 43.440 125.600 43.540 125.770 ;
        RECT 44.710 125.770 46.420 125.800 ;
        RECT 37.210 124.160 39.250 124.330 ;
        RECT 36.540 123.810 38.900 123.980 ;
        RECT 36.540 123.490 36.710 123.810 ;
        RECT 39.080 123.630 39.250 124.160 ;
        RECT 33.840 122.890 35.650 123.060 ;
        RECT 35.830 123.320 36.710 123.490 ;
        RECT 33.840 122.530 34.010 122.890 ;
        RECT 32.980 122.360 34.010 122.530 ;
        RECT 34.190 122.660 35.140 122.710 ;
        RECT 34.190 122.490 34.220 122.660 ;
        RECT 34.390 122.490 34.580 122.660 ;
        RECT 34.750 122.490 34.940 122.660 ;
        RECT 35.110 122.490 35.140 122.660 ;
        RECT 34.190 122.410 35.140 122.490 ;
        RECT 35.830 122.410 36.080 123.320 ;
        RECT 36.890 122.660 37.840 123.490 ;
        RECT 38.240 123.460 39.250 123.630 ;
        RECT 39.750 124.490 39.960 124.670 ;
        RECT 39.750 124.160 41.120 124.490 ;
        RECT 38.240 122.990 38.490 123.460 ;
        RECT 38.670 122.660 39.570 123.280 ;
        RECT 39.750 123.160 40.000 124.160 ;
        RECT 36.890 122.490 36.920 122.660 ;
        RECT 37.090 122.490 37.280 122.660 ;
        RECT 37.450 122.490 37.640 122.660 ;
        RECT 37.810 122.490 37.840 122.660 ;
        RECT 38.840 122.490 39.030 122.660 ;
        RECT 39.200 122.490 39.390 122.660 ;
        RECT 39.560 122.490 39.570 122.660 ;
        RECT 36.890 122.460 37.840 122.490 ;
        RECT 38.670 122.460 39.570 122.490 ;
        RECT 40.180 122.660 41.120 123.970 ;
        RECT 40.180 122.490 40.200 122.660 ;
        RECT 40.370 122.490 40.560 122.660 ;
        RECT 40.730 122.490 40.920 122.660 ;
        RECT 41.090 122.490 41.120 122.660 ;
        RECT 40.180 122.430 41.120 122.490 ;
      LAYER li1 ;
        RECT 41.300 122.430 41.640 125.500 ;
      LAYER li1 ;
        RECT 41.930 125.320 43.540 125.600 ;
        RECT 42.240 124.920 43.540 125.320 ;
        RECT 42.240 124.140 42.570 124.920 ;
        RECT 42.780 123.480 43.110 124.470 ;
        RECT 42.010 122.610 43.460 123.480 ;
        RECT 42.010 122.440 42.260 122.610 ;
        RECT 42.430 122.440 42.620 122.610 ;
        RECT 42.790 122.440 43.060 122.610 ;
        RECT 43.230 122.440 43.460 122.610 ;
        RECT 42.010 122.410 43.460 122.440 ;
      LAYER li1 ;
        RECT 44.270 122.410 44.540 125.670 ;
      LAYER li1 ;
        RECT 44.710 125.600 44.760 125.770 ;
        RECT 44.930 125.600 45.120 125.770 ;
        RECT 45.290 125.600 45.480 125.770 ;
        RECT 45.650 125.600 45.840 125.770 ;
        RECT 46.010 125.600 46.200 125.770 ;
        RECT 46.370 125.600 46.420 125.770 ;
        RECT 47.980 125.770 49.290 125.800 ;
        RECT 44.710 124.920 46.420 125.600 ;
        RECT 46.850 125.540 47.800 125.710 ;
        RECT 46.850 124.740 47.020 125.540 ;
        RECT 44.750 124.570 47.020 124.740 ;
      LAYER li1 ;
        RECT 47.200 124.590 47.370 125.360 ;
      LAYER li1 ;
        RECT 47.550 124.840 47.800 125.540 ;
        RECT 47.980 125.600 48.010 125.770 ;
        RECT 48.180 125.600 48.370 125.770 ;
        RECT 48.540 125.600 48.730 125.770 ;
        RECT 48.900 125.600 49.090 125.770 ;
        RECT 49.260 125.600 49.290 125.770 ;
        RECT 47.980 124.840 49.290 125.600 ;
        RECT 50.020 125.780 52.750 125.810 ;
        RECT 50.020 125.610 50.190 125.780 ;
        RECT 50.360 125.610 50.630 125.780 ;
        RECT 50.800 125.610 51.040 125.780 ;
        RECT 51.210 125.610 51.470 125.780 ;
        RECT 51.640 125.610 51.910 125.780 ;
        RECT 52.080 125.610 52.320 125.780 ;
        RECT 52.490 125.610 52.750 125.780 ;
        RECT 50.020 124.810 52.750 125.610 ;
        RECT 53.860 125.780 56.590 125.810 ;
        RECT 53.860 125.610 54.030 125.780 ;
        RECT 54.200 125.610 54.470 125.780 ;
        RECT 54.640 125.610 54.880 125.780 ;
        RECT 55.050 125.610 55.310 125.780 ;
        RECT 55.480 125.610 55.750 125.780 ;
        RECT 55.920 125.610 56.160 125.780 ;
        RECT 56.330 125.610 56.590 125.780 ;
        RECT 58.630 125.770 59.880 125.800 ;
        RECT 61.060 125.780 63.790 125.810 ;
        RECT 53.860 124.810 56.590 125.610 ;
        RECT 44.750 124.410 45.080 124.570 ;
        RECT 44.720 122.660 45.620 123.990 ;
        RECT 44.720 122.490 44.730 122.660 ;
        RECT 44.900 122.490 45.090 122.660 ;
        RECT 45.260 122.490 45.450 122.660 ;
        RECT 45.800 122.530 45.970 123.990 ;
      LAYER li1 ;
        RECT 46.150 122.910 46.480 124.390 ;
      LAYER li1 ;
        RECT 46.660 122.710 46.990 124.570 ;
      LAYER li1 ;
        RECT 47.190 124.420 47.370 124.590 ;
        RECT 47.650 124.420 48.810 124.660 ;
      LAYER li1 ;
        RECT 47.440 124.070 49.330 124.240 ;
        RECT 50.180 124.140 50.510 124.810 ;
        RECT 47.440 122.530 47.690 124.070 ;
        RECT 44.720 122.410 45.620 122.490 ;
        RECT 45.800 122.360 47.690 122.530 ;
        RECT 47.870 122.660 48.820 123.890 ;
        RECT 47.870 122.490 47.900 122.660 ;
        RECT 48.070 122.490 48.260 122.660 ;
        RECT 48.430 122.490 48.620 122.660 ;
        RECT 48.790 122.490 48.820 122.660 ;
        RECT 47.870 122.410 48.820 122.490 ;
        RECT 49.000 122.430 49.330 124.070 ;
        RECT 50.910 123.490 51.240 124.470 ;
        RECT 51.460 124.140 51.790 124.810 ;
        RECT 52.190 123.490 52.520 124.470 ;
        RECT 54.020 124.140 54.350 124.810 ;
        RECT 54.750 123.490 55.080 124.470 ;
        RECT 55.300 124.140 55.630 124.810 ;
        RECT 56.030 123.490 56.360 124.470 ;
      LAYER li1 ;
        RECT 58.200 123.990 58.450 125.670 ;
      LAYER li1 ;
        RECT 58.800 125.600 58.990 125.770 ;
        RECT 59.160 125.600 59.350 125.770 ;
        RECT 59.520 125.600 59.710 125.770 ;
        RECT 58.630 125.230 59.880 125.600 ;
        RECT 60.060 125.050 60.310 125.670 ;
        RECT 58.760 124.880 60.310 125.050 ;
        RECT 58.760 124.420 59.090 124.880 ;
        RECT 49.940 122.610 52.680 123.490 ;
        RECT 49.940 122.440 50.150 122.610 ;
        RECT 50.320 122.440 50.590 122.610 ;
        RECT 50.760 122.440 51.000 122.610 ;
        RECT 51.170 122.440 51.430 122.610 ;
        RECT 51.600 122.440 51.870 122.610 ;
        RECT 52.040 122.440 52.280 122.610 ;
        RECT 52.450 122.440 52.680 122.610 ;
        RECT 49.940 122.420 52.680 122.440 ;
        RECT 53.780 122.610 56.520 123.490 ;
        RECT 53.780 122.440 53.990 122.610 ;
        RECT 54.160 122.440 54.430 122.610 ;
        RECT 54.600 122.440 54.840 122.610 ;
        RECT 55.010 122.440 55.270 122.610 ;
        RECT 55.440 122.440 55.710 122.610 ;
        RECT 55.880 122.440 56.120 122.610 ;
        RECT 56.290 122.440 56.520 122.610 ;
        RECT 53.780 122.420 56.520 122.440 ;
      LAYER li1 ;
        RECT 58.200 122.410 58.630 123.990 ;
      LAYER li1 ;
        RECT 58.810 122.660 59.370 123.990 ;
      LAYER li1 ;
        RECT 59.550 122.910 59.880 124.700 ;
      LAYER li1 ;
        RECT 60.060 123.160 60.310 124.880 ;
        RECT 61.060 125.610 61.230 125.780 ;
        RECT 61.400 125.610 61.670 125.780 ;
        RECT 61.840 125.610 62.080 125.780 ;
        RECT 62.250 125.610 62.510 125.780 ;
        RECT 62.680 125.610 62.950 125.780 ;
        RECT 63.120 125.610 63.360 125.780 ;
        RECT 63.530 125.610 63.790 125.780 ;
        RECT 61.060 124.810 63.790 125.610 ;
        RECT 64.900 125.780 67.630 125.810 ;
        RECT 64.900 125.610 65.070 125.780 ;
        RECT 65.240 125.610 65.510 125.780 ;
        RECT 65.680 125.610 65.920 125.780 ;
        RECT 66.090 125.610 66.350 125.780 ;
        RECT 66.520 125.610 66.790 125.780 ;
        RECT 66.960 125.610 67.200 125.780 ;
        RECT 67.370 125.610 67.630 125.780 ;
        RECT 64.900 124.810 67.630 125.610 ;
        RECT 68.740 125.780 71.470 125.810 ;
        RECT 68.740 125.610 68.910 125.780 ;
        RECT 69.080 125.610 69.350 125.780 ;
        RECT 69.520 125.610 69.760 125.780 ;
        RECT 69.930 125.610 70.190 125.780 ;
        RECT 70.360 125.610 70.630 125.780 ;
        RECT 70.800 125.610 71.040 125.780 ;
        RECT 71.210 125.610 71.470 125.780 ;
        RECT 68.740 124.810 71.470 125.610 ;
        RECT 72.170 125.770 73.780 125.800 ;
        RECT 72.170 125.600 72.220 125.770 ;
        RECT 72.390 125.600 72.660 125.770 ;
        RECT 72.830 125.600 73.100 125.770 ;
        RECT 73.270 125.600 73.510 125.770 ;
        RECT 73.680 125.600 73.780 125.770 ;
        RECT 72.170 125.320 73.780 125.600 ;
        RECT 72.480 124.920 73.780 125.320 ;
        RECT 74.970 125.770 75.560 125.800 ;
        RECT 74.970 125.600 75.000 125.770 ;
        RECT 75.170 125.600 75.360 125.770 ;
        RECT 75.530 125.600 75.560 125.770 ;
        RECT 76.240 125.770 77.190 125.800 ;
        RECT 61.220 124.140 61.550 124.810 ;
        RECT 61.950 123.490 62.280 124.470 ;
        RECT 62.500 124.140 62.830 124.810 ;
        RECT 63.230 123.490 63.560 124.470 ;
        RECT 65.060 124.140 65.390 124.810 ;
        RECT 65.790 123.490 66.120 124.470 ;
        RECT 66.340 124.140 66.670 124.810 ;
        RECT 67.070 123.490 67.400 124.470 ;
        RECT 68.900 124.140 69.230 124.810 ;
        RECT 69.630 123.490 69.960 124.470 ;
        RECT 70.180 124.140 70.510 124.810 ;
        RECT 70.910 123.490 71.240 124.470 ;
        RECT 72.480 124.140 72.810 124.920 ;
        RECT 74.970 124.840 75.560 125.600 ;
      LAYER li1 ;
        RECT 75.810 124.740 76.060 125.670 ;
      LAYER li1 ;
        RECT 76.240 125.600 76.270 125.770 ;
        RECT 76.440 125.600 76.630 125.770 ;
        RECT 76.800 125.600 76.990 125.770 ;
        RECT 77.160 125.600 77.190 125.770 ;
        RECT 78.820 125.780 81.550 125.810 ;
        RECT 76.240 124.920 77.190 125.600 ;
      LAYER li1 ;
        RECT 77.370 124.740 77.640 125.670 ;
      LAYER li1 ;
        RECT 78.820 125.610 78.990 125.780 ;
        RECT 79.160 125.610 79.430 125.780 ;
        RECT 79.600 125.610 79.840 125.780 ;
        RECT 80.010 125.610 80.270 125.780 ;
        RECT 80.440 125.610 80.710 125.780 ;
        RECT 80.880 125.610 81.120 125.780 ;
        RECT 81.290 125.610 81.550 125.780 ;
        RECT 78.820 124.810 81.550 125.610 ;
        RECT 82.660 125.780 85.390 125.810 ;
        RECT 82.660 125.610 82.830 125.780 ;
        RECT 83.000 125.610 83.270 125.780 ;
        RECT 83.440 125.610 83.680 125.780 ;
        RECT 83.850 125.610 84.110 125.780 ;
        RECT 84.280 125.610 84.550 125.780 ;
        RECT 84.720 125.610 84.960 125.780 ;
        RECT 85.130 125.610 85.390 125.780 ;
        RECT 82.660 124.810 85.390 125.610 ;
        RECT 86.500 125.780 89.230 125.810 ;
        RECT 86.500 125.610 86.670 125.780 ;
        RECT 86.840 125.610 87.110 125.780 ;
        RECT 87.280 125.610 87.520 125.780 ;
        RECT 87.690 125.610 87.950 125.780 ;
        RECT 88.120 125.610 88.390 125.780 ;
        RECT 88.560 125.610 88.800 125.780 ;
        RECT 88.970 125.610 89.230 125.780 ;
        RECT 86.500 124.810 89.230 125.610 ;
        RECT 90.810 125.770 91.400 125.800 ;
        RECT 90.810 125.600 90.840 125.770 ;
        RECT 91.010 125.600 91.200 125.770 ;
        RECT 91.370 125.600 91.400 125.770 ;
        RECT 92.330 125.770 93.940 125.800 ;
        RECT 94.640 125.770 95.530 125.800 ;
        RECT 90.810 124.840 91.400 125.600 ;
        RECT 58.810 122.490 58.820 122.660 ;
        RECT 58.990 122.490 59.180 122.660 ;
        RECT 59.350 122.490 59.370 122.660 ;
        RECT 58.810 122.410 59.370 122.490 ;
        RECT 60.980 122.610 63.720 123.490 ;
        RECT 60.980 122.440 61.190 122.610 ;
        RECT 61.360 122.440 61.630 122.610 ;
        RECT 61.800 122.440 62.040 122.610 ;
        RECT 62.210 122.440 62.470 122.610 ;
        RECT 62.640 122.440 62.910 122.610 ;
        RECT 63.080 122.440 63.320 122.610 ;
        RECT 63.490 122.440 63.720 122.610 ;
        RECT 60.980 122.420 63.720 122.440 ;
        RECT 64.820 122.610 67.560 123.490 ;
        RECT 64.820 122.440 65.030 122.610 ;
        RECT 65.200 122.440 65.470 122.610 ;
        RECT 65.640 122.440 65.880 122.610 ;
        RECT 66.050 122.440 66.310 122.610 ;
        RECT 66.480 122.440 66.750 122.610 ;
        RECT 66.920 122.440 67.160 122.610 ;
        RECT 67.330 122.440 67.560 122.610 ;
        RECT 64.820 122.420 67.560 122.440 ;
        RECT 68.660 122.610 71.400 123.490 ;
        RECT 73.020 123.480 73.350 124.470 ;
      LAYER li1 ;
        RECT 75.010 124.050 75.310 124.640 ;
        RECT 75.810 124.570 77.640 124.740 ;
        RECT 75.490 124.050 76.680 124.390 ;
      LAYER li1 ;
        RECT 68.660 122.440 68.870 122.610 ;
        RECT 69.040 122.440 69.310 122.610 ;
        RECT 69.480 122.440 69.720 122.610 ;
        RECT 69.890 122.440 70.150 122.610 ;
        RECT 70.320 122.440 70.590 122.610 ;
        RECT 70.760 122.440 71.000 122.610 ;
        RECT 71.170 122.440 71.400 122.610 ;
        RECT 68.660 122.420 71.400 122.440 ;
        RECT 72.250 122.610 73.700 123.480 ;
        RECT 72.250 122.440 72.500 122.610 ;
        RECT 72.670 122.440 72.860 122.610 ;
        RECT 73.030 122.440 73.300 122.610 ;
        RECT 73.470 122.440 73.700 122.610 ;
        RECT 72.250 122.410 73.700 122.440 ;
        RECT 74.970 122.660 76.640 123.870 ;
      LAYER li1 ;
        RECT 76.860 122.910 77.190 124.390 ;
      LAYER li1 ;
        RECT 74.970 122.490 75.000 122.660 ;
        RECT 75.170 122.490 75.360 122.660 ;
        RECT 75.530 122.490 75.720 122.660 ;
        RECT 75.890 122.490 76.080 122.660 ;
        RECT 76.250 122.490 76.440 122.660 ;
        RECT 76.610 122.490 76.640 122.660 ;
        RECT 74.970 122.410 76.640 122.490 ;
      LAYER li1 ;
        RECT 77.370 122.410 77.640 124.570 ;
      LAYER li1 ;
        RECT 78.980 124.140 79.310 124.810 ;
        RECT 79.710 123.490 80.040 124.470 ;
        RECT 80.260 124.140 80.590 124.810 ;
        RECT 80.990 123.490 81.320 124.470 ;
        RECT 82.820 124.140 83.150 124.810 ;
        RECT 83.550 123.490 83.880 124.470 ;
        RECT 84.100 124.140 84.430 124.810 ;
        RECT 84.830 123.490 85.160 124.470 ;
        RECT 86.660 124.140 86.990 124.810 ;
        RECT 87.390 123.490 87.720 124.470 ;
        RECT 87.940 124.140 88.270 124.810 ;
        RECT 88.670 123.490 89.000 124.470 ;
      LAYER li1 ;
        RECT 90.850 124.230 91.560 124.620 ;
        RECT 91.740 123.990 92.070 125.670 ;
      LAYER li1 ;
        RECT 92.330 125.600 92.380 125.770 ;
        RECT 92.550 125.600 92.820 125.770 ;
        RECT 92.990 125.600 93.260 125.770 ;
        RECT 93.430 125.600 93.670 125.770 ;
        RECT 93.840 125.600 93.940 125.770 ;
        RECT 92.330 125.320 93.940 125.600 ;
        RECT 92.640 124.920 93.940 125.320 ;
        RECT 92.640 124.140 92.970 124.920 ;
        RECT 78.740 122.610 81.480 123.490 ;
        RECT 78.740 122.440 78.950 122.610 ;
        RECT 79.120 122.440 79.390 122.610 ;
        RECT 79.560 122.440 79.800 122.610 ;
        RECT 79.970 122.440 80.230 122.610 ;
        RECT 80.400 122.440 80.670 122.610 ;
        RECT 80.840 122.440 81.080 122.610 ;
        RECT 81.250 122.440 81.480 122.610 ;
        RECT 78.740 122.420 81.480 122.440 ;
        RECT 82.580 122.610 85.320 123.490 ;
        RECT 82.580 122.440 82.790 122.610 ;
        RECT 82.960 122.440 83.230 122.610 ;
        RECT 83.400 122.440 83.640 122.610 ;
        RECT 83.810 122.440 84.070 122.610 ;
        RECT 84.240 122.440 84.510 122.610 ;
        RECT 84.680 122.440 84.920 122.610 ;
        RECT 85.090 122.440 85.320 122.610 ;
        RECT 82.580 122.420 85.320 122.440 ;
        RECT 86.420 122.610 89.160 123.490 ;
        RECT 86.420 122.440 86.630 122.610 ;
        RECT 86.800 122.440 87.070 122.610 ;
        RECT 87.240 122.440 87.480 122.610 ;
        RECT 87.650 122.440 87.910 122.610 ;
        RECT 88.080 122.440 88.350 122.610 ;
        RECT 88.520 122.440 88.760 122.610 ;
        RECT 88.930 122.440 89.160 122.610 ;
        RECT 86.420 122.420 89.160 122.440 ;
        RECT 90.810 122.660 91.400 123.990 ;
        RECT 90.810 122.490 90.840 122.660 ;
        RECT 91.010 122.490 91.200 122.660 ;
        RECT 91.370 122.490 91.400 122.660 ;
        RECT 90.810 122.410 91.400 122.490 ;
      LAYER li1 ;
        RECT 91.680 122.410 92.070 123.990 ;
      LAYER li1 ;
        RECT 93.180 123.480 93.510 124.470 ;
        RECT 92.410 122.610 93.860 123.480 ;
        RECT 92.410 122.440 92.660 122.610 ;
        RECT 92.830 122.440 93.020 122.610 ;
        RECT 93.190 122.440 93.460 122.610 ;
        RECT 93.630 122.440 93.860 122.610 ;
        RECT 92.410 122.410 93.860 122.440 ;
      LAYER li1 ;
        RECT 94.210 122.410 94.460 125.670 ;
      LAYER li1 ;
        RECT 94.810 125.600 95.000 125.770 ;
        RECT 95.170 125.600 95.360 125.770 ;
        RECT 95.830 125.730 97.760 125.900 ;
        RECT 94.640 124.920 95.530 125.600 ;
        RECT 95.830 125.300 96.160 125.730 ;
        RECT 96.610 125.290 96.940 125.550 ;
        RECT 96.340 125.120 96.940 125.290 ;
        RECT 97.430 125.140 97.760 125.730 ;
        RECT 97.970 125.770 99.270 125.800 ;
        RECT 97.970 125.600 98.000 125.770 ;
        RECT 98.170 125.600 98.360 125.770 ;
        RECT 98.530 125.600 98.720 125.770 ;
        RECT 98.890 125.600 99.080 125.770 ;
        RECT 99.250 125.600 99.270 125.770 ;
        RECT 97.970 125.120 99.270 125.600 ;
        RECT 99.530 125.770 101.140 125.800 ;
        RECT 99.530 125.600 99.580 125.770 ;
        RECT 99.750 125.600 100.020 125.770 ;
        RECT 100.190 125.600 100.460 125.770 ;
        RECT 100.630 125.600 100.870 125.770 ;
        RECT 101.040 125.600 101.140 125.770 ;
        RECT 99.530 125.320 101.140 125.600 ;
        RECT 95.710 124.950 96.510 125.120 ;
        RECT 95.710 124.740 95.880 124.950 ;
      LAYER li1 ;
        RECT 97.120 124.940 97.790 124.960 ;
        RECT 96.690 124.770 98.960 124.940 ;
      LAYER li1 ;
        RECT 94.670 124.570 95.880 124.740 ;
      LAYER li1 ;
        RECT 96.060 124.600 96.860 124.770 ;
      LAYER li1 ;
        RECT 94.670 123.870 95.000 124.570 ;
      LAYER li1 ;
        RECT 96.060 124.390 96.230 124.600 ;
        RECT 95.500 124.110 96.230 124.390 ;
        RECT 95.670 124.050 95.840 124.110 ;
        RECT 96.410 124.050 96.840 124.420 ;
        RECT 97.040 124.050 97.330 124.590 ;
        RECT 97.570 124.260 98.280 124.590 ;
        RECT 98.630 124.150 98.960 124.770 ;
      LAYER li1 ;
        RECT 99.840 124.920 101.140 125.320 ;
        RECT 101.440 125.730 103.250 125.900 ;
        RECT 99.840 124.140 100.170 124.920 ;
        RECT 101.440 124.810 101.770 125.730 ;
      LAYER li1 ;
        RECT 102.020 124.810 102.550 125.550 ;
      LAYER li1 ;
        RECT 97.510 123.870 97.760 123.990 ;
        RECT 94.670 123.700 97.760 123.870 ;
        RECT 94.640 122.660 97.330 123.520 ;
        RECT 94.810 122.490 95.000 122.660 ;
        RECT 95.170 122.490 95.360 122.660 ;
        RECT 95.530 122.490 95.720 122.660 ;
        RECT 95.890 122.490 96.080 122.660 ;
        RECT 96.250 122.490 96.440 122.660 ;
        RECT 96.610 122.490 96.800 122.660 ;
        RECT 96.970 122.490 97.160 122.660 ;
        RECT 94.640 122.410 97.330 122.490 ;
        RECT 97.510 122.410 97.760 123.700 ;
        RECT 97.940 122.660 99.250 123.970 ;
        RECT 100.380 123.480 100.710 124.470 ;
      LAYER li1 ;
        RECT 101.410 124.300 101.830 124.630 ;
        RECT 102.020 124.240 102.190 124.810 ;
      LAYER li1 ;
        RECT 103.080 124.710 103.250 125.730 ;
        RECT 103.430 125.770 104.530 125.800 ;
        RECT 103.430 125.600 103.480 125.770 ;
        RECT 103.650 125.600 103.840 125.770 ;
        RECT 104.010 125.600 104.200 125.770 ;
        RECT 104.370 125.600 104.530 125.770 ;
        RECT 105.290 125.770 106.900 125.800 ;
        RECT 103.430 124.890 104.530 125.600 ;
        RECT 104.700 124.710 104.950 125.640 ;
        RECT 105.290 125.600 105.340 125.770 ;
        RECT 105.510 125.600 105.780 125.770 ;
        RECT 105.950 125.600 106.220 125.770 ;
        RECT 106.390 125.600 106.630 125.770 ;
        RECT 106.800 125.600 106.900 125.770 ;
        RECT 105.290 125.320 106.900 125.600 ;
      LAYER li1 ;
        RECT 102.370 124.420 102.880 124.630 ;
      LAYER li1 ;
        RECT 103.080 124.540 104.950 124.710 ;
        RECT 105.600 124.920 106.900 125.320 ;
        RECT 107.130 125.770 107.720 125.800 ;
        RECT 107.130 125.600 107.160 125.770 ;
        RECT 107.330 125.600 107.520 125.770 ;
        RECT 107.690 125.600 107.720 125.770 ;
        RECT 108.650 125.770 110.260 125.800 ;
      LAYER li1 ;
        RECT 102.020 124.070 103.080 124.240 ;
        RECT 102.810 123.990 103.080 124.070 ;
        RECT 103.530 124.050 104.040 124.360 ;
        RECT 104.290 124.050 105.000 124.360 ;
      LAYER li1 ;
        RECT 105.600 124.140 105.930 124.920 ;
        RECT 107.130 124.840 107.720 125.600 ;
        RECT 97.940 122.490 97.970 122.660 ;
        RECT 98.140 122.490 98.330 122.660 ;
        RECT 98.500 122.490 98.690 122.660 ;
        RECT 98.860 122.490 99.050 122.660 ;
        RECT 99.220 122.490 99.250 122.660 ;
        RECT 97.940 122.430 99.250 122.490 ;
        RECT 99.610 122.610 101.060 123.480 ;
        RECT 99.610 122.440 99.860 122.610 ;
        RECT 100.030 122.440 100.220 122.610 ;
        RECT 100.390 122.440 100.660 122.610 ;
        RECT 100.830 122.440 101.060 122.610 ;
        RECT 99.610 122.410 101.060 122.440 ;
        RECT 101.370 122.660 102.630 123.890 ;
      LAYER li1 ;
        RECT 102.810 122.910 103.330 123.990 ;
      LAYER li1 ;
        RECT 101.370 122.490 101.380 122.660 ;
        RECT 101.550 122.490 101.740 122.660 ;
        RECT 101.910 122.490 102.100 122.660 ;
        RECT 102.270 122.490 102.460 122.660 ;
        RECT 101.370 122.410 102.630 122.490 ;
      LAYER li1 ;
        RECT 103.160 122.410 103.330 122.910 ;
      LAYER li1 ;
        RECT 103.590 122.660 104.900 123.870 ;
        RECT 106.140 123.480 106.470 124.470 ;
      LAYER li1 ;
        RECT 107.170 124.230 107.880 124.620 ;
        RECT 108.060 123.990 108.390 125.670 ;
      LAYER li1 ;
        RECT 108.650 125.600 108.700 125.770 ;
        RECT 108.870 125.600 109.140 125.770 ;
        RECT 109.310 125.600 109.580 125.770 ;
        RECT 109.750 125.600 109.990 125.770 ;
        RECT 110.160 125.600 110.260 125.770 ;
        RECT 111.920 125.770 112.870 125.800 ;
        RECT 108.650 125.320 110.260 125.600 ;
        RECT 108.960 124.920 110.260 125.320 ;
        RECT 108.960 124.140 109.290 124.920 ;
        RECT 103.590 122.490 103.620 122.660 ;
        RECT 103.790 122.490 103.980 122.660 ;
        RECT 104.150 122.490 104.340 122.660 ;
        RECT 104.510 122.490 104.700 122.660 ;
        RECT 104.870 122.490 104.900 122.660 ;
        RECT 103.590 122.410 104.900 122.490 ;
        RECT 105.370 122.610 106.820 123.480 ;
        RECT 105.370 122.440 105.620 122.610 ;
        RECT 105.790 122.440 105.980 122.610 ;
        RECT 106.150 122.440 106.420 122.610 ;
        RECT 106.590 122.440 106.820 122.610 ;
        RECT 105.370 122.410 106.820 122.440 ;
        RECT 107.130 122.660 107.720 123.990 ;
        RECT 107.130 122.490 107.160 122.660 ;
        RECT 107.330 122.490 107.520 122.660 ;
        RECT 107.690 122.490 107.720 122.660 ;
        RECT 107.130 122.410 107.720 122.490 ;
      LAYER li1 ;
        RECT 108.000 122.410 108.390 123.990 ;
      LAYER li1 ;
        RECT 109.500 123.480 109.830 124.470 ;
        RECT 111.470 123.810 111.740 125.670 ;
        RECT 111.920 125.600 111.950 125.770 ;
        RECT 112.120 125.600 112.310 125.770 ;
        RECT 112.480 125.600 112.670 125.770 ;
        RECT 112.840 125.600 112.870 125.770 ;
        RECT 113.560 125.770 114.150 125.800 ;
        RECT 111.920 125.170 112.870 125.600 ;
        RECT 113.050 125.170 113.380 125.670 ;
      LAYER li1 ;
        RECT 111.920 124.020 112.250 124.990 ;
      LAYER li1 ;
        RECT 112.600 123.810 112.930 124.310 ;
        RECT 111.470 123.640 112.930 123.810 ;
        RECT 108.730 122.610 110.180 123.480 ;
        RECT 111.470 122.710 111.800 123.640 ;
        RECT 108.730 122.440 108.980 122.610 ;
        RECT 109.150 122.440 109.340 122.610 ;
        RECT 109.510 122.440 109.780 122.610 ;
        RECT 109.950 122.440 110.180 122.610 ;
        RECT 111.990 122.660 112.580 123.440 ;
        RECT 111.990 122.490 112.020 122.660 ;
        RECT 112.190 122.490 112.380 122.660 ;
        RECT 112.550 122.490 112.580 122.660 ;
        RECT 111.990 122.460 112.580 122.490 ;
        RECT 112.760 122.530 112.930 123.640 ;
        RECT 113.110 124.250 113.380 125.170 ;
        RECT 113.560 125.600 113.590 125.770 ;
        RECT 113.760 125.600 113.950 125.770 ;
        RECT 114.120 125.600 114.150 125.770 ;
        RECT 118.520 125.770 119.470 125.800 ;
        RECT 113.560 124.920 114.150 125.600 ;
      LAYER li1 ;
        RECT 114.430 125.540 117.370 125.710 ;
        RECT 114.430 125.330 114.600 125.540 ;
        RECT 114.390 125.160 114.600 125.330 ;
        RECT 114.430 124.550 114.600 125.160 ;
      LAYER li1 ;
        RECT 113.110 124.020 113.640 124.250 ;
        RECT 113.110 122.710 113.360 124.020 ;
      LAYER li1 ;
        RECT 114.060 123.680 114.600 124.550 ;
        RECT 114.780 124.060 115.110 125.360 ;
      LAYER li1 ;
        RECT 115.290 124.840 115.560 125.340 ;
        RECT 116.010 125.090 116.340 125.340 ;
        RECT 116.010 124.920 117.020 125.090 ;
        RECT 115.290 123.850 115.460 124.840 ;
        RECT 116.340 124.250 116.670 124.740 ;
        RECT 115.240 123.680 115.460 123.850 ;
        RECT 115.640 124.020 116.670 124.250 ;
        RECT 116.850 124.690 117.020 124.920 ;
      LAYER li1 ;
        RECT 117.200 125.040 117.370 125.540 ;
      LAYER li1 ;
        RECT 118.520 125.600 118.550 125.770 ;
        RECT 118.720 125.600 118.910 125.770 ;
        RECT 119.080 125.600 119.270 125.770 ;
        RECT 119.440 125.600 119.470 125.770 ;
        RECT 118.520 125.220 119.470 125.600 ;
      LAYER li1 ;
        RECT 119.650 125.730 122.310 125.900 ;
        RECT 119.650 125.040 119.820 125.730 ;
        RECT 117.200 124.870 119.820 125.040 ;
      LAYER li1 ;
        RECT 116.850 124.520 119.470 124.690 ;
        RECT 115.240 123.500 115.410 123.680 ;
        RECT 115.640 123.500 115.810 124.020 ;
        RECT 116.850 123.840 117.020 124.520 ;
      LAYER li1 ;
        RECT 119.650 124.340 119.820 124.870 ;
      LAYER li1 ;
        RECT 113.600 123.330 115.410 123.500 ;
        RECT 113.600 122.710 113.850 123.330 ;
        RECT 114.030 122.980 115.060 123.150 ;
        RECT 114.030 122.530 114.200 122.980 ;
        RECT 108.730 122.410 110.180 122.440 ;
        RECT 112.760 122.360 114.200 122.530 ;
        RECT 114.380 122.660 114.710 122.800 ;
        RECT 114.380 122.490 114.410 122.660 ;
        RECT 114.580 122.490 114.710 122.660 ;
        RECT 114.380 122.460 114.710 122.490 ;
        RECT 114.890 122.530 115.060 122.980 ;
        RECT 115.240 122.710 115.410 123.330 ;
        RECT 115.590 123.170 115.810 123.500 ;
        RECT 115.990 123.670 117.020 123.840 ;
        RECT 117.200 123.990 117.530 124.340 ;
      LAYER li1 ;
        RECT 117.970 124.170 119.820 124.340 ;
      LAYER li1 ;
        RECT 120.000 124.840 120.330 125.550 ;
        RECT 120.790 125.380 121.960 125.550 ;
        RECT 120.790 124.840 121.120 125.380 ;
        RECT 120.000 123.990 120.260 124.840 ;
        RECT 121.330 124.580 121.610 125.080 ;
        RECT 117.200 123.820 120.260 123.990 ;
        RECT 115.990 122.970 116.160 123.670 ;
        RECT 116.850 123.640 117.020 123.670 ;
        RECT 116.340 123.290 116.670 123.490 ;
        RECT 116.850 123.470 118.620 123.640 ;
        RECT 116.340 123.170 118.110 123.290 ;
        RECT 116.460 123.120 118.110 123.170 ;
        RECT 115.940 122.710 116.270 122.970 ;
        RECT 116.460 122.530 116.630 123.120 ;
        RECT 114.890 122.360 116.630 122.530 ;
        RECT 116.810 122.660 117.760 122.940 ;
        RECT 116.810 122.490 116.840 122.660 ;
        RECT 117.010 122.490 117.200 122.660 ;
        RECT 117.370 122.490 117.560 122.660 ;
        RECT 117.730 122.490 117.760 122.660 ;
        RECT 116.810 122.460 117.760 122.490 ;
        RECT 117.940 122.530 118.110 123.120 ;
        RECT 118.290 122.710 118.620 123.470 ;
        RECT 119.930 123.240 120.260 123.820 ;
        RECT 120.440 124.410 121.610 124.580 ;
        RECT 120.440 123.060 120.610 124.410 ;
        RECT 120.990 123.730 121.320 124.230 ;
        RECT 121.790 123.980 121.960 125.380 ;
      LAYER li1 ;
        RECT 122.140 125.070 122.310 125.730 ;
      LAYER li1 ;
        RECT 122.490 125.770 123.440 125.800 ;
        RECT 122.490 125.600 122.520 125.770 ;
        RECT 122.690 125.600 122.880 125.770 ;
        RECT 123.050 125.600 123.240 125.770 ;
        RECT 123.410 125.600 123.440 125.770 ;
        RECT 125.100 125.770 126.050 125.800 ;
        RECT 122.490 125.250 123.440 125.600 ;
        RECT 123.980 125.170 124.310 125.670 ;
        RECT 125.100 125.600 125.130 125.770 ;
        RECT 125.300 125.600 125.490 125.770 ;
        RECT 125.660 125.600 125.850 125.770 ;
        RECT 126.020 125.600 126.050 125.770 ;
      LAYER li1 ;
        RECT 122.140 124.900 123.150 125.070 ;
      LAYER li1 ;
        RECT 122.170 124.330 122.500 124.720 ;
      LAYER li1 ;
        RECT 122.820 124.510 123.150 124.900 ;
      LAYER li1 ;
        RECT 123.980 124.330 124.210 125.170 ;
        RECT 124.590 124.670 124.920 125.170 ;
        RECT 125.100 124.670 126.050 125.600 ;
        RECT 127.300 125.780 130.030 125.810 ;
        RECT 127.300 125.610 127.470 125.780 ;
        RECT 127.640 125.610 127.910 125.780 ;
        RECT 128.080 125.610 128.320 125.780 ;
        RECT 128.490 125.610 128.750 125.780 ;
        RECT 128.920 125.610 129.190 125.780 ;
        RECT 129.360 125.610 129.600 125.780 ;
        RECT 129.770 125.610 130.030 125.780 ;
        RECT 122.170 124.160 124.210 124.330 ;
        RECT 121.500 123.810 123.860 123.980 ;
        RECT 121.500 123.490 121.670 123.810 ;
        RECT 124.040 123.630 124.210 124.160 ;
        RECT 118.800 122.890 120.610 123.060 ;
        RECT 120.790 123.320 121.670 123.490 ;
        RECT 118.800 122.530 118.970 122.890 ;
        RECT 117.940 122.360 118.970 122.530 ;
        RECT 119.150 122.660 120.100 122.710 ;
        RECT 119.150 122.490 119.180 122.660 ;
        RECT 119.350 122.490 119.540 122.660 ;
        RECT 119.710 122.490 119.900 122.660 ;
        RECT 120.070 122.490 120.100 122.660 ;
        RECT 119.150 122.410 120.100 122.490 ;
        RECT 120.790 122.410 121.040 123.320 ;
        RECT 121.850 122.660 122.800 123.490 ;
        RECT 123.200 123.460 124.210 123.630 ;
        RECT 124.710 124.490 124.920 124.670 ;
        RECT 124.710 124.160 126.080 124.490 ;
        RECT 123.200 122.990 123.450 123.460 ;
        RECT 123.630 122.660 124.530 123.280 ;
        RECT 124.710 123.160 124.960 124.160 ;
        RECT 121.850 122.490 121.880 122.660 ;
        RECT 122.050 122.490 122.240 122.660 ;
        RECT 122.410 122.490 122.600 122.660 ;
        RECT 122.770 122.490 122.800 122.660 ;
        RECT 123.800 122.490 123.990 122.660 ;
        RECT 124.160 122.490 124.350 122.660 ;
        RECT 124.520 122.490 124.530 122.660 ;
        RECT 121.850 122.460 122.800 122.490 ;
        RECT 123.630 122.460 124.530 122.490 ;
        RECT 125.140 122.660 126.080 123.970 ;
        RECT 125.140 122.490 125.160 122.660 ;
        RECT 125.330 122.490 125.520 122.660 ;
        RECT 125.690 122.490 125.880 122.660 ;
        RECT 126.050 122.490 126.080 122.660 ;
        RECT 125.140 122.430 126.080 122.490 ;
      LAYER li1 ;
        RECT 126.260 122.430 126.600 125.500 ;
      LAYER li1 ;
        RECT 127.300 124.810 130.030 125.610 ;
        RECT 131.140 125.780 133.870 125.810 ;
        RECT 131.140 125.610 131.310 125.780 ;
        RECT 131.480 125.610 131.750 125.780 ;
        RECT 131.920 125.610 132.160 125.780 ;
        RECT 132.330 125.610 132.590 125.780 ;
        RECT 132.760 125.610 133.030 125.780 ;
        RECT 133.200 125.610 133.440 125.780 ;
        RECT 133.610 125.610 133.870 125.780 ;
        RECT 131.140 124.810 133.870 125.610 ;
        RECT 134.980 125.780 137.710 125.810 ;
        RECT 134.980 125.610 135.150 125.780 ;
        RECT 135.320 125.610 135.590 125.780 ;
        RECT 135.760 125.610 136.000 125.780 ;
        RECT 136.170 125.610 136.430 125.780 ;
        RECT 136.600 125.610 136.870 125.780 ;
        RECT 137.040 125.610 137.280 125.780 ;
        RECT 137.450 125.610 137.710 125.780 ;
        RECT 134.980 124.810 137.710 125.610 ;
        RECT 138.820 125.780 141.550 125.810 ;
        RECT 138.820 125.610 138.990 125.780 ;
        RECT 139.160 125.610 139.430 125.780 ;
        RECT 139.600 125.610 139.840 125.780 ;
        RECT 140.010 125.610 140.270 125.780 ;
        RECT 140.440 125.610 140.710 125.780 ;
        RECT 140.880 125.610 141.120 125.780 ;
        RECT 141.290 125.610 141.550 125.780 ;
        RECT 138.820 124.810 141.550 125.610 ;
        RECT 127.460 124.140 127.790 124.810 ;
        RECT 128.190 123.490 128.520 124.470 ;
        RECT 128.740 124.140 129.070 124.810 ;
        RECT 129.470 123.490 129.800 124.470 ;
        RECT 131.300 124.140 131.630 124.810 ;
        RECT 132.030 123.490 132.360 124.470 ;
        RECT 132.580 124.140 132.910 124.810 ;
        RECT 133.310 123.490 133.640 124.470 ;
        RECT 135.140 124.140 135.470 124.810 ;
        RECT 135.870 123.490 136.200 124.470 ;
        RECT 136.420 124.140 136.750 124.810 ;
        RECT 137.150 123.490 137.480 124.470 ;
        RECT 138.980 124.140 139.310 124.810 ;
        RECT 139.710 123.490 140.040 124.470 ;
        RECT 140.260 124.140 140.590 124.810 ;
        RECT 140.990 123.490 141.320 124.470 ;
        RECT 127.220 122.610 129.960 123.490 ;
        RECT 127.220 122.440 127.430 122.610 ;
        RECT 127.600 122.440 127.870 122.610 ;
        RECT 128.040 122.440 128.280 122.610 ;
        RECT 128.450 122.440 128.710 122.610 ;
        RECT 128.880 122.440 129.150 122.610 ;
        RECT 129.320 122.440 129.560 122.610 ;
        RECT 129.730 122.440 129.960 122.610 ;
        RECT 127.220 122.420 129.960 122.440 ;
        RECT 131.060 122.610 133.800 123.490 ;
        RECT 131.060 122.440 131.270 122.610 ;
        RECT 131.440 122.440 131.710 122.610 ;
        RECT 131.880 122.440 132.120 122.610 ;
        RECT 132.290 122.440 132.550 122.610 ;
        RECT 132.720 122.440 132.990 122.610 ;
        RECT 133.160 122.440 133.400 122.610 ;
        RECT 133.570 122.440 133.800 122.610 ;
        RECT 131.060 122.420 133.800 122.440 ;
        RECT 134.900 122.610 137.640 123.490 ;
        RECT 134.900 122.440 135.110 122.610 ;
        RECT 135.280 122.440 135.550 122.610 ;
        RECT 135.720 122.440 135.960 122.610 ;
        RECT 136.130 122.440 136.390 122.610 ;
        RECT 136.560 122.440 136.830 122.610 ;
        RECT 137.000 122.440 137.240 122.610 ;
        RECT 137.410 122.440 137.640 122.610 ;
        RECT 134.900 122.420 137.640 122.440 ;
        RECT 138.740 122.610 141.480 123.490 ;
        RECT 138.740 122.440 138.950 122.610 ;
        RECT 139.120 122.440 139.390 122.610 ;
        RECT 139.560 122.440 139.800 122.610 ;
        RECT 139.970 122.440 140.230 122.610 ;
        RECT 140.400 122.440 140.670 122.610 ;
        RECT 140.840 122.440 141.080 122.610 ;
        RECT 141.250 122.440 141.480 122.610 ;
        RECT 138.740 122.420 141.480 122.440 ;
        RECT 5.760 122.010 5.920 122.190 ;
        RECT 6.090 122.010 6.400 122.190 ;
        RECT 6.570 122.010 6.880 122.190 ;
        RECT 7.050 122.010 7.360 122.190 ;
        RECT 7.530 122.020 7.840 122.190 ;
        RECT 8.010 122.020 8.320 122.190 ;
        RECT 7.530 122.010 7.680 122.020 ;
        RECT 8.160 122.010 8.320 122.020 ;
        RECT 8.490 122.010 8.800 122.190 ;
        RECT 8.970 122.010 9.280 122.190 ;
        RECT 9.450 122.010 9.760 122.190 ;
        RECT 9.930 122.010 10.240 122.190 ;
        RECT 10.410 122.180 10.560 122.190 ;
        RECT 11.040 122.180 11.200 122.190 ;
        RECT 10.410 122.010 10.720 122.180 ;
        RECT 10.890 122.010 11.200 122.180 ;
        RECT 11.370 122.010 11.680 122.190 ;
        RECT 11.850 122.010 12.160 122.190 ;
        RECT 12.330 122.010 12.640 122.190 ;
        RECT 12.810 122.010 13.120 122.190 ;
        RECT 13.290 122.010 13.600 122.190 ;
        RECT 13.770 122.010 14.080 122.190 ;
        RECT 14.250 122.010 14.560 122.190 ;
        RECT 14.730 122.010 15.040 122.190 ;
        RECT 15.210 122.010 15.520 122.190 ;
        RECT 15.690 122.010 16.000 122.190 ;
        RECT 16.170 122.010 16.480 122.190 ;
        RECT 16.650 122.010 16.960 122.190 ;
        RECT 17.130 122.010 17.440 122.190 ;
        RECT 17.610 122.010 17.920 122.190 ;
        RECT 18.090 122.010 18.400 122.190 ;
        RECT 18.570 122.010 18.880 122.190 ;
        RECT 19.050 122.010 19.360 122.190 ;
        RECT 19.530 122.010 19.840 122.190 ;
        RECT 20.010 122.010 20.320 122.190 ;
        RECT 20.490 122.010 20.800 122.190 ;
        RECT 20.970 122.010 21.280 122.190 ;
        RECT 21.450 122.010 21.760 122.190 ;
        RECT 21.930 122.010 22.240 122.190 ;
        RECT 22.410 122.010 22.720 122.190 ;
        RECT 22.890 122.010 23.200 122.190 ;
        RECT 23.370 122.010 23.680 122.190 ;
        RECT 23.850 122.010 24.160 122.190 ;
        RECT 24.330 122.010 24.640 122.190 ;
        RECT 24.810 122.010 25.120 122.190 ;
        RECT 25.290 122.010 25.600 122.190 ;
        RECT 25.770 122.010 26.080 122.190 ;
        RECT 26.250 122.010 26.560 122.190 ;
        RECT 26.730 122.010 27.040 122.190 ;
        RECT 27.210 122.010 27.520 122.190 ;
        RECT 27.690 122.010 28.000 122.190 ;
        RECT 28.170 122.020 28.320 122.190 ;
        RECT 28.800 122.020 28.960 122.190 ;
        RECT 28.170 122.010 28.480 122.020 ;
        RECT 28.650 122.010 28.960 122.020 ;
        RECT 29.130 122.010 29.440 122.190 ;
        RECT 29.610 122.010 29.920 122.190 ;
        RECT 30.090 122.010 30.400 122.190 ;
        RECT 30.570 122.010 30.880 122.190 ;
        RECT 31.050 122.010 31.360 122.190 ;
        RECT 31.530 122.010 31.840 122.190 ;
        RECT 32.010 122.010 32.320 122.190 ;
        RECT 32.490 122.010 32.800 122.190 ;
        RECT 32.970 122.010 33.280 122.190 ;
        RECT 33.450 122.010 33.760 122.190 ;
        RECT 33.930 122.010 34.240 122.190 ;
        RECT 34.410 122.010 34.720 122.190 ;
        RECT 34.890 122.010 35.200 122.190 ;
        RECT 35.370 122.010 35.680 122.190 ;
        RECT 35.850 122.010 36.160 122.190 ;
        RECT 36.330 122.010 36.640 122.190 ;
        RECT 36.810 122.010 37.120 122.190 ;
        RECT 37.290 122.010 37.600 122.190 ;
        RECT 37.770 122.010 38.080 122.190 ;
        RECT 38.250 122.010 38.560 122.190 ;
        RECT 38.730 122.010 39.040 122.190 ;
        RECT 39.210 122.010 39.520 122.190 ;
        RECT 39.690 122.010 40.000 122.190 ;
        RECT 40.170 122.010 40.480 122.190 ;
        RECT 40.650 122.010 40.960 122.190 ;
        RECT 41.130 122.010 41.440 122.190 ;
        RECT 41.610 122.010 41.920 122.190 ;
        RECT 42.090 122.010 42.400 122.190 ;
        RECT 42.570 122.010 42.880 122.190 ;
        RECT 43.050 122.020 43.200 122.190 ;
        RECT 43.680 122.020 43.840 122.190 ;
        RECT 44.010 122.020 44.320 122.190 ;
        RECT 43.050 122.010 43.360 122.020 ;
        RECT 43.530 122.010 43.680 122.020 ;
        RECT 44.160 122.010 44.320 122.020 ;
        RECT 44.490 122.010 44.800 122.190 ;
        RECT 44.970 122.010 45.280 122.190 ;
        RECT 45.450 122.010 45.760 122.190 ;
        RECT 45.930 122.010 46.240 122.190 ;
        RECT 46.410 122.010 46.720 122.190 ;
        RECT 46.890 122.010 47.200 122.190 ;
        RECT 47.370 122.010 47.680 122.190 ;
        RECT 47.850 122.010 48.160 122.190 ;
        RECT 48.330 122.010 48.640 122.190 ;
        RECT 48.810 122.010 49.120 122.190 ;
        RECT 49.290 122.010 49.600 122.190 ;
        RECT 49.770 122.020 49.920 122.190 ;
        RECT 50.400 122.020 50.560 122.190 ;
        RECT 49.770 122.010 50.080 122.020 ;
        RECT 50.250 122.010 50.560 122.020 ;
        RECT 50.730 122.010 51.040 122.190 ;
        RECT 51.210 122.010 51.520 122.190 ;
        RECT 51.690 122.010 52.000 122.190 ;
        RECT 52.170 122.010 52.480 122.190 ;
        RECT 52.650 122.010 52.960 122.190 ;
        RECT 53.130 122.010 53.440 122.190 ;
        RECT 53.610 122.010 53.920 122.190 ;
        RECT 54.090 122.010 54.400 122.190 ;
        RECT 54.570 122.010 54.880 122.190 ;
        RECT 55.050 122.010 55.360 122.190 ;
        RECT 55.530 122.010 55.840 122.190 ;
        RECT 56.010 122.010 56.320 122.190 ;
        RECT 56.490 122.010 56.800 122.190 ;
        RECT 56.970 122.010 57.280 122.190 ;
        RECT 57.450 122.010 57.760 122.190 ;
        RECT 57.930 122.010 58.240 122.190 ;
        RECT 58.410 122.010 58.720 122.190 ;
        RECT 58.890 122.010 59.200 122.190 ;
        RECT 59.370 122.010 59.680 122.190 ;
        RECT 59.850 122.010 60.160 122.190 ;
        RECT 60.330 122.010 60.640 122.190 ;
        RECT 60.810 122.010 61.120 122.190 ;
        RECT 61.290 122.010 61.600 122.190 ;
        RECT 61.770 122.010 62.080 122.190 ;
        RECT 62.250 122.010 62.560 122.190 ;
        RECT 62.730 122.010 63.040 122.190 ;
        RECT 63.210 122.010 63.520 122.190 ;
        RECT 63.690 122.010 64.000 122.190 ;
        RECT 64.170 122.010 64.480 122.190 ;
        RECT 64.650 122.010 64.960 122.190 ;
        RECT 65.130 122.010 65.440 122.190 ;
        RECT 65.610 122.010 65.920 122.190 ;
        RECT 66.090 122.010 66.400 122.190 ;
        RECT 66.570 122.010 66.880 122.190 ;
        RECT 67.050 122.180 67.200 122.190 ;
        RECT 67.680 122.180 67.840 122.190 ;
        RECT 67.050 122.010 67.360 122.180 ;
        RECT 67.530 122.010 67.840 122.180 ;
        RECT 68.010 122.010 68.320 122.190 ;
        RECT 68.490 122.010 68.800 122.190 ;
        RECT 68.970 122.010 69.280 122.190 ;
        RECT 69.450 122.010 69.760 122.190 ;
        RECT 69.930 122.010 70.240 122.190 ;
        RECT 70.410 122.010 70.720 122.190 ;
        RECT 70.890 122.010 71.200 122.190 ;
        RECT 71.370 122.010 71.680 122.190 ;
        RECT 71.850 122.010 72.160 122.190 ;
        RECT 72.330 122.010 72.640 122.190 ;
        RECT 72.810 122.010 73.120 122.190 ;
        RECT 73.290 122.010 73.600 122.190 ;
        RECT 73.770 122.010 74.080 122.190 ;
        RECT 74.250 122.010 74.560 122.190 ;
        RECT 74.730 122.010 75.040 122.190 ;
        RECT 75.210 122.010 75.520 122.190 ;
        RECT 75.690 122.010 76.000 122.190 ;
        RECT 76.170 122.010 76.480 122.190 ;
        RECT 76.650 122.010 76.960 122.190 ;
        RECT 77.130 122.010 77.440 122.190 ;
        RECT 77.610 122.010 77.920 122.190 ;
        RECT 78.090 122.010 78.400 122.190 ;
        RECT 78.570 122.010 78.880 122.190 ;
        RECT 79.050 122.010 79.360 122.190 ;
        RECT 79.530 122.010 79.840 122.190 ;
        RECT 80.010 122.010 80.320 122.190 ;
        RECT 80.490 122.010 80.800 122.190 ;
        RECT 80.970 122.010 81.280 122.190 ;
        RECT 81.450 122.010 81.760 122.190 ;
        RECT 81.930 122.010 82.240 122.190 ;
        RECT 82.410 122.010 82.720 122.190 ;
        RECT 82.890 122.010 83.200 122.190 ;
        RECT 83.370 122.010 83.680 122.190 ;
        RECT 83.850 122.010 84.160 122.190 ;
        RECT 84.330 122.010 84.640 122.190 ;
        RECT 84.810 122.010 85.120 122.190 ;
        RECT 85.290 122.010 85.600 122.190 ;
        RECT 85.770 122.010 86.080 122.190 ;
        RECT 86.250 122.010 86.560 122.190 ;
        RECT 86.730 122.010 87.040 122.190 ;
        RECT 87.210 122.010 87.520 122.190 ;
        RECT 87.690 122.010 88.000 122.190 ;
        RECT 88.170 122.010 88.480 122.190 ;
        RECT 88.650 122.010 88.960 122.190 ;
        RECT 89.130 122.010 89.440 122.190 ;
        RECT 89.610 122.010 89.920 122.190 ;
        RECT 90.090 122.010 90.400 122.190 ;
        RECT 90.570 122.010 90.880 122.190 ;
        RECT 91.050 122.010 91.360 122.190 ;
        RECT 91.530 122.010 91.840 122.190 ;
        RECT 92.010 122.010 92.320 122.190 ;
        RECT 92.490 122.010 92.800 122.190 ;
        RECT 92.970 122.010 93.280 122.190 ;
        RECT 93.450 122.010 93.760 122.190 ;
        RECT 93.930 122.010 94.240 122.190 ;
        RECT 94.410 122.010 94.720 122.190 ;
        RECT 94.890 122.010 95.200 122.190 ;
        RECT 95.370 122.010 95.680 122.190 ;
        RECT 95.850 122.010 96.160 122.190 ;
        RECT 96.330 122.010 96.640 122.190 ;
        RECT 96.810 122.010 97.120 122.190 ;
        RECT 97.290 122.010 97.600 122.190 ;
        RECT 97.770 122.010 98.080 122.190 ;
        RECT 98.250 122.010 98.560 122.190 ;
        RECT 98.730 122.010 99.040 122.190 ;
        RECT 99.210 122.010 99.520 122.190 ;
        RECT 99.690 122.010 100.000 122.190 ;
        RECT 100.170 122.020 100.320 122.190 ;
        RECT 100.800 122.020 100.960 122.190 ;
        RECT 100.170 122.010 100.480 122.020 ;
        RECT 100.650 122.010 100.960 122.020 ;
        RECT 101.130 122.010 101.440 122.190 ;
        RECT 101.610 122.010 101.920 122.190 ;
        RECT 102.090 122.010 102.400 122.190 ;
        RECT 102.570 122.010 102.880 122.190 ;
        RECT 103.050 122.010 103.360 122.190 ;
        RECT 103.530 122.010 103.840 122.190 ;
        RECT 104.010 122.010 104.320 122.190 ;
        RECT 104.490 122.010 104.800 122.190 ;
        RECT 104.970 122.010 105.280 122.190 ;
        RECT 105.450 122.010 105.760 122.190 ;
        RECT 105.930 122.010 106.240 122.190 ;
        RECT 106.410 122.010 106.720 122.190 ;
        RECT 106.890 122.010 107.200 122.190 ;
        RECT 107.370 122.010 107.680 122.190 ;
        RECT 107.850 122.010 108.160 122.190 ;
        RECT 108.330 122.010 108.640 122.190 ;
        RECT 108.810 122.010 109.120 122.190 ;
        RECT 109.290 122.010 109.600 122.190 ;
        RECT 109.770 122.010 110.080 122.190 ;
        RECT 110.250 122.010 110.560 122.190 ;
        RECT 110.730 122.010 111.040 122.190 ;
        RECT 111.210 122.010 111.520 122.190 ;
        RECT 111.690 122.010 112.000 122.190 ;
        RECT 112.170 122.010 112.480 122.190 ;
        RECT 112.650 122.010 112.960 122.190 ;
        RECT 113.130 122.010 113.440 122.190 ;
        RECT 113.610 122.010 113.920 122.190 ;
        RECT 114.090 122.010 114.400 122.190 ;
        RECT 114.570 122.010 114.880 122.190 ;
        RECT 115.050 122.010 115.360 122.190 ;
        RECT 115.530 122.010 115.840 122.190 ;
        RECT 116.010 122.010 116.320 122.190 ;
        RECT 116.490 122.010 116.800 122.190 ;
        RECT 116.970 122.010 117.280 122.190 ;
        RECT 117.450 122.010 117.760 122.190 ;
        RECT 117.930 122.010 118.240 122.190 ;
        RECT 118.410 122.010 118.720 122.190 ;
        RECT 118.890 122.010 119.200 122.190 ;
        RECT 119.370 122.010 119.680 122.190 ;
        RECT 119.850 122.010 120.160 122.190 ;
        RECT 120.330 122.010 120.640 122.190 ;
        RECT 120.810 122.010 121.120 122.190 ;
        RECT 121.290 122.010 121.600 122.190 ;
        RECT 121.770 122.010 122.080 122.190 ;
        RECT 122.250 122.010 122.560 122.190 ;
        RECT 122.730 122.010 123.040 122.190 ;
        RECT 123.210 122.010 123.520 122.190 ;
        RECT 123.690 122.010 124.000 122.190 ;
        RECT 124.170 122.010 124.480 122.190 ;
        RECT 124.650 122.010 124.960 122.190 ;
        RECT 125.130 122.010 125.440 122.190 ;
        RECT 125.610 122.010 125.920 122.190 ;
        RECT 126.090 122.010 126.400 122.190 ;
        RECT 126.570 122.010 126.880 122.190 ;
        RECT 127.050 122.010 127.360 122.190 ;
        RECT 127.530 122.010 127.840 122.190 ;
        RECT 128.010 122.010 128.320 122.190 ;
        RECT 128.490 122.010 128.800 122.190 ;
        RECT 128.970 122.010 129.280 122.190 ;
        RECT 129.450 122.010 129.760 122.190 ;
        RECT 129.930 122.010 130.240 122.190 ;
        RECT 130.410 122.010 130.720 122.190 ;
        RECT 130.890 122.010 131.200 122.190 ;
        RECT 131.370 122.010 131.680 122.190 ;
        RECT 131.850 122.010 132.160 122.190 ;
        RECT 132.330 122.010 132.640 122.190 ;
        RECT 132.810 122.010 133.120 122.190 ;
        RECT 133.290 122.010 133.600 122.190 ;
        RECT 133.770 122.010 134.080 122.190 ;
        RECT 134.250 122.010 134.560 122.190 ;
        RECT 134.730 122.010 135.040 122.190 ;
        RECT 135.210 122.010 135.520 122.190 ;
        RECT 135.690 122.010 136.000 122.190 ;
        RECT 136.170 122.010 136.480 122.190 ;
        RECT 136.650 122.010 136.960 122.190 ;
        RECT 137.130 122.010 137.440 122.190 ;
        RECT 137.610 122.010 137.920 122.190 ;
        RECT 138.090 122.010 138.400 122.190 ;
        RECT 138.570 122.010 138.880 122.190 ;
        RECT 139.050 122.010 139.360 122.190 ;
        RECT 139.530 122.010 139.840 122.190 ;
        RECT 140.010 122.010 140.320 122.190 ;
        RECT 140.490 122.010 140.800 122.190 ;
        RECT 140.970 122.010 141.280 122.190 ;
        RECT 141.450 122.180 141.600 122.190 ;
        RECT 141.450 122.010 141.760 122.180 ;
        RECT 141.930 122.010 142.080 122.180 ;
        RECT 6.260 121.760 9.000 121.780 ;
        RECT 6.260 121.590 6.470 121.760 ;
        RECT 6.640 121.590 6.910 121.760 ;
        RECT 7.080 121.590 7.320 121.760 ;
        RECT 7.490 121.590 7.750 121.760 ;
        RECT 7.920 121.590 8.190 121.760 ;
        RECT 8.360 121.590 8.600 121.760 ;
        RECT 8.770 121.590 9.000 121.760 ;
        RECT 6.260 120.710 9.000 121.590 ;
        RECT 11.130 121.710 11.720 121.790 ;
        RECT 11.130 121.540 11.160 121.710 ;
        RECT 11.330 121.540 11.520 121.710 ;
        RECT 11.690 121.540 11.720 121.710 ;
        RECT 6.500 119.390 6.830 120.060 ;
        RECT 7.230 119.730 7.560 120.710 ;
        RECT 7.780 119.390 8.110 120.060 ;
        RECT 8.510 119.730 8.840 120.710 ;
        RECT 11.130 120.210 11.720 121.540 ;
      LAYER li1 ;
        RECT 12.000 120.210 12.390 121.790 ;
      LAYER li1 ;
        RECT 12.980 121.760 15.720 121.780 ;
        RECT 12.980 121.590 13.190 121.760 ;
        RECT 13.360 121.590 13.630 121.760 ;
        RECT 13.800 121.590 14.040 121.760 ;
        RECT 14.210 121.590 14.470 121.760 ;
        RECT 14.640 121.590 14.910 121.760 ;
        RECT 15.080 121.590 15.320 121.760 ;
        RECT 15.490 121.590 15.720 121.760 ;
        RECT 12.980 120.710 15.720 121.590 ;
        RECT 16.820 121.760 19.560 121.780 ;
        RECT 16.820 121.590 17.030 121.760 ;
        RECT 17.200 121.590 17.470 121.760 ;
        RECT 17.640 121.590 17.880 121.760 ;
        RECT 18.050 121.590 18.310 121.760 ;
        RECT 18.480 121.590 18.750 121.760 ;
        RECT 18.920 121.590 19.160 121.760 ;
        RECT 19.330 121.590 19.560 121.760 ;
        RECT 16.820 120.710 19.560 121.590 ;
        RECT 6.340 118.390 9.070 119.390 ;
        RECT 11.130 118.400 11.720 119.360 ;
      LAYER li1 ;
        RECT 12.060 118.530 12.390 120.210 ;
      LAYER li1 ;
        RECT 13.220 119.390 13.550 120.060 ;
        RECT 13.950 119.730 14.280 120.710 ;
        RECT 14.500 119.390 14.830 120.060 ;
        RECT 15.230 119.730 15.560 120.710 ;
        RECT 17.060 119.390 17.390 120.060 ;
        RECT 17.790 119.730 18.120 120.710 ;
        RECT 18.340 119.390 18.670 120.060 ;
        RECT 19.070 119.730 19.400 120.710 ;
        RECT 13.060 118.390 15.790 119.390 ;
        RECT 16.900 118.390 19.630 119.390 ;
      LAYER li1 ;
        RECT 20.270 118.530 20.540 121.790 ;
      LAYER li1 ;
        RECT 20.720 121.710 21.620 121.790 ;
        RECT 20.720 121.540 20.730 121.710 ;
        RECT 20.900 121.540 21.090 121.710 ;
        RECT 21.260 121.540 21.450 121.710 ;
        RECT 21.800 121.670 23.690 121.840 ;
        RECT 20.720 120.210 21.620 121.540 ;
        RECT 21.800 120.210 21.970 121.670 ;
      LAYER li1 ;
        RECT 22.150 119.810 22.480 121.290 ;
      LAYER li1 ;
        RECT 20.750 119.630 21.080 119.790 ;
        RECT 22.660 119.630 22.990 121.490 ;
        RECT 23.440 120.130 23.690 121.670 ;
        RECT 23.870 121.710 24.820 121.790 ;
        RECT 23.870 121.540 23.900 121.710 ;
        RECT 24.070 121.540 24.260 121.710 ;
        RECT 24.430 121.540 24.620 121.710 ;
        RECT 24.790 121.540 24.820 121.710 ;
        RECT 23.870 120.310 24.820 121.540 ;
        RECT 25.000 120.130 25.330 121.770 ;
        RECT 25.690 121.760 27.140 121.790 ;
        RECT 25.690 121.590 25.940 121.760 ;
        RECT 26.110 121.590 26.300 121.760 ;
        RECT 26.470 121.590 26.740 121.760 ;
        RECT 26.910 121.590 27.140 121.760 ;
        RECT 25.690 120.720 27.140 121.590 ;
        RECT 23.440 119.960 25.330 120.130 ;
        RECT 20.750 119.460 23.020 119.630 ;
        RECT 20.710 118.400 22.420 119.280 ;
        RECT 22.850 118.660 23.020 119.460 ;
      LAYER li1 ;
        RECT 23.200 119.040 23.370 119.780 ;
        RECT 23.650 119.540 24.810 119.780 ;
        RECT 24.990 119.540 25.320 119.780 ;
        RECT 23.190 118.870 23.370 119.040 ;
        RECT 23.200 118.840 23.370 118.870 ;
      LAYER li1 ;
        RECT 23.550 118.660 23.800 119.360 ;
        RECT 22.850 118.490 23.800 118.660 ;
        RECT 23.980 118.400 25.290 119.360 ;
        RECT 25.920 119.280 26.250 120.060 ;
        RECT 26.460 119.730 26.790 120.720 ;
        RECT 25.920 118.880 27.220 119.280 ;
        RECT 25.610 118.400 27.220 118.880 ;
      LAYER li1 ;
        RECT 28.910 118.530 29.180 121.790 ;
      LAYER li1 ;
        RECT 29.360 121.710 30.260 121.790 ;
        RECT 29.360 121.540 29.370 121.710 ;
        RECT 29.540 121.540 29.730 121.710 ;
        RECT 29.900 121.540 30.090 121.710 ;
        RECT 30.440 121.670 32.330 121.840 ;
        RECT 29.360 120.210 30.260 121.540 ;
        RECT 30.440 120.210 30.610 121.670 ;
      LAYER li1 ;
        RECT 30.790 119.810 31.120 121.290 ;
      LAYER li1 ;
        RECT 29.390 119.630 29.720 119.790 ;
        RECT 31.300 119.630 31.630 121.490 ;
        RECT 32.080 120.130 32.330 121.670 ;
        RECT 32.510 121.710 33.460 121.790 ;
        RECT 32.510 121.540 32.540 121.710 ;
        RECT 32.710 121.540 32.900 121.710 ;
        RECT 33.070 121.540 33.260 121.710 ;
        RECT 33.430 121.540 33.460 121.710 ;
        RECT 32.510 120.310 33.460 121.540 ;
        RECT 33.640 120.130 33.970 121.770 ;
        RECT 34.330 121.760 35.780 121.790 ;
        RECT 34.330 121.590 34.580 121.760 ;
        RECT 34.750 121.590 34.940 121.760 ;
        RECT 35.110 121.590 35.380 121.760 ;
        RECT 35.550 121.590 35.780 121.760 ;
        RECT 34.330 120.720 35.780 121.590 ;
        RECT 32.080 119.960 33.970 120.130 ;
        RECT 29.390 119.460 31.660 119.630 ;
      LAYER li1 ;
        RECT 31.830 119.610 32.010 119.780 ;
      LAYER li1 ;
        RECT 29.350 118.400 31.060 119.280 ;
        RECT 31.490 118.660 31.660 119.460 ;
      LAYER li1 ;
        RECT 31.840 118.840 32.010 119.610 ;
        RECT 32.290 119.540 33.450 119.780 ;
        RECT 33.630 119.540 33.960 119.780 ;
      LAYER li1 ;
        RECT 32.190 118.660 32.440 119.360 ;
        RECT 31.490 118.490 32.440 118.660 ;
        RECT 32.620 118.400 33.930 119.360 ;
        RECT 34.560 119.280 34.890 120.060 ;
        RECT 35.100 119.730 35.430 120.720 ;
      LAYER li1 ;
        RECT 36.120 120.210 36.550 121.790 ;
      LAYER li1 ;
        RECT 36.730 121.710 37.290 121.790 ;
        RECT 36.730 121.540 36.740 121.710 ;
        RECT 36.910 121.540 37.100 121.710 ;
        RECT 37.270 121.540 37.290 121.710 ;
        RECT 36.730 120.210 37.290 121.540 ;
        RECT 38.900 121.760 41.640 121.780 ;
        RECT 38.900 121.590 39.110 121.760 ;
        RECT 39.280 121.590 39.550 121.760 ;
        RECT 39.720 121.590 39.960 121.760 ;
        RECT 40.130 121.590 40.390 121.760 ;
        RECT 40.560 121.590 40.830 121.760 ;
        RECT 41.000 121.590 41.240 121.760 ;
        RECT 41.410 121.590 41.640 121.760 ;
        RECT 34.560 118.880 35.860 119.280 ;
        RECT 34.250 118.400 35.860 118.880 ;
      LAYER li1 ;
        RECT 36.120 118.530 36.370 120.210 ;
      LAYER li1 ;
        RECT 36.680 119.320 37.010 119.780 ;
      LAYER li1 ;
        RECT 37.470 119.500 37.800 121.290 ;
      LAYER li1 ;
        RECT 37.980 119.320 38.230 121.040 ;
        RECT 38.900 120.710 41.640 121.590 ;
        RECT 39.140 119.390 39.470 120.060 ;
        RECT 39.870 119.730 40.200 120.710 ;
        RECT 40.420 119.390 40.750 120.060 ;
        RECT 41.150 119.730 41.480 120.710 ;
      LAYER li1 ;
        RECT 43.800 120.210 44.230 121.790 ;
      LAYER li1 ;
        RECT 44.410 121.710 44.970 121.790 ;
        RECT 44.410 121.540 44.420 121.710 ;
        RECT 44.590 121.540 44.780 121.710 ;
        RECT 44.950 121.540 44.970 121.710 ;
        RECT 44.410 120.210 44.970 121.540 ;
        RECT 46.580 121.760 49.320 121.780 ;
        RECT 46.580 121.590 46.790 121.760 ;
        RECT 46.960 121.590 47.230 121.760 ;
        RECT 47.400 121.590 47.640 121.760 ;
        RECT 47.810 121.590 48.070 121.760 ;
        RECT 48.240 121.590 48.510 121.760 ;
        RECT 48.680 121.590 48.920 121.760 ;
        RECT 49.090 121.590 49.320 121.760 ;
        RECT 36.680 119.150 38.230 119.320 ;
        RECT 36.550 118.400 37.800 118.970 ;
        RECT 37.980 118.530 38.230 119.150 ;
        RECT 38.980 118.390 41.710 119.390 ;
      LAYER li1 ;
        RECT 43.800 118.530 44.050 120.210 ;
      LAYER li1 ;
        RECT 44.360 119.320 44.690 119.780 ;
      LAYER li1 ;
        RECT 45.150 119.500 45.480 121.290 ;
      LAYER li1 ;
        RECT 45.660 119.320 45.910 121.040 ;
        RECT 46.580 120.710 49.320 121.590 ;
        RECT 46.820 119.390 47.150 120.060 ;
        RECT 47.550 119.730 47.880 120.710 ;
        RECT 48.100 119.390 48.430 120.060 ;
        RECT 48.830 119.730 49.160 120.710 ;
        RECT 50.520 119.500 50.770 121.770 ;
        RECT 50.950 121.710 51.900 121.790 ;
        RECT 50.950 121.540 50.980 121.710 ;
        RECT 51.150 121.540 51.340 121.710 ;
        RECT 51.510 121.540 51.700 121.710 ;
        RECT 51.870 121.540 51.900 121.710 ;
        RECT 50.950 120.960 51.900 121.540 ;
        RECT 52.080 120.980 52.410 121.770 ;
        RECT 52.090 120.480 52.410 120.980 ;
        RECT 52.640 121.710 52.890 121.740 ;
        RECT 52.640 121.540 52.670 121.710 ;
        RECT 52.840 121.540 52.890 121.710 ;
        RECT 52.640 120.660 52.890 121.540 ;
        RECT 53.070 120.480 53.240 121.790 ;
        RECT 56.010 121.710 56.340 121.740 ;
        RECT 52.090 120.310 53.240 120.480 ;
        RECT 53.420 121.320 55.410 121.650 ;
        RECT 51.580 119.500 51.910 119.930 ;
        RECT 44.360 119.150 45.910 119.320 ;
        RECT 44.230 118.400 45.480 118.970 ;
        RECT 45.660 118.530 45.910 119.150 ;
        RECT 46.660 118.390 49.390 119.390 ;
        RECT 50.520 119.330 51.910 119.500 ;
        RECT 50.520 118.650 50.780 119.330 ;
        RECT 50.970 118.400 51.560 119.150 ;
        RECT 51.740 118.470 51.910 119.330 ;
        RECT 52.090 118.650 52.340 120.310 ;
      LAYER li1 ;
        RECT 52.910 119.560 53.240 120.130 ;
      LAYER li1 ;
        RECT 53.420 119.380 53.590 121.320 ;
        RECT 52.520 119.210 53.590 119.380 ;
        RECT 52.520 118.470 52.690 119.210 ;
        RECT 53.770 119.030 53.940 121.140 ;
        RECT 54.120 119.120 54.290 121.320 ;
        RECT 54.470 120.640 54.800 121.140 ;
        RECT 54.470 119.170 54.640 120.640 ;
        RECT 55.240 120.360 55.410 121.320 ;
        RECT 55.590 120.710 55.830 121.590 ;
        RECT 56.010 121.540 56.040 121.710 ;
        RECT 56.210 121.540 56.340 121.710 ;
        RECT 56.010 120.890 56.340 121.540 ;
        RECT 57.480 121.710 58.430 121.740 ;
        RECT 57.480 121.540 57.510 121.710 ;
        RECT 57.680 121.540 57.870 121.710 ;
        RECT 58.040 121.540 58.230 121.710 ;
        RECT 58.400 121.540 58.430 121.710 ;
        RECT 56.970 120.880 57.300 121.140 ;
        RECT 56.520 120.710 57.300 120.880 ;
        RECT 57.480 120.710 58.430 121.540 ;
        RECT 59.100 121.630 60.230 121.840 ;
        RECT 60.410 121.710 61.360 121.740 ;
        RECT 59.100 120.880 59.270 121.630 ;
        RECT 60.410 121.540 60.440 121.710 ;
        RECT 60.610 121.540 60.800 121.710 ;
        RECT 60.970 121.540 61.160 121.710 ;
        RECT 61.330 121.540 61.360 121.710 ;
        RECT 59.450 121.060 60.060 121.450 ;
        RECT 59.100 120.710 59.710 120.880 ;
        RECT 55.590 120.540 56.690 120.710 ;
        RECT 56.870 120.360 59.360 120.530 ;
        RECT 54.820 120.010 55.060 120.200 ;
        RECT 55.240 120.190 57.040 120.360 ;
        RECT 57.220 120.010 58.850 120.180 ;
        RECT 59.030 120.120 59.360 120.360 ;
        RECT 54.820 119.840 57.390 120.010 ;
        RECT 58.680 119.910 58.850 120.010 ;
        RECT 59.540 119.910 59.710 120.710 ;
        RECT 54.820 119.530 55.060 119.840 ;
        RECT 55.540 119.350 56.270 119.660 ;
      LAYER li1 ;
        RECT 57.570 119.590 58.500 119.830 ;
      LAYER li1 ;
        RECT 51.740 118.300 52.690 118.470 ;
        RECT 52.870 118.400 53.410 119.030 ;
        RECT 53.590 118.530 53.940 119.030 ;
        RECT 54.470 119.000 56.720 119.170 ;
        RECT 54.470 118.530 54.720 119.000 ;
        RECT 55.260 118.400 56.210 118.820 ;
        RECT 56.390 118.300 56.720 119.000 ;
        RECT 57.200 118.400 58.150 119.410 ;
      LAYER li1 ;
        RECT 58.330 119.040 58.500 119.590 ;
      LAYER li1 ;
        RECT 58.680 119.740 59.710 119.910 ;
        RECT 59.890 120.520 60.060 121.060 ;
        RECT 60.410 120.700 61.360 121.540 ;
        RECT 61.700 121.290 61.950 121.790 ;
        RECT 62.130 121.710 63.080 121.770 ;
        RECT 65.530 121.760 66.980 121.790 ;
        RECT 62.130 121.540 62.160 121.710 ;
        RECT 62.330 121.540 62.520 121.710 ;
        RECT 62.690 121.540 62.880 121.710 ;
        RECT 63.050 121.540 63.080 121.710 ;
        RECT 62.130 121.390 63.080 121.540 ;
        RECT 63.700 121.710 64.640 121.740 ;
        RECT 63.700 121.540 63.720 121.710 ;
        RECT 63.890 121.540 64.080 121.710 ;
        RECT 64.250 121.540 64.440 121.710 ;
        RECT 64.610 121.540 64.640 121.710 ;
        RECT 61.780 121.210 61.950 121.290 ;
        RECT 61.780 121.040 62.960 121.210 ;
        RECT 61.810 120.710 62.140 120.860 ;
        RECT 61.810 120.520 62.610 120.710 ;
        RECT 59.890 120.350 62.610 120.520 ;
        RECT 58.680 119.580 59.190 119.740 ;
        RECT 59.890 119.510 60.060 120.350 ;
        RECT 60.710 119.860 61.040 120.170 ;
        RECT 62.280 120.040 62.610 120.350 ;
        RECT 62.790 119.860 62.960 121.040 ;
        RECT 60.710 119.690 62.960 119.860 ;
        RECT 63.270 120.430 63.520 121.400 ;
        RECT 63.700 120.610 64.640 121.540 ;
        RECT 65.530 121.590 65.780 121.760 ;
        RECT 65.950 121.590 66.140 121.760 ;
        RECT 66.310 121.590 66.580 121.760 ;
        RECT 66.750 121.590 66.980 121.760 ;
        RECT 65.530 120.720 66.980 121.590 ;
        RECT 67.770 121.710 68.360 121.790 ;
        RECT 67.770 121.540 67.800 121.710 ;
        RECT 67.970 121.540 68.160 121.710 ;
        RECT 68.330 121.540 68.360 121.710 ;
        RECT 63.270 120.260 64.640 120.430 ;
        RECT 60.710 119.580 61.040 119.690 ;
        RECT 59.430 119.220 60.060 119.510 ;
      LAYER li1 ;
        RECT 61.290 119.040 61.560 119.070 ;
        RECT 58.330 118.870 61.560 119.040 ;
        RECT 58.690 118.590 61.560 118.870 ;
      LAYER li1 ;
        RECT 61.740 118.400 62.330 119.510 ;
        RECT 62.520 119.010 62.850 119.690 ;
        RECT 63.270 119.510 63.480 120.260 ;
        RECT 64.310 119.760 64.640 120.260 ;
        RECT 63.150 119.010 63.480 119.510 ;
        RECT 63.660 118.400 64.610 119.510 ;
        RECT 65.760 119.280 66.090 120.060 ;
        RECT 66.300 119.730 66.630 120.720 ;
        RECT 67.770 120.210 68.360 121.540 ;
      LAYER li1 ;
        RECT 68.640 120.210 69.030 121.790 ;
      LAYER li1 ;
        RECT 69.620 121.760 72.360 121.780 ;
        RECT 69.620 121.590 69.830 121.760 ;
        RECT 70.000 121.590 70.270 121.760 ;
        RECT 70.440 121.590 70.680 121.760 ;
        RECT 70.850 121.590 71.110 121.760 ;
        RECT 71.280 121.590 71.550 121.760 ;
        RECT 71.720 121.590 71.960 121.760 ;
        RECT 72.130 121.590 72.360 121.760 ;
        RECT 69.620 120.710 72.360 121.590 ;
        RECT 65.760 118.880 67.060 119.280 ;
        RECT 65.450 118.400 67.060 118.880 ;
        RECT 67.770 118.400 68.360 119.360 ;
      LAYER li1 ;
        RECT 68.700 118.530 69.030 120.210 ;
      LAYER li1 ;
        RECT 69.860 119.390 70.190 120.060 ;
        RECT 70.590 119.730 70.920 120.710 ;
        RECT 71.140 119.390 71.470 120.060 ;
        RECT 71.870 119.730 72.200 120.710 ;
      LAYER li1 ;
        RECT 74.040 120.210 74.470 121.790 ;
      LAYER li1 ;
        RECT 74.650 121.710 75.210 121.790 ;
        RECT 74.650 121.540 74.660 121.710 ;
        RECT 74.830 121.540 75.020 121.710 ;
        RECT 75.190 121.540 75.210 121.710 ;
        RECT 74.650 120.210 75.210 121.540 ;
        RECT 76.570 121.760 78.020 121.790 ;
        RECT 76.570 121.590 76.820 121.760 ;
        RECT 76.990 121.590 77.180 121.760 ;
        RECT 77.350 121.590 77.620 121.760 ;
        RECT 77.790 121.590 78.020 121.760 ;
        RECT 69.700 118.390 72.430 119.390 ;
      LAYER li1 ;
        RECT 74.040 118.530 74.290 120.210 ;
      LAYER li1 ;
        RECT 74.600 119.320 74.930 119.780 ;
      LAYER li1 ;
        RECT 75.390 119.500 75.720 121.290 ;
      LAYER li1 ;
        RECT 75.900 119.320 76.150 121.040 ;
        RECT 76.570 120.720 78.020 121.590 ;
        RECT 78.330 121.710 80.000 121.790 ;
        RECT 78.330 121.540 78.360 121.710 ;
        RECT 78.530 121.540 78.720 121.710 ;
        RECT 78.890 121.540 79.080 121.710 ;
        RECT 79.250 121.540 79.440 121.710 ;
        RECT 79.610 121.540 79.800 121.710 ;
        RECT 79.970 121.540 80.000 121.710 ;
        RECT 74.600 119.150 76.150 119.320 ;
        RECT 74.470 118.400 75.720 118.970 ;
        RECT 75.900 118.530 76.150 119.150 ;
        RECT 76.800 119.280 77.130 120.060 ;
        RECT 77.340 119.730 77.670 120.720 ;
        RECT 78.330 120.330 80.000 121.540 ;
      LAYER li1 ;
        RECT 78.370 119.810 79.560 120.150 ;
        RECT 79.740 119.810 80.070 120.150 ;
        RECT 80.260 119.630 80.520 121.790 ;
      LAYER li1 ;
        RECT 80.890 121.760 82.340 121.790 ;
        RECT 80.890 121.590 81.140 121.760 ;
        RECT 81.310 121.590 81.500 121.760 ;
        RECT 81.670 121.590 81.940 121.760 ;
        RECT 82.110 121.590 82.340 121.760 ;
        RECT 80.890 120.720 82.340 121.590 ;
        RECT 82.650 121.710 83.240 121.790 ;
        RECT 82.650 121.540 82.680 121.710 ;
        RECT 82.850 121.540 83.040 121.710 ;
        RECT 83.210 121.540 83.240 121.710 ;
      LAYER li1 ;
        RECT 79.440 119.460 80.520 119.630 ;
      LAYER li1 ;
        RECT 76.800 118.880 78.100 119.280 ;
        RECT 76.490 118.400 78.100 118.880 ;
        RECT 78.330 118.400 79.260 119.360 ;
      LAYER li1 ;
        RECT 79.440 118.530 79.770 119.460 ;
      LAYER li1 ;
        RECT 81.120 119.280 81.450 120.060 ;
        RECT 81.660 119.730 81.990 120.720 ;
        RECT 82.650 120.210 83.240 121.540 ;
      LAYER li1 ;
        RECT 83.520 120.210 83.910 121.790 ;
      LAYER li1 ;
        RECT 84.250 121.760 85.700 121.790 ;
        RECT 84.250 121.590 84.500 121.760 ;
        RECT 84.670 121.590 84.860 121.760 ;
        RECT 85.030 121.590 85.300 121.760 ;
        RECT 85.470 121.590 85.700 121.760 ;
        RECT 84.250 120.720 85.700 121.590 ;
        RECT 86.010 121.710 86.960 121.790 ;
        RECT 86.010 121.540 86.040 121.710 ;
        RECT 86.210 121.540 86.400 121.710 ;
        RECT 86.570 121.540 86.760 121.710 ;
        RECT 86.930 121.540 86.960 121.710 ;
      LAYER li1 ;
        RECT 82.690 119.580 83.400 119.970 ;
      LAYER li1 ;
        RECT 79.960 118.400 80.550 119.280 ;
        RECT 81.120 118.880 82.420 119.280 ;
        RECT 80.810 118.400 82.420 118.880 ;
        RECT 82.650 118.400 83.240 119.360 ;
      LAYER li1 ;
        RECT 83.580 118.530 83.910 120.210 ;
      LAYER li1 ;
        RECT 84.480 119.280 84.810 120.060 ;
        RECT 85.020 119.730 85.350 120.720 ;
        RECT 86.010 120.210 86.960 121.540 ;
      LAYER li1 ;
        RECT 86.050 119.580 86.940 119.970 ;
        RECT 87.140 119.730 87.390 121.790 ;
      LAYER li1 ;
        RECT 87.580 121.710 88.170 121.790 ;
        RECT 87.580 121.540 87.610 121.710 ;
        RECT 87.780 121.540 87.970 121.710 ;
        RECT 88.140 121.540 88.170 121.710 ;
        RECT 87.580 120.210 88.170 121.540 ;
        RECT 88.570 121.760 90.020 121.790 ;
        RECT 88.570 121.590 88.820 121.760 ;
        RECT 88.990 121.590 89.180 121.760 ;
        RECT 89.350 121.590 89.620 121.760 ;
        RECT 89.790 121.590 90.020 121.760 ;
        RECT 88.570 120.720 90.020 121.590 ;
        RECT 90.330 121.710 92.000 121.790 ;
        RECT 90.330 121.540 90.360 121.710 ;
        RECT 90.530 121.540 90.720 121.710 ;
        RECT 90.890 121.540 91.080 121.710 ;
        RECT 91.250 121.540 91.440 121.710 ;
        RECT 91.610 121.540 91.800 121.710 ;
        RECT 91.970 121.540 92.000 121.710 ;
      LAYER li1 ;
        RECT 87.140 119.560 87.720 119.730 ;
        RECT 87.500 119.380 87.720 119.560 ;
      LAYER li1 ;
        RECT 84.480 118.880 85.780 119.280 ;
        RECT 84.170 118.400 85.780 118.880 ;
        RECT 86.010 118.400 87.320 119.380 ;
      LAYER li1 ;
        RECT 87.500 119.210 88.100 119.380 ;
        RECT 87.770 119.040 88.100 119.210 ;
      LAYER li1 ;
        RECT 88.800 119.280 89.130 120.060 ;
        RECT 89.340 119.730 89.670 120.720 ;
        RECT 90.330 120.330 92.000 121.540 ;
      LAYER li1 ;
        RECT 90.370 119.810 91.560 120.150 ;
        RECT 91.740 119.810 92.070 120.150 ;
        RECT 92.260 119.630 92.520 121.790 ;
      LAYER li1 ;
        RECT 92.890 121.760 94.340 121.790 ;
        RECT 92.890 121.590 93.140 121.760 ;
        RECT 93.310 121.590 93.500 121.760 ;
        RECT 93.670 121.590 93.940 121.760 ;
        RECT 94.110 121.590 94.340 121.760 ;
        RECT 92.890 120.720 94.340 121.590 ;
        RECT 94.710 121.670 96.520 121.840 ;
      LAYER li1 ;
        RECT 91.440 119.460 92.520 119.630 ;
        RECT 87.770 118.870 88.160 119.040 ;
      LAYER li1 ;
        RECT 88.800 118.880 90.100 119.280 ;
      LAYER li1 ;
        RECT 87.770 118.550 88.100 118.870 ;
      LAYER li1 ;
        RECT 88.490 118.400 90.100 118.880 ;
        RECT 90.330 118.400 91.260 119.360 ;
      LAYER li1 ;
        RECT 91.440 118.530 91.770 119.460 ;
      LAYER li1 ;
        RECT 93.120 119.280 93.450 120.060 ;
        RECT 93.660 119.730 93.990 120.720 ;
        RECT 94.710 120.210 95.040 121.670 ;
      LAYER li1 ;
        RECT 95.490 120.210 95.850 121.490 ;
        RECT 94.690 119.540 95.400 119.870 ;
      LAYER li1 ;
        RECT 91.960 118.400 92.550 119.280 ;
        RECT 93.120 118.880 94.420 119.280 ;
        RECT 92.810 118.400 94.420 118.880 ;
        RECT 94.650 118.400 95.240 119.360 ;
      LAYER li1 ;
        RECT 95.650 119.010 95.850 120.210 ;
      LAYER li1 ;
        RECT 96.270 120.130 96.520 121.670 ;
        RECT 96.700 121.710 97.650 121.790 ;
        RECT 96.700 121.540 96.730 121.710 ;
        RECT 96.900 121.540 97.090 121.710 ;
        RECT 97.260 121.540 97.450 121.710 ;
        RECT 97.620 121.540 97.650 121.710 ;
        RECT 96.700 120.310 97.650 121.540 ;
        RECT 97.830 120.130 98.160 121.790 ;
        RECT 98.650 121.760 100.100 121.790 ;
        RECT 98.650 121.590 98.900 121.760 ;
        RECT 99.070 121.590 99.260 121.760 ;
        RECT 99.430 121.590 99.700 121.760 ;
        RECT 99.870 121.590 100.100 121.760 ;
        RECT 98.650 120.720 100.100 121.590 ;
        RECT 100.890 121.710 101.480 121.790 ;
        RECT 100.890 121.540 100.920 121.710 ;
        RECT 101.090 121.540 101.280 121.710 ;
        RECT 101.450 121.540 101.480 121.710 ;
        RECT 96.270 119.960 98.160 120.130 ;
      LAYER li1 ;
        RECT 96.030 119.540 96.360 119.780 ;
        RECT 96.610 119.540 97.320 119.780 ;
        RECT 97.500 119.540 98.280 119.780 ;
        RECT 96.270 119.010 96.520 119.360 ;
        RECT 95.650 118.840 96.520 119.010 ;
        RECT 96.270 118.530 96.520 118.840 ;
      LAYER li1 ;
        RECT 96.700 118.400 98.310 119.360 ;
        RECT 98.880 119.280 99.210 120.060 ;
        RECT 99.420 119.730 99.750 120.720 ;
        RECT 100.890 120.210 101.480 121.540 ;
      LAYER li1 ;
        RECT 101.760 120.210 102.150 121.790 ;
      LAYER li1 ;
        RECT 102.490 121.760 103.940 121.790 ;
        RECT 102.490 121.590 102.740 121.760 ;
        RECT 102.910 121.590 103.100 121.760 ;
        RECT 103.270 121.590 103.540 121.760 ;
        RECT 103.710 121.590 103.940 121.760 ;
        RECT 102.490 120.720 103.940 121.590 ;
        RECT 104.250 121.710 105.510 121.790 ;
        RECT 104.250 121.540 104.260 121.710 ;
        RECT 104.430 121.540 104.620 121.710 ;
        RECT 104.790 121.540 104.980 121.710 ;
        RECT 105.150 121.540 105.340 121.710 ;
      LAYER li1 ;
        RECT 100.930 119.580 101.640 119.970 ;
      LAYER li1 ;
        RECT 98.880 118.880 100.180 119.280 ;
        RECT 98.570 118.400 100.180 118.880 ;
        RECT 100.890 118.400 101.480 119.360 ;
      LAYER li1 ;
        RECT 101.820 118.530 102.150 120.210 ;
      LAYER li1 ;
        RECT 102.720 119.280 103.050 120.060 ;
        RECT 103.260 119.730 103.590 120.720 ;
        RECT 104.250 120.310 105.510 121.540 ;
      LAYER li1 ;
        RECT 106.040 121.290 106.210 121.790 ;
        RECT 105.690 120.210 106.210 121.290 ;
      LAYER li1 ;
        RECT 106.470 121.710 107.780 121.790 ;
        RECT 106.470 121.540 106.500 121.710 ;
        RECT 106.670 121.540 106.860 121.710 ;
        RECT 107.030 121.540 107.220 121.710 ;
        RECT 107.390 121.540 107.580 121.710 ;
        RECT 107.750 121.540 107.780 121.710 ;
        RECT 106.470 120.330 107.780 121.540 ;
        RECT 108.500 121.760 111.240 121.780 ;
        RECT 108.500 121.590 108.710 121.760 ;
        RECT 108.880 121.590 109.150 121.760 ;
        RECT 109.320 121.590 109.560 121.760 ;
        RECT 109.730 121.590 109.990 121.760 ;
        RECT 110.160 121.590 110.430 121.760 ;
        RECT 110.600 121.590 110.840 121.760 ;
        RECT 111.010 121.590 111.240 121.760 ;
        RECT 108.500 120.710 111.240 121.590 ;
        RECT 112.340 121.760 115.080 121.780 ;
        RECT 112.340 121.590 112.550 121.760 ;
        RECT 112.720 121.590 112.990 121.760 ;
        RECT 113.160 121.590 113.400 121.760 ;
        RECT 113.570 121.590 113.830 121.760 ;
        RECT 114.000 121.590 114.270 121.760 ;
        RECT 114.440 121.590 114.680 121.760 ;
        RECT 114.850 121.590 115.080 121.760 ;
        RECT 112.340 120.710 115.080 121.590 ;
        RECT 116.180 121.760 118.920 121.780 ;
        RECT 116.180 121.590 116.390 121.760 ;
        RECT 116.560 121.590 116.830 121.760 ;
        RECT 117.000 121.590 117.240 121.760 ;
        RECT 117.410 121.590 117.670 121.760 ;
        RECT 117.840 121.590 118.110 121.760 ;
        RECT 118.280 121.590 118.520 121.760 ;
        RECT 118.690 121.590 118.920 121.760 ;
        RECT 116.180 120.710 118.920 121.590 ;
        RECT 120.020 121.760 122.760 121.780 ;
        RECT 120.020 121.590 120.230 121.760 ;
        RECT 120.400 121.590 120.670 121.760 ;
        RECT 120.840 121.590 121.080 121.760 ;
        RECT 121.250 121.590 121.510 121.760 ;
        RECT 121.680 121.590 121.950 121.760 ;
        RECT 122.120 121.590 122.360 121.760 ;
        RECT 122.530 121.590 122.760 121.760 ;
        RECT 120.020 120.710 122.760 121.590 ;
        RECT 123.860 121.760 126.600 121.780 ;
        RECT 123.860 121.590 124.070 121.760 ;
        RECT 124.240 121.590 124.510 121.760 ;
        RECT 124.680 121.590 124.920 121.760 ;
        RECT 125.090 121.590 125.350 121.760 ;
        RECT 125.520 121.590 125.790 121.760 ;
        RECT 125.960 121.590 126.200 121.760 ;
        RECT 126.370 121.590 126.600 121.760 ;
        RECT 123.860 120.710 126.600 121.590 ;
        RECT 127.700 121.760 130.440 121.780 ;
        RECT 127.700 121.590 127.910 121.760 ;
        RECT 128.080 121.590 128.350 121.760 ;
        RECT 128.520 121.590 128.760 121.760 ;
        RECT 128.930 121.590 129.190 121.760 ;
        RECT 129.360 121.590 129.630 121.760 ;
        RECT 129.800 121.590 130.040 121.760 ;
        RECT 130.210 121.590 130.440 121.760 ;
        RECT 127.700 120.710 130.440 121.590 ;
        RECT 131.540 121.760 134.280 121.780 ;
        RECT 131.540 121.590 131.750 121.760 ;
        RECT 131.920 121.590 132.190 121.760 ;
        RECT 132.360 121.590 132.600 121.760 ;
        RECT 132.770 121.590 133.030 121.760 ;
        RECT 133.200 121.590 133.470 121.760 ;
        RECT 133.640 121.590 133.880 121.760 ;
        RECT 134.050 121.590 134.280 121.760 ;
        RECT 131.540 120.710 134.280 121.590 ;
        RECT 135.380 121.760 138.120 121.780 ;
        RECT 135.380 121.590 135.590 121.760 ;
        RECT 135.760 121.590 136.030 121.760 ;
        RECT 136.200 121.590 136.440 121.760 ;
        RECT 136.610 121.590 136.870 121.760 ;
        RECT 137.040 121.590 137.310 121.760 ;
        RECT 137.480 121.590 137.720 121.760 ;
        RECT 137.890 121.590 138.120 121.760 ;
        RECT 135.380 120.710 138.120 121.590 ;
        RECT 138.970 121.760 140.420 121.790 ;
        RECT 138.970 121.590 139.220 121.760 ;
        RECT 139.390 121.590 139.580 121.760 ;
        RECT 139.750 121.590 140.020 121.760 ;
        RECT 140.190 121.590 140.420 121.760 ;
        RECT 138.970 120.720 140.420 121.590 ;
      LAYER li1 ;
        RECT 105.690 120.130 105.960 120.210 ;
        RECT 104.900 119.960 105.960 120.130 ;
        RECT 104.290 119.570 104.710 119.900 ;
        RECT 104.900 119.390 105.070 119.960 ;
        RECT 106.410 119.840 106.920 120.150 ;
        RECT 107.170 119.840 107.880 120.150 ;
        RECT 105.250 119.570 105.760 119.780 ;
      LAYER li1 ;
        RECT 105.960 119.490 107.830 119.660 ;
        RECT 102.720 118.880 104.020 119.280 ;
        RECT 102.410 118.400 104.020 118.880 ;
        RECT 104.320 118.470 104.650 119.390 ;
      LAYER li1 ;
        RECT 104.900 118.650 105.430 119.390 ;
      LAYER li1 ;
        RECT 105.960 118.470 106.130 119.490 ;
        RECT 104.320 118.300 106.130 118.470 ;
        RECT 106.310 118.400 107.410 119.310 ;
        RECT 107.580 118.560 107.830 119.490 ;
        RECT 108.740 119.390 109.070 120.060 ;
        RECT 109.470 119.730 109.800 120.710 ;
        RECT 110.020 119.390 110.350 120.060 ;
        RECT 110.750 119.730 111.080 120.710 ;
        RECT 112.580 119.390 112.910 120.060 ;
        RECT 113.310 119.730 113.640 120.710 ;
        RECT 113.860 119.390 114.190 120.060 ;
        RECT 114.590 119.730 114.920 120.710 ;
        RECT 116.420 119.390 116.750 120.060 ;
        RECT 117.150 119.730 117.480 120.710 ;
        RECT 117.700 119.390 118.030 120.060 ;
        RECT 118.430 119.730 118.760 120.710 ;
        RECT 120.260 119.390 120.590 120.060 ;
        RECT 120.990 119.730 121.320 120.710 ;
        RECT 121.540 119.390 121.870 120.060 ;
        RECT 122.270 119.730 122.600 120.710 ;
        RECT 124.100 119.390 124.430 120.060 ;
        RECT 124.830 119.730 125.160 120.710 ;
        RECT 125.380 119.390 125.710 120.060 ;
        RECT 126.110 119.730 126.440 120.710 ;
        RECT 127.940 119.390 128.270 120.060 ;
        RECT 128.670 119.730 129.000 120.710 ;
        RECT 129.220 119.390 129.550 120.060 ;
        RECT 129.950 119.730 130.280 120.710 ;
        RECT 131.780 119.390 132.110 120.060 ;
        RECT 132.510 119.730 132.840 120.710 ;
        RECT 133.060 119.390 133.390 120.060 ;
        RECT 133.790 119.730 134.120 120.710 ;
        RECT 135.620 119.390 135.950 120.060 ;
        RECT 136.350 119.730 136.680 120.710 ;
        RECT 136.900 119.390 137.230 120.060 ;
        RECT 137.630 119.730 137.960 120.710 ;
        RECT 108.580 118.390 111.310 119.390 ;
        RECT 112.420 118.390 115.150 119.390 ;
        RECT 116.260 118.390 118.990 119.390 ;
        RECT 120.100 118.390 122.830 119.390 ;
        RECT 123.940 118.390 126.670 119.390 ;
        RECT 127.780 118.390 130.510 119.390 ;
        RECT 131.620 118.390 134.350 119.390 ;
        RECT 135.460 118.390 138.190 119.390 ;
        RECT 139.200 119.280 139.530 120.060 ;
        RECT 139.740 119.730 140.070 120.720 ;
        RECT 139.200 118.880 140.500 119.280 ;
        RECT 138.890 118.400 140.500 118.880 ;
        RECT 5.760 117.940 5.920 118.120 ;
        RECT 6.090 117.940 6.400 118.120 ;
        RECT 6.570 117.940 6.880 118.120 ;
        RECT 7.050 117.940 7.360 118.120 ;
        RECT 7.530 117.940 7.840 118.120 ;
        RECT 8.010 117.940 8.320 118.120 ;
        RECT 8.490 117.940 8.800 118.120 ;
        RECT 8.970 117.940 9.280 118.120 ;
        RECT 9.450 117.940 9.760 118.120 ;
        RECT 9.930 117.940 10.240 118.120 ;
        RECT 10.410 117.940 10.560 118.120 ;
        RECT 11.040 117.940 11.200 118.120 ;
        RECT 11.370 117.940 11.680 118.120 ;
        RECT 11.850 117.940 12.160 118.120 ;
        RECT 12.330 117.940 12.640 118.120 ;
        RECT 12.810 117.940 13.120 118.120 ;
        RECT 13.290 117.940 13.600 118.120 ;
        RECT 13.770 117.940 14.080 118.120 ;
        RECT 14.250 117.940 14.560 118.120 ;
        RECT 14.730 117.940 15.040 118.120 ;
        RECT 15.210 117.940 15.520 118.120 ;
        RECT 15.690 117.940 16.000 118.120 ;
        RECT 16.170 117.940 16.480 118.120 ;
        RECT 16.650 117.940 16.960 118.120 ;
        RECT 17.130 117.940 17.440 118.120 ;
        RECT 17.610 117.940 17.920 118.120 ;
        RECT 18.090 117.940 18.400 118.120 ;
        RECT 18.570 117.940 18.880 118.120 ;
        RECT 19.050 117.940 19.360 118.120 ;
        RECT 19.530 117.940 19.840 118.120 ;
        RECT 20.010 117.940 20.320 118.120 ;
        RECT 20.490 117.940 20.800 118.120 ;
        RECT 20.970 117.940 21.280 118.120 ;
        RECT 21.450 117.940 21.760 118.120 ;
        RECT 21.930 117.940 22.240 118.120 ;
        RECT 22.410 117.940 22.720 118.120 ;
        RECT 22.890 117.940 23.200 118.120 ;
        RECT 23.370 117.940 23.680 118.120 ;
        RECT 23.850 117.940 24.160 118.120 ;
        RECT 24.330 117.940 24.640 118.120 ;
        RECT 24.810 117.940 25.120 118.120 ;
        RECT 25.290 117.940 25.600 118.120 ;
        RECT 25.770 117.940 26.080 118.120 ;
        RECT 26.250 117.940 26.560 118.120 ;
        RECT 26.730 117.940 27.040 118.120 ;
        RECT 27.210 117.940 27.520 118.120 ;
        RECT 27.690 117.940 28.000 118.120 ;
        RECT 28.170 117.940 28.320 118.120 ;
        RECT 28.800 117.940 28.960 118.120 ;
        RECT 29.130 117.940 29.440 118.120 ;
        RECT 29.610 117.940 29.920 118.120 ;
        RECT 30.090 117.940 30.400 118.120 ;
        RECT 30.570 117.940 30.880 118.120 ;
        RECT 31.050 117.940 31.360 118.120 ;
        RECT 31.530 117.940 31.840 118.120 ;
        RECT 32.010 117.940 32.320 118.120 ;
        RECT 32.490 117.940 32.800 118.120 ;
        RECT 32.970 117.940 33.280 118.120 ;
        RECT 33.450 117.940 33.760 118.120 ;
        RECT 33.930 117.940 34.240 118.120 ;
        RECT 34.410 117.940 34.720 118.120 ;
        RECT 34.890 117.940 35.200 118.120 ;
        RECT 35.370 117.940 35.680 118.120 ;
        RECT 35.850 117.940 36.160 118.120 ;
        RECT 36.330 117.940 36.640 118.120 ;
        RECT 36.810 117.940 37.120 118.120 ;
        RECT 37.290 117.940 37.600 118.120 ;
        RECT 37.770 117.940 38.080 118.120 ;
        RECT 38.250 117.940 38.560 118.120 ;
        RECT 38.730 117.940 39.040 118.120 ;
        RECT 39.210 117.940 39.520 118.120 ;
        RECT 39.690 117.940 40.000 118.120 ;
        RECT 40.170 117.940 40.480 118.120 ;
        RECT 40.650 117.940 40.960 118.120 ;
        RECT 41.130 117.940 41.440 118.120 ;
        RECT 41.610 117.940 41.920 118.120 ;
        RECT 42.090 117.940 42.400 118.120 ;
        RECT 42.570 117.940 42.880 118.120 ;
        RECT 43.050 117.940 43.200 118.120 ;
        RECT 43.680 117.940 43.840 118.120 ;
        RECT 44.010 117.940 44.320 118.120 ;
        RECT 44.490 117.940 44.800 118.120 ;
        RECT 44.970 117.940 45.280 118.120 ;
        RECT 45.450 117.940 45.760 118.120 ;
        RECT 45.930 117.940 46.240 118.120 ;
        RECT 46.410 117.940 46.720 118.120 ;
        RECT 46.890 117.940 47.200 118.120 ;
        RECT 47.370 117.940 47.680 118.120 ;
        RECT 47.850 117.940 48.160 118.120 ;
        RECT 48.330 117.940 48.640 118.120 ;
        RECT 48.810 117.940 49.120 118.120 ;
        RECT 49.290 117.940 49.600 118.120 ;
        RECT 49.770 117.940 49.920 118.120 ;
        RECT 50.400 117.940 50.560 118.120 ;
        RECT 50.730 117.940 51.040 118.120 ;
        RECT 51.210 117.940 51.520 118.120 ;
        RECT 51.690 117.940 52.000 118.120 ;
        RECT 52.170 117.940 52.480 118.120 ;
        RECT 52.650 117.940 52.960 118.120 ;
        RECT 53.130 117.940 53.440 118.120 ;
        RECT 53.610 117.940 53.920 118.120 ;
        RECT 54.090 117.940 54.400 118.120 ;
        RECT 54.570 117.940 54.880 118.120 ;
        RECT 55.050 117.940 55.360 118.120 ;
        RECT 55.530 117.940 55.840 118.120 ;
        RECT 56.010 117.940 56.320 118.120 ;
        RECT 56.490 117.940 56.800 118.120 ;
        RECT 56.970 117.940 57.280 118.120 ;
        RECT 57.450 117.940 57.760 118.120 ;
        RECT 57.930 117.940 58.240 118.120 ;
        RECT 58.410 117.940 58.720 118.120 ;
        RECT 58.890 117.940 59.200 118.120 ;
        RECT 59.370 117.940 59.680 118.120 ;
        RECT 59.850 117.940 60.160 118.120 ;
        RECT 60.330 117.940 60.640 118.120 ;
        RECT 60.810 117.940 61.120 118.120 ;
        RECT 61.290 117.940 61.600 118.120 ;
        RECT 61.770 117.940 62.080 118.120 ;
        RECT 62.250 117.940 62.560 118.120 ;
        RECT 62.730 117.940 63.040 118.120 ;
        RECT 63.210 117.940 63.520 118.120 ;
        RECT 63.690 117.940 64.000 118.120 ;
        RECT 64.170 117.940 64.480 118.120 ;
        RECT 64.650 117.940 64.960 118.120 ;
        RECT 65.130 117.940 65.440 118.120 ;
        RECT 65.610 117.940 65.920 118.120 ;
        RECT 66.090 117.940 66.400 118.120 ;
        RECT 66.570 117.940 66.880 118.120 ;
        RECT 67.050 117.940 67.200 118.120 ;
        RECT 67.680 117.940 67.840 118.120 ;
        RECT 68.010 117.940 68.320 118.120 ;
        RECT 68.490 117.940 68.800 118.120 ;
        RECT 68.970 117.940 69.280 118.120 ;
        RECT 69.450 117.940 69.760 118.120 ;
        RECT 69.930 117.940 70.240 118.120 ;
        RECT 70.410 117.940 70.720 118.120 ;
        RECT 70.890 117.940 71.200 118.120 ;
        RECT 71.370 117.940 71.680 118.120 ;
        RECT 71.850 117.940 72.160 118.120 ;
        RECT 72.330 117.940 72.640 118.120 ;
        RECT 72.810 117.940 73.120 118.120 ;
        RECT 73.290 117.940 73.600 118.120 ;
        RECT 73.770 117.940 74.080 118.120 ;
        RECT 74.250 117.940 74.560 118.120 ;
        RECT 74.730 117.940 75.040 118.120 ;
        RECT 75.210 117.940 75.520 118.120 ;
        RECT 75.690 117.940 76.000 118.120 ;
        RECT 76.170 117.940 76.480 118.120 ;
        RECT 76.650 117.940 76.960 118.120 ;
        RECT 77.130 117.940 77.440 118.120 ;
        RECT 77.610 117.940 77.920 118.120 ;
        RECT 78.090 117.940 78.400 118.120 ;
        RECT 78.570 117.940 78.880 118.120 ;
        RECT 79.050 117.940 79.360 118.120 ;
        RECT 79.530 117.940 79.840 118.120 ;
        RECT 80.010 117.940 80.320 118.120 ;
        RECT 80.490 117.940 80.800 118.120 ;
        RECT 80.970 117.940 81.280 118.120 ;
        RECT 81.450 117.940 81.760 118.120 ;
        RECT 81.930 117.940 82.240 118.120 ;
        RECT 82.410 117.940 82.720 118.120 ;
        RECT 82.890 117.940 83.200 118.120 ;
        RECT 83.370 117.940 83.680 118.120 ;
        RECT 83.850 117.940 84.160 118.120 ;
        RECT 84.330 117.940 84.640 118.120 ;
        RECT 84.810 117.940 85.120 118.120 ;
        RECT 85.290 117.940 85.600 118.120 ;
        RECT 85.770 117.940 86.080 118.120 ;
        RECT 86.250 117.940 86.560 118.120 ;
        RECT 86.730 117.940 87.040 118.120 ;
        RECT 87.210 117.940 87.520 118.120 ;
        RECT 87.690 117.940 88.000 118.120 ;
        RECT 88.170 117.940 88.480 118.120 ;
        RECT 88.650 117.940 88.960 118.120 ;
        RECT 89.130 117.940 89.440 118.120 ;
        RECT 89.610 117.940 89.920 118.120 ;
        RECT 90.090 117.940 90.400 118.120 ;
        RECT 90.570 117.940 90.880 118.120 ;
        RECT 91.050 117.940 91.360 118.120 ;
        RECT 91.530 117.940 91.840 118.120 ;
        RECT 92.010 117.940 92.320 118.120 ;
        RECT 92.490 117.940 92.800 118.120 ;
        RECT 92.970 117.940 93.280 118.120 ;
        RECT 93.450 117.940 93.760 118.120 ;
        RECT 93.930 117.940 94.240 118.120 ;
        RECT 94.410 117.940 94.720 118.120 ;
        RECT 94.890 117.940 95.200 118.120 ;
        RECT 95.370 117.940 95.680 118.120 ;
        RECT 95.850 117.940 96.160 118.120 ;
        RECT 96.330 117.940 96.640 118.120 ;
        RECT 96.810 117.940 97.120 118.120 ;
        RECT 97.290 117.940 97.600 118.120 ;
        RECT 97.770 117.940 98.080 118.120 ;
        RECT 98.250 117.940 98.560 118.120 ;
        RECT 98.730 117.940 99.040 118.120 ;
        RECT 99.210 117.940 99.520 118.120 ;
        RECT 99.690 117.940 100.000 118.120 ;
        RECT 100.170 117.940 100.320 118.120 ;
        RECT 100.800 117.940 100.960 118.120 ;
        RECT 101.130 117.940 101.440 118.120 ;
        RECT 101.610 117.940 101.920 118.120 ;
        RECT 102.090 117.940 102.400 118.120 ;
        RECT 102.570 117.940 102.880 118.120 ;
        RECT 103.050 117.940 103.360 118.120 ;
        RECT 103.530 117.940 103.840 118.120 ;
        RECT 104.010 117.940 104.320 118.120 ;
        RECT 104.490 117.940 104.800 118.120 ;
        RECT 104.970 117.940 105.280 118.120 ;
        RECT 105.450 117.940 105.760 118.120 ;
        RECT 105.930 117.940 106.240 118.120 ;
        RECT 106.410 117.940 106.720 118.120 ;
        RECT 106.890 117.940 107.200 118.120 ;
        RECT 107.370 117.940 107.680 118.120 ;
        RECT 107.850 117.940 108.160 118.120 ;
        RECT 108.330 117.940 108.640 118.120 ;
        RECT 108.810 117.940 109.120 118.120 ;
        RECT 109.290 117.940 109.600 118.120 ;
        RECT 109.770 117.940 110.080 118.120 ;
        RECT 110.250 117.940 110.560 118.120 ;
        RECT 110.730 117.940 111.040 118.120 ;
        RECT 111.210 117.940 111.520 118.120 ;
        RECT 111.690 117.940 112.000 118.120 ;
        RECT 112.170 117.940 112.480 118.120 ;
        RECT 112.650 117.940 112.960 118.120 ;
        RECT 113.130 117.940 113.440 118.120 ;
        RECT 113.610 117.940 113.920 118.120 ;
        RECT 114.090 117.940 114.400 118.120 ;
        RECT 114.570 117.940 114.880 118.120 ;
        RECT 115.050 117.940 115.360 118.120 ;
        RECT 115.530 117.940 115.840 118.120 ;
        RECT 116.010 117.940 116.320 118.120 ;
        RECT 116.490 117.940 116.800 118.120 ;
        RECT 116.970 117.940 117.280 118.120 ;
        RECT 117.450 117.940 117.760 118.120 ;
        RECT 117.930 117.940 118.240 118.120 ;
        RECT 118.410 117.940 118.720 118.120 ;
        RECT 118.890 117.940 119.200 118.120 ;
        RECT 119.370 117.940 119.680 118.120 ;
        RECT 119.850 117.940 120.160 118.120 ;
        RECT 120.330 117.940 120.640 118.120 ;
        RECT 120.810 117.940 121.120 118.120 ;
        RECT 121.290 117.940 121.600 118.120 ;
        RECT 121.770 117.940 122.080 118.120 ;
        RECT 122.250 117.940 122.560 118.120 ;
        RECT 122.730 117.940 123.040 118.120 ;
        RECT 123.210 117.940 123.520 118.120 ;
        RECT 123.690 117.940 124.000 118.120 ;
        RECT 124.170 117.940 124.480 118.120 ;
        RECT 124.650 117.940 124.960 118.120 ;
        RECT 125.130 117.940 125.440 118.120 ;
        RECT 125.610 117.940 125.920 118.120 ;
        RECT 126.090 117.940 126.400 118.120 ;
        RECT 126.570 117.940 126.880 118.120 ;
        RECT 127.050 117.940 127.360 118.120 ;
        RECT 127.530 117.940 127.840 118.120 ;
        RECT 128.010 117.940 128.320 118.120 ;
        RECT 128.490 117.940 128.800 118.120 ;
        RECT 128.970 117.940 129.280 118.120 ;
        RECT 129.450 117.940 129.760 118.120 ;
        RECT 129.930 117.940 130.240 118.120 ;
        RECT 130.410 117.940 130.720 118.120 ;
        RECT 130.890 117.940 131.200 118.120 ;
        RECT 131.370 117.940 131.680 118.120 ;
        RECT 131.850 117.940 132.160 118.120 ;
        RECT 132.330 117.940 132.640 118.120 ;
        RECT 132.810 117.940 133.120 118.120 ;
        RECT 133.290 117.940 133.600 118.120 ;
        RECT 133.770 117.940 134.080 118.120 ;
        RECT 134.250 117.940 134.560 118.120 ;
        RECT 134.730 117.940 135.040 118.120 ;
        RECT 135.210 117.940 135.520 118.120 ;
        RECT 135.690 117.940 136.000 118.120 ;
        RECT 136.170 117.940 136.480 118.120 ;
        RECT 136.650 117.940 136.960 118.120 ;
        RECT 137.130 117.940 137.440 118.120 ;
        RECT 137.610 117.940 137.920 118.120 ;
        RECT 138.090 117.940 138.400 118.120 ;
        RECT 138.570 117.940 138.880 118.120 ;
        RECT 139.050 117.940 139.360 118.120 ;
        RECT 139.530 117.940 139.840 118.120 ;
        RECT 140.010 117.940 140.320 118.120 ;
        RECT 140.490 117.940 140.800 118.120 ;
        RECT 140.970 117.940 141.280 118.120 ;
        RECT 141.450 117.940 141.600 118.120 ;
        RECT 6.340 117.640 9.070 117.670 ;
        RECT 6.340 117.470 6.510 117.640 ;
        RECT 6.680 117.470 6.950 117.640 ;
        RECT 7.120 117.470 7.360 117.640 ;
        RECT 7.530 117.470 7.790 117.640 ;
        RECT 7.960 117.470 8.230 117.640 ;
        RECT 8.400 117.470 8.640 117.640 ;
        RECT 8.810 117.470 9.070 117.640 ;
        RECT 6.340 116.670 9.070 117.470 ;
        RECT 10.180 117.640 12.910 117.670 ;
        RECT 10.180 117.470 10.350 117.640 ;
        RECT 10.520 117.470 10.790 117.640 ;
        RECT 10.960 117.470 11.200 117.640 ;
        RECT 11.370 117.470 11.630 117.640 ;
        RECT 11.800 117.470 12.070 117.640 ;
        RECT 12.240 117.470 12.480 117.640 ;
        RECT 12.650 117.470 12.910 117.640 ;
        RECT 14.470 117.630 15.720 117.660 ;
        RECT 16.900 117.640 19.630 117.670 ;
        RECT 10.180 116.670 12.910 117.470 ;
        RECT 6.500 116.000 6.830 116.670 ;
        RECT 7.230 115.350 7.560 116.330 ;
        RECT 7.780 116.000 8.110 116.670 ;
        RECT 8.510 115.350 8.840 116.330 ;
        RECT 10.340 116.000 10.670 116.670 ;
        RECT 11.070 115.350 11.400 116.330 ;
        RECT 11.620 116.000 11.950 116.670 ;
        RECT 12.350 115.350 12.680 116.330 ;
      LAYER li1 ;
        RECT 14.040 115.850 14.290 117.530 ;
      LAYER li1 ;
        RECT 14.640 117.460 14.830 117.630 ;
        RECT 15.000 117.460 15.190 117.630 ;
        RECT 15.360 117.460 15.550 117.630 ;
        RECT 14.470 117.090 15.720 117.460 ;
        RECT 15.900 116.910 16.150 117.530 ;
        RECT 14.600 116.740 16.150 116.910 ;
        RECT 14.600 116.280 14.930 116.740 ;
        RECT 6.260 114.470 9.000 115.350 ;
        RECT 6.260 114.300 6.470 114.470 ;
        RECT 6.640 114.300 6.910 114.470 ;
        RECT 7.080 114.300 7.320 114.470 ;
        RECT 7.490 114.300 7.750 114.470 ;
        RECT 7.920 114.300 8.190 114.470 ;
        RECT 8.360 114.300 8.600 114.470 ;
        RECT 8.770 114.300 9.000 114.470 ;
        RECT 6.260 114.280 9.000 114.300 ;
        RECT 10.100 114.470 12.840 115.350 ;
        RECT 10.100 114.300 10.310 114.470 ;
        RECT 10.480 114.300 10.750 114.470 ;
        RECT 10.920 114.300 11.160 114.470 ;
        RECT 11.330 114.300 11.590 114.470 ;
        RECT 11.760 114.300 12.030 114.470 ;
        RECT 12.200 114.300 12.440 114.470 ;
        RECT 12.610 114.300 12.840 114.470 ;
        RECT 10.100 114.280 12.840 114.300 ;
      LAYER li1 ;
        RECT 14.040 114.270 14.470 115.850 ;
      LAYER li1 ;
        RECT 14.650 114.520 15.210 115.850 ;
      LAYER li1 ;
        RECT 15.390 114.770 15.720 116.560 ;
      LAYER li1 ;
        RECT 15.900 115.020 16.150 116.740 ;
        RECT 16.900 117.470 17.070 117.640 ;
        RECT 17.240 117.470 17.510 117.640 ;
        RECT 17.680 117.470 17.920 117.640 ;
        RECT 18.090 117.470 18.350 117.640 ;
        RECT 18.520 117.470 18.790 117.640 ;
        RECT 18.960 117.470 19.200 117.640 ;
        RECT 19.370 117.470 19.630 117.640 ;
        RECT 16.900 116.670 19.630 117.470 ;
        RECT 20.740 117.640 23.470 117.670 ;
        RECT 20.740 117.470 20.910 117.640 ;
        RECT 21.080 117.470 21.350 117.640 ;
        RECT 21.520 117.470 21.760 117.640 ;
        RECT 21.930 117.470 22.190 117.640 ;
        RECT 22.360 117.470 22.630 117.640 ;
        RECT 22.800 117.470 23.040 117.640 ;
        RECT 23.210 117.470 23.470 117.640 ;
        RECT 20.740 116.670 23.470 117.470 ;
        RECT 25.050 117.630 25.640 117.660 ;
        RECT 25.050 117.460 25.080 117.630 ;
        RECT 25.250 117.460 25.440 117.630 ;
        RECT 25.610 117.460 25.640 117.630 ;
        RECT 26.980 117.640 29.710 117.670 ;
        RECT 25.050 116.700 25.640 117.460 ;
        RECT 17.060 116.000 17.390 116.670 ;
        RECT 17.790 115.350 18.120 116.330 ;
        RECT 18.340 116.000 18.670 116.670 ;
        RECT 19.070 115.350 19.400 116.330 ;
        RECT 20.900 116.000 21.230 116.670 ;
        RECT 21.630 115.350 21.960 116.330 ;
        RECT 22.180 116.000 22.510 116.670 ;
        RECT 22.910 115.350 23.240 116.330 ;
      LAYER li1 ;
        RECT 25.090 116.090 25.800 116.480 ;
        RECT 25.980 115.850 26.310 117.530 ;
      LAYER li1 ;
        RECT 26.980 117.470 27.150 117.640 ;
        RECT 27.320 117.470 27.590 117.640 ;
        RECT 27.760 117.470 28.000 117.640 ;
        RECT 28.170 117.470 28.430 117.640 ;
        RECT 28.600 117.470 28.870 117.640 ;
        RECT 29.040 117.470 29.280 117.640 ;
        RECT 29.450 117.470 29.710 117.640 ;
        RECT 26.980 116.670 29.710 117.470 ;
        RECT 30.820 117.640 33.550 117.670 ;
        RECT 30.820 117.470 30.990 117.640 ;
        RECT 31.160 117.470 31.430 117.640 ;
        RECT 31.600 117.470 31.840 117.640 ;
        RECT 32.010 117.470 32.270 117.640 ;
        RECT 32.440 117.470 32.710 117.640 ;
        RECT 32.880 117.470 33.120 117.640 ;
        RECT 33.290 117.470 33.550 117.640 ;
        RECT 30.820 116.670 33.550 117.470 ;
        RECT 34.660 117.640 37.390 117.670 ;
        RECT 34.660 117.470 34.830 117.640 ;
        RECT 35.000 117.470 35.270 117.640 ;
        RECT 35.440 117.470 35.680 117.640 ;
        RECT 35.850 117.470 36.110 117.640 ;
        RECT 36.280 117.470 36.550 117.640 ;
        RECT 36.720 117.470 36.960 117.640 ;
        RECT 37.130 117.470 37.390 117.640 ;
        RECT 34.660 116.670 37.390 117.470 ;
        RECT 38.500 117.640 41.230 117.670 ;
        RECT 38.500 117.470 38.670 117.640 ;
        RECT 38.840 117.470 39.110 117.640 ;
        RECT 39.280 117.470 39.520 117.640 ;
        RECT 39.690 117.470 39.950 117.640 ;
        RECT 40.120 117.470 40.390 117.640 ;
        RECT 40.560 117.470 40.800 117.640 ;
        RECT 40.970 117.470 41.230 117.640 ;
        RECT 38.500 116.670 41.230 117.470 ;
        RECT 42.880 117.590 44.690 117.760 ;
        RECT 42.880 116.670 43.210 117.590 ;
      LAYER li1 ;
        RECT 43.460 116.670 43.990 117.410 ;
      LAYER li1 ;
        RECT 27.140 116.000 27.470 116.670 ;
        RECT 14.650 114.350 14.660 114.520 ;
        RECT 14.830 114.350 15.020 114.520 ;
        RECT 15.190 114.350 15.210 114.520 ;
        RECT 14.650 114.270 15.210 114.350 ;
        RECT 16.820 114.470 19.560 115.350 ;
        RECT 16.820 114.300 17.030 114.470 ;
        RECT 17.200 114.300 17.470 114.470 ;
        RECT 17.640 114.300 17.880 114.470 ;
        RECT 18.050 114.300 18.310 114.470 ;
        RECT 18.480 114.300 18.750 114.470 ;
        RECT 18.920 114.300 19.160 114.470 ;
        RECT 19.330 114.300 19.560 114.470 ;
        RECT 16.820 114.280 19.560 114.300 ;
        RECT 20.660 114.470 23.400 115.350 ;
        RECT 20.660 114.300 20.870 114.470 ;
        RECT 21.040 114.300 21.310 114.470 ;
        RECT 21.480 114.300 21.720 114.470 ;
        RECT 21.890 114.300 22.150 114.470 ;
        RECT 22.320 114.300 22.590 114.470 ;
        RECT 22.760 114.300 23.000 114.470 ;
        RECT 23.170 114.300 23.400 114.470 ;
        RECT 20.660 114.280 23.400 114.300 ;
        RECT 25.050 114.520 25.640 115.850 ;
        RECT 25.050 114.350 25.080 114.520 ;
        RECT 25.250 114.350 25.440 114.520 ;
        RECT 25.610 114.350 25.640 114.520 ;
        RECT 25.050 114.270 25.640 114.350 ;
      LAYER li1 ;
        RECT 25.920 114.270 26.310 115.850 ;
      LAYER li1 ;
        RECT 27.870 115.350 28.200 116.330 ;
        RECT 28.420 116.000 28.750 116.670 ;
        RECT 29.150 115.350 29.480 116.330 ;
        RECT 30.980 116.000 31.310 116.670 ;
        RECT 31.710 115.350 32.040 116.330 ;
        RECT 32.260 116.000 32.590 116.670 ;
        RECT 32.990 115.350 33.320 116.330 ;
        RECT 34.820 116.000 35.150 116.670 ;
        RECT 35.550 115.350 35.880 116.330 ;
        RECT 36.100 116.000 36.430 116.670 ;
        RECT 36.830 115.350 37.160 116.330 ;
        RECT 38.660 116.000 38.990 116.670 ;
        RECT 39.390 115.350 39.720 116.330 ;
        RECT 39.940 116.000 40.270 116.670 ;
        RECT 40.670 115.350 41.000 116.330 ;
      LAYER li1 ;
        RECT 42.850 116.160 43.270 116.490 ;
        RECT 43.460 116.100 43.630 116.670 ;
      LAYER li1 ;
        RECT 44.520 116.570 44.690 117.590 ;
        RECT 44.870 117.630 45.970 117.660 ;
        RECT 44.870 117.460 44.920 117.630 ;
        RECT 45.090 117.460 45.280 117.630 ;
        RECT 45.450 117.460 45.640 117.630 ;
        RECT 45.810 117.460 45.970 117.630 ;
        RECT 46.730 117.630 48.340 117.660 ;
        RECT 44.870 116.750 45.970 117.460 ;
        RECT 46.140 116.570 46.390 117.500 ;
        RECT 46.730 117.460 46.780 117.630 ;
        RECT 46.950 117.460 47.220 117.630 ;
        RECT 47.390 117.460 47.660 117.630 ;
        RECT 47.830 117.460 48.070 117.630 ;
        RECT 48.240 117.460 48.340 117.630 ;
        RECT 46.730 117.180 48.340 117.460 ;
      LAYER li1 ;
        RECT 43.810 116.280 44.320 116.490 ;
      LAYER li1 ;
        RECT 44.520 116.400 46.390 116.570 ;
        RECT 47.040 116.780 48.340 117.180 ;
        RECT 48.570 117.630 49.520 117.660 ;
        RECT 48.570 117.460 48.600 117.630 ;
        RECT 48.770 117.460 48.960 117.630 ;
        RECT 49.130 117.460 49.320 117.630 ;
        RECT 49.490 117.460 49.520 117.630 ;
        RECT 50.130 117.630 51.080 117.660 ;
      LAYER li1 ;
        RECT 43.460 115.930 44.520 116.100 ;
        RECT 44.250 115.850 44.520 115.930 ;
        RECT 44.970 115.910 45.480 116.220 ;
        RECT 45.730 115.910 46.440 116.220 ;
      LAYER li1 ;
        RECT 47.040 116.000 47.370 116.780 ;
        RECT 48.570 116.700 49.520 117.460 ;
      LAYER li1 ;
        RECT 49.700 116.820 49.950 117.530 ;
      LAYER li1 ;
        RECT 50.130 117.460 50.160 117.630 ;
        RECT 50.330 117.460 50.520 117.630 ;
        RECT 50.690 117.460 50.880 117.630 ;
        RECT 51.050 117.460 51.080 117.630 ;
        RECT 51.690 117.630 52.640 117.660 ;
        RECT 50.130 117.000 51.080 117.460 ;
      LAYER li1 ;
        RECT 51.260 116.820 51.510 117.530 ;
        RECT 49.700 116.650 51.510 116.820 ;
      LAYER li1 ;
        RECT 51.690 117.460 51.720 117.630 ;
        RECT 51.890 117.460 52.080 117.630 ;
        RECT 52.250 117.460 52.440 117.630 ;
        RECT 52.610 117.460 52.640 117.630 ;
        RECT 53.450 117.630 55.060 117.660 ;
        RECT 56.710 117.630 57.960 117.660 ;
        RECT 58.730 117.630 60.340 117.660 ;
        RECT 61.030 117.630 62.280 117.660 ;
        RECT 63.460 117.640 66.190 117.670 ;
        RECT 51.690 116.780 52.640 117.460 ;
      LAYER li1 ;
        RECT 49.700 116.480 49.870 116.650 ;
      LAYER li1 ;
        RECT 52.820 116.600 53.150 117.530 ;
        RECT 53.450 117.460 53.500 117.630 ;
        RECT 53.670 117.460 53.940 117.630 ;
        RECT 54.110 117.460 54.380 117.630 ;
        RECT 54.550 117.460 54.790 117.630 ;
        RECT 54.960 117.460 55.060 117.630 ;
        RECT 53.450 117.180 55.060 117.460 ;
        RECT 26.900 114.470 29.640 115.350 ;
        RECT 26.900 114.300 27.110 114.470 ;
        RECT 27.280 114.300 27.550 114.470 ;
        RECT 27.720 114.300 27.960 114.470 ;
        RECT 28.130 114.300 28.390 114.470 ;
        RECT 28.560 114.300 28.830 114.470 ;
        RECT 29.000 114.300 29.240 114.470 ;
        RECT 29.410 114.300 29.640 114.470 ;
        RECT 26.900 114.280 29.640 114.300 ;
        RECT 30.740 114.470 33.480 115.350 ;
        RECT 30.740 114.300 30.950 114.470 ;
        RECT 31.120 114.300 31.390 114.470 ;
        RECT 31.560 114.300 31.800 114.470 ;
        RECT 31.970 114.300 32.230 114.470 ;
        RECT 32.400 114.300 32.670 114.470 ;
        RECT 32.840 114.300 33.080 114.470 ;
        RECT 33.250 114.300 33.480 114.470 ;
        RECT 30.740 114.280 33.480 114.300 ;
        RECT 34.580 114.470 37.320 115.350 ;
        RECT 34.580 114.300 34.790 114.470 ;
        RECT 34.960 114.300 35.230 114.470 ;
        RECT 35.400 114.300 35.640 114.470 ;
        RECT 35.810 114.300 36.070 114.470 ;
        RECT 36.240 114.300 36.510 114.470 ;
        RECT 36.680 114.300 36.920 114.470 ;
        RECT 37.090 114.300 37.320 114.470 ;
        RECT 34.580 114.280 37.320 114.300 ;
        RECT 38.420 114.470 41.160 115.350 ;
        RECT 38.420 114.300 38.630 114.470 ;
        RECT 38.800 114.300 39.070 114.470 ;
        RECT 39.240 114.300 39.480 114.470 ;
        RECT 39.650 114.300 39.910 114.470 ;
        RECT 40.080 114.300 40.350 114.470 ;
        RECT 40.520 114.300 40.760 114.470 ;
        RECT 40.930 114.300 41.160 114.470 ;
        RECT 38.420 114.280 41.160 114.300 ;
        RECT 42.810 114.520 44.070 115.750 ;
      LAYER li1 ;
        RECT 44.250 114.770 44.770 115.850 ;
      LAYER li1 ;
        RECT 42.810 114.350 42.820 114.520 ;
        RECT 42.990 114.350 43.180 114.520 ;
        RECT 43.350 114.350 43.540 114.520 ;
        RECT 43.710 114.350 43.900 114.520 ;
        RECT 42.810 114.270 44.070 114.350 ;
      LAYER li1 ;
        RECT 44.600 114.270 44.770 114.770 ;
      LAYER li1 ;
        RECT 45.030 114.520 46.340 115.730 ;
        RECT 47.580 115.340 47.910 116.330 ;
      LAYER li1 ;
        RECT 48.610 116.250 49.870 116.480 ;
      LAYER li1 ;
        RECT 51.910 116.470 53.150 116.600 ;
        RECT 50.050 116.430 53.150 116.470 ;
        RECT 50.050 116.300 52.080 116.430 ;
      LAYER li1 ;
        RECT 49.700 116.120 49.870 116.250 ;
        RECT 49.700 115.950 51.590 116.120 ;
      LAYER li1 ;
        RECT 45.030 114.350 45.060 114.520 ;
        RECT 45.230 114.350 45.420 114.520 ;
        RECT 45.590 114.350 45.780 114.520 ;
        RECT 45.950 114.350 46.140 114.520 ;
        RECT 46.310 114.350 46.340 114.520 ;
        RECT 45.030 114.270 46.340 114.350 ;
        RECT 46.810 114.470 48.260 115.340 ;
        RECT 46.810 114.300 47.060 114.470 ;
        RECT 47.230 114.300 47.420 114.470 ;
        RECT 47.590 114.300 47.860 114.470 ;
        RECT 48.030 114.300 48.260 114.470 ;
        RECT 46.810 114.270 48.260 114.300 ;
        RECT 48.570 114.520 49.520 115.850 ;
        RECT 48.570 114.350 48.600 114.520 ;
        RECT 48.770 114.350 48.960 114.520 ;
        RECT 49.130 114.350 49.320 114.520 ;
        RECT 49.490 114.350 49.520 114.520 ;
        RECT 48.570 114.270 49.520 114.350 ;
      LAYER li1 ;
        RECT 49.700 114.270 49.950 115.950 ;
      LAYER li1 ;
        RECT 50.130 114.520 51.080 115.770 ;
        RECT 50.130 114.350 50.160 114.520 ;
        RECT 50.330 114.350 50.520 114.520 ;
        RECT 50.690 114.350 50.880 114.520 ;
        RECT 51.050 114.350 51.080 114.520 ;
        RECT 50.130 114.270 51.080 114.350 ;
      LAYER li1 ;
        RECT 51.260 114.270 51.590 115.950 ;
        RECT 52.370 115.910 52.700 116.250 ;
      LAYER li1 ;
        RECT 51.770 114.520 52.720 115.730 ;
        RECT 51.770 114.350 51.800 114.520 ;
        RECT 51.970 114.350 52.160 114.520 ;
        RECT 52.330 114.350 52.520 114.520 ;
        RECT 52.690 114.350 52.720 114.520 ;
        RECT 51.770 114.270 52.720 114.350 ;
        RECT 52.900 114.270 53.150 116.430 ;
        RECT 53.760 116.780 55.060 117.180 ;
        RECT 53.760 116.000 54.090 116.780 ;
        RECT 54.300 115.340 54.630 116.330 ;
      LAYER li1 ;
        RECT 56.280 115.850 56.530 117.530 ;
      LAYER li1 ;
        RECT 56.880 117.460 57.070 117.630 ;
        RECT 57.240 117.460 57.430 117.630 ;
        RECT 57.600 117.460 57.790 117.630 ;
        RECT 56.710 117.090 57.960 117.460 ;
        RECT 58.140 116.910 58.390 117.530 ;
        RECT 58.730 117.460 58.780 117.630 ;
        RECT 58.950 117.460 59.220 117.630 ;
        RECT 59.390 117.460 59.660 117.630 ;
        RECT 59.830 117.460 60.070 117.630 ;
        RECT 60.240 117.460 60.340 117.630 ;
        RECT 58.730 117.180 60.340 117.460 ;
        RECT 56.840 116.740 58.390 116.910 ;
        RECT 56.840 116.280 57.170 116.740 ;
        RECT 53.530 114.470 54.980 115.340 ;
        RECT 53.530 114.300 53.780 114.470 ;
        RECT 53.950 114.300 54.140 114.470 ;
        RECT 54.310 114.300 54.580 114.470 ;
        RECT 54.750 114.300 54.980 114.470 ;
        RECT 53.530 114.270 54.980 114.300 ;
      LAYER li1 ;
        RECT 56.280 114.270 56.710 115.850 ;
      LAYER li1 ;
        RECT 56.890 114.520 57.450 115.850 ;
      LAYER li1 ;
        RECT 57.630 114.770 57.960 116.560 ;
      LAYER li1 ;
        RECT 58.140 115.020 58.390 116.740 ;
        RECT 59.040 116.780 60.340 117.180 ;
        RECT 59.040 116.000 59.370 116.780 ;
        RECT 59.580 115.340 59.910 116.330 ;
      LAYER li1 ;
        RECT 60.600 115.850 60.850 117.530 ;
      LAYER li1 ;
        RECT 61.200 117.460 61.390 117.630 ;
        RECT 61.560 117.460 61.750 117.630 ;
        RECT 61.920 117.460 62.110 117.630 ;
        RECT 61.030 117.090 62.280 117.460 ;
        RECT 62.460 116.910 62.710 117.530 ;
        RECT 61.160 116.740 62.710 116.910 ;
        RECT 61.160 116.280 61.490 116.740 ;
        RECT 56.890 114.350 56.900 114.520 ;
        RECT 57.070 114.350 57.260 114.520 ;
        RECT 57.430 114.350 57.450 114.520 ;
        RECT 56.890 114.270 57.450 114.350 ;
        RECT 58.810 114.470 60.260 115.340 ;
        RECT 58.810 114.300 59.060 114.470 ;
        RECT 59.230 114.300 59.420 114.470 ;
        RECT 59.590 114.300 59.860 114.470 ;
        RECT 60.030 114.300 60.260 114.470 ;
        RECT 58.810 114.270 60.260 114.300 ;
      LAYER li1 ;
        RECT 60.600 114.270 61.030 115.850 ;
      LAYER li1 ;
        RECT 61.210 114.520 61.770 115.850 ;
      LAYER li1 ;
        RECT 61.950 114.770 62.280 116.560 ;
      LAYER li1 ;
        RECT 62.460 115.020 62.710 116.740 ;
        RECT 63.460 117.470 63.630 117.640 ;
        RECT 63.800 117.470 64.070 117.640 ;
        RECT 64.240 117.470 64.480 117.640 ;
        RECT 64.650 117.470 64.910 117.640 ;
        RECT 65.080 117.470 65.350 117.640 ;
        RECT 65.520 117.470 65.760 117.640 ;
        RECT 65.930 117.470 66.190 117.640 ;
        RECT 67.270 117.630 68.520 117.660 ;
        RECT 69.290 117.630 70.900 117.660 ;
        RECT 63.460 116.670 66.190 117.470 ;
        RECT 63.620 116.000 63.950 116.670 ;
        RECT 64.350 115.350 64.680 116.330 ;
        RECT 64.900 116.000 65.230 116.670 ;
        RECT 65.630 115.350 65.960 116.330 ;
      LAYER li1 ;
        RECT 66.840 115.850 67.090 117.530 ;
      LAYER li1 ;
        RECT 67.440 117.460 67.630 117.630 ;
        RECT 67.800 117.460 67.990 117.630 ;
        RECT 68.160 117.460 68.350 117.630 ;
        RECT 67.270 117.090 68.520 117.460 ;
        RECT 68.700 116.910 68.950 117.530 ;
        RECT 69.290 117.460 69.340 117.630 ;
        RECT 69.510 117.460 69.780 117.630 ;
        RECT 69.950 117.460 70.220 117.630 ;
        RECT 70.390 117.460 70.630 117.630 ;
        RECT 70.800 117.460 70.900 117.630 ;
        RECT 71.600 117.630 72.550 117.660 ;
        RECT 69.290 117.180 70.900 117.460 ;
        RECT 67.400 116.740 68.950 116.910 ;
        RECT 67.400 116.280 67.730 116.740 ;
        RECT 61.210 114.350 61.220 114.520 ;
        RECT 61.390 114.350 61.580 114.520 ;
        RECT 61.750 114.350 61.770 114.520 ;
        RECT 61.210 114.270 61.770 114.350 ;
        RECT 63.380 114.470 66.120 115.350 ;
        RECT 63.380 114.300 63.590 114.470 ;
        RECT 63.760 114.300 64.030 114.470 ;
        RECT 64.200 114.300 64.440 114.470 ;
        RECT 64.610 114.300 64.870 114.470 ;
        RECT 65.040 114.300 65.310 114.470 ;
        RECT 65.480 114.300 65.720 114.470 ;
        RECT 65.890 114.300 66.120 114.470 ;
        RECT 63.380 114.280 66.120 114.300 ;
      LAYER li1 ;
        RECT 66.840 114.270 67.270 115.850 ;
      LAYER li1 ;
        RECT 67.450 114.520 68.010 115.850 ;
      LAYER li1 ;
        RECT 68.190 114.770 68.520 116.560 ;
      LAYER li1 ;
        RECT 68.700 115.020 68.950 116.740 ;
        RECT 69.600 116.780 70.900 117.180 ;
        RECT 69.600 116.000 69.930 116.780 ;
        RECT 70.140 115.340 70.470 116.330 ;
        RECT 71.150 115.670 71.420 117.530 ;
        RECT 71.600 117.460 71.630 117.630 ;
        RECT 71.800 117.460 71.990 117.630 ;
        RECT 72.160 117.460 72.350 117.630 ;
        RECT 72.520 117.460 72.550 117.630 ;
        RECT 73.240 117.630 73.830 117.660 ;
        RECT 71.600 117.030 72.550 117.460 ;
        RECT 72.730 117.030 73.060 117.530 ;
      LAYER li1 ;
        RECT 71.600 115.880 71.930 116.850 ;
      LAYER li1 ;
        RECT 72.280 115.670 72.610 116.170 ;
        RECT 71.150 115.500 72.610 115.670 ;
        RECT 67.450 114.350 67.460 114.520 ;
        RECT 67.630 114.350 67.820 114.520 ;
        RECT 67.990 114.350 68.010 114.520 ;
        RECT 67.450 114.270 68.010 114.350 ;
        RECT 69.370 114.470 70.820 115.340 ;
        RECT 71.150 114.570 71.480 115.500 ;
        RECT 69.370 114.300 69.620 114.470 ;
        RECT 69.790 114.300 69.980 114.470 ;
        RECT 70.150 114.300 70.420 114.470 ;
        RECT 70.590 114.300 70.820 114.470 ;
        RECT 71.670 114.520 72.260 115.300 ;
        RECT 71.670 114.350 71.700 114.520 ;
        RECT 71.870 114.350 72.060 114.520 ;
        RECT 72.230 114.350 72.260 114.520 ;
        RECT 71.670 114.320 72.260 114.350 ;
        RECT 72.440 114.390 72.610 115.500 ;
        RECT 72.790 116.110 73.060 117.030 ;
        RECT 73.240 117.460 73.270 117.630 ;
        RECT 73.440 117.460 73.630 117.630 ;
        RECT 73.800 117.460 73.830 117.630 ;
        RECT 78.200 117.630 79.150 117.660 ;
        RECT 73.240 116.780 73.830 117.460 ;
      LAYER li1 ;
        RECT 74.110 117.400 77.050 117.570 ;
        RECT 74.110 116.410 74.280 117.400 ;
      LAYER li1 ;
        RECT 72.790 115.880 73.320 116.110 ;
        RECT 72.790 114.570 73.040 115.880 ;
      LAYER li1 ;
        RECT 73.740 115.540 74.280 116.410 ;
        RECT 74.460 115.920 74.790 117.220 ;
      LAYER li1 ;
        RECT 74.970 116.700 75.240 117.200 ;
        RECT 75.690 116.950 76.020 117.200 ;
        RECT 75.690 116.780 76.700 116.950 ;
        RECT 74.970 115.710 75.140 116.700 ;
        RECT 76.020 116.110 76.350 116.600 ;
        RECT 74.920 115.540 75.140 115.710 ;
        RECT 75.320 115.880 76.350 116.110 ;
        RECT 76.530 116.550 76.700 116.780 ;
      LAYER li1 ;
        RECT 76.880 116.900 77.050 117.400 ;
      LAYER li1 ;
        RECT 78.200 117.460 78.230 117.630 ;
        RECT 78.400 117.460 78.590 117.630 ;
        RECT 78.760 117.460 78.950 117.630 ;
        RECT 79.120 117.460 79.150 117.630 ;
        RECT 78.200 117.080 79.150 117.460 ;
      LAYER li1 ;
        RECT 79.330 117.590 81.990 117.760 ;
        RECT 79.330 116.900 79.500 117.590 ;
        RECT 76.880 116.730 79.500 116.900 ;
      LAYER li1 ;
        RECT 76.530 116.380 79.150 116.550 ;
        RECT 74.920 115.360 75.090 115.540 ;
        RECT 75.320 115.360 75.490 115.880 ;
        RECT 76.530 115.700 76.700 116.380 ;
      LAYER li1 ;
        RECT 79.330 116.200 79.500 116.730 ;
      LAYER li1 ;
        RECT 73.280 115.190 75.090 115.360 ;
        RECT 73.280 114.570 73.530 115.190 ;
        RECT 73.710 114.840 74.740 115.010 ;
        RECT 73.710 114.390 73.880 114.840 ;
        RECT 69.370 114.270 70.820 114.300 ;
        RECT 72.440 114.220 73.880 114.390 ;
        RECT 74.060 114.520 74.390 114.660 ;
        RECT 74.060 114.350 74.090 114.520 ;
        RECT 74.260 114.350 74.390 114.520 ;
        RECT 74.060 114.320 74.390 114.350 ;
        RECT 74.570 114.390 74.740 114.840 ;
        RECT 74.920 114.570 75.090 115.190 ;
        RECT 75.270 115.030 75.490 115.360 ;
        RECT 75.670 115.530 76.700 115.700 ;
        RECT 76.880 115.850 77.210 116.200 ;
      LAYER li1 ;
        RECT 77.650 116.030 79.500 116.200 ;
      LAYER li1 ;
        RECT 79.680 116.700 80.010 117.410 ;
        RECT 80.470 117.240 81.640 117.410 ;
        RECT 80.470 116.700 80.800 117.240 ;
        RECT 79.680 115.850 79.940 116.700 ;
        RECT 81.010 116.440 81.290 116.940 ;
        RECT 76.880 115.680 79.940 115.850 ;
        RECT 75.670 114.830 75.840 115.530 ;
        RECT 76.530 115.500 76.700 115.530 ;
        RECT 76.020 115.150 76.350 115.350 ;
        RECT 76.530 115.330 78.300 115.500 ;
        RECT 76.020 115.030 77.790 115.150 ;
        RECT 76.140 114.980 77.790 115.030 ;
        RECT 75.620 114.570 75.950 114.830 ;
        RECT 76.140 114.390 76.310 114.980 ;
        RECT 74.570 114.220 76.310 114.390 ;
        RECT 76.490 114.520 77.440 114.800 ;
        RECT 76.490 114.350 76.520 114.520 ;
        RECT 76.690 114.350 76.880 114.520 ;
        RECT 77.050 114.350 77.240 114.520 ;
        RECT 77.410 114.350 77.440 114.520 ;
        RECT 76.490 114.320 77.440 114.350 ;
        RECT 77.620 114.390 77.790 114.980 ;
        RECT 77.970 114.570 78.300 115.330 ;
        RECT 79.610 115.100 79.940 115.680 ;
        RECT 80.120 116.270 81.290 116.440 ;
        RECT 80.120 114.920 80.290 116.270 ;
        RECT 80.670 115.590 81.000 116.090 ;
        RECT 81.470 115.840 81.640 117.240 ;
      LAYER li1 ;
        RECT 81.820 116.930 81.990 117.590 ;
      LAYER li1 ;
        RECT 82.170 117.630 83.120 117.660 ;
        RECT 82.170 117.460 82.200 117.630 ;
        RECT 82.370 117.460 82.560 117.630 ;
        RECT 82.730 117.460 82.920 117.630 ;
        RECT 83.090 117.460 83.120 117.630 ;
        RECT 84.780 117.630 85.730 117.660 ;
        RECT 82.170 117.110 83.120 117.460 ;
        RECT 83.660 117.030 83.990 117.530 ;
        RECT 84.780 117.460 84.810 117.630 ;
        RECT 84.980 117.460 85.170 117.630 ;
        RECT 85.340 117.460 85.530 117.630 ;
        RECT 85.700 117.460 85.730 117.630 ;
      LAYER li1 ;
        RECT 81.820 116.760 82.830 116.930 ;
      LAYER li1 ;
        RECT 81.850 116.190 82.180 116.580 ;
      LAYER li1 ;
        RECT 82.500 116.370 82.830 116.760 ;
      LAYER li1 ;
        RECT 83.660 116.190 83.890 117.030 ;
        RECT 84.270 116.530 84.600 117.030 ;
        RECT 84.780 116.530 85.730 117.460 ;
        RECT 86.570 117.630 88.180 117.660 ;
        RECT 89.350 117.630 90.600 117.660 ;
        RECT 91.370 117.630 92.980 117.660 ;
        RECT 93.680 117.630 94.570 117.660 ;
        RECT 86.570 117.460 86.620 117.630 ;
        RECT 86.790 117.460 87.060 117.630 ;
        RECT 87.230 117.460 87.500 117.630 ;
        RECT 87.670 117.460 87.910 117.630 ;
        RECT 88.080 117.460 88.180 117.630 ;
        RECT 81.850 116.020 83.890 116.190 ;
        RECT 81.180 115.670 83.540 115.840 ;
        RECT 81.180 115.350 81.350 115.670 ;
        RECT 83.720 115.490 83.890 116.020 ;
        RECT 78.480 114.750 80.290 114.920 ;
        RECT 80.470 115.180 81.350 115.350 ;
        RECT 78.480 114.390 78.650 114.750 ;
        RECT 77.620 114.220 78.650 114.390 ;
        RECT 78.830 114.520 79.780 114.570 ;
        RECT 78.830 114.350 78.860 114.520 ;
        RECT 79.030 114.350 79.220 114.520 ;
        RECT 79.390 114.350 79.580 114.520 ;
        RECT 79.750 114.350 79.780 114.520 ;
        RECT 78.830 114.270 79.780 114.350 ;
        RECT 80.470 114.270 80.720 115.180 ;
        RECT 81.530 114.520 82.480 115.350 ;
        RECT 82.880 115.320 83.890 115.490 ;
        RECT 84.390 116.350 84.600 116.530 ;
        RECT 84.390 116.020 85.760 116.350 ;
        RECT 82.880 114.850 83.130 115.320 ;
        RECT 83.310 114.520 84.210 115.140 ;
        RECT 84.390 115.020 84.640 116.020 ;
        RECT 81.530 114.350 81.560 114.520 ;
        RECT 81.730 114.350 81.920 114.520 ;
        RECT 82.090 114.350 82.280 114.520 ;
        RECT 82.450 114.350 82.480 114.520 ;
        RECT 83.480 114.350 83.670 114.520 ;
        RECT 83.840 114.350 84.030 114.520 ;
        RECT 84.200 114.350 84.210 114.520 ;
        RECT 81.530 114.320 82.480 114.350 ;
        RECT 83.310 114.320 84.210 114.350 ;
        RECT 84.820 114.520 85.760 115.830 ;
        RECT 84.820 114.350 84.840 114.520 ;
        RECT 85.010 114.350 85.200 114.520 ;
        RECT 85.370 114.350 85.560 114.520 ;
        RECT 85.730 114.350 85.760 114.520 ;
        RECT 84.820 114.290 85.760 114.350 ;
      LAYER li1 ;
        RECT 85.940 114.290 86.280 117.360 ;
      LAYER li1 ;
        RECT 86.570 117.180 88.180 117.460 ;
        RECT 86.880 116.780 88.180 117.180 ;
        RECT 86.880 116.000 87.210 116.780 ;
        RECT 87.420 115.340 87.750 116.330 ;
      LAYER li1 ;
        RECT 88.920 115.850 89.170 117.530 ;
      LAYER li1 ;
        RECT 89.520 117.460 89.710 117.630 ;
        RECT 89.880 117.460 90.070 117.630 ;
        RECT 90.240 117.460 90.430 117.630 ;
        RECT 89.350 117.090 90.600 117.460 ;
        RECT 90.780 116.910 91.030 117.530 ;
        RECT 91.370 117.460 91.420 117.630 ;
        RECT 91.590 117.460 91.860 117.630 ;
        RECT 92.030 117.460 92.300 117.630 ;
        RECT 92.470 117.460 92.710 117.630 ;
        RECT 92.880 117.460 92.980 117.630 ;
        RECT 91.370 117.180 92.980 117.460 ;
        RECT 89.480 116.740 91.030 116.910 ;
        RECT 89.480 116.280 89.810 116.740 ;
        RECT 86.650 114.470 88.100 115.340 ;
        RECT 86.650 114.300 86.900 114.470 ;
        RECT 87.070 114.300 87.260 114.470 ;
        RECT 87.430 114.300 87.700 114.470 ;
        RECT 87.870 114.300 88.100 114.470 ;
        RECT 86.650 114.270 88.100 114.300 ;
      LAYER li1 ;
        RECT 88.920 114.270 89.350 115.850 ;
      LAYER li1 ;
        RECT 89.530 114.520 90.090 115.850 ;
      LAYER li1 ;
        RECT 90.270 114.770 90.600 116.560 ;
      LAYER li1 ;
        RECT 90.780 115.020 91.030 116.740 ;
        RECT 91.680 116.780 92.980 117.180 ;
        RECT 91.680 116.000 92.010 116.780 ;
        RECT 92.220 115.340 92.550 116.330 ;
        RECT 89.530 114.350 89.540 114.520 ;
        RECT 89.710 114.350 89.900 114.520 ;
        RECT 90.070 114.350 90.090 114.520 ;
        RECT 89.530 114.270 90.090 114.350 ;
        RECT 91.450 114.470 92.900 115.340 ;
        RECT 91.450 114.300 91.700 114.470 ;
        RECT 91.870 114.300 92.060 114.470 ;
        RECT 92.230 114.300 92.500 114.470 ;
        RECT 92.670 114.300 92.900 114.470 ;
        RECT 91.450 114.270 92.900 114.300 ;
      LAYER li1 ;
        RECT 93.250 114.270 93.500 117.530 ;
      LAYER li1 ;
        RECT 93.850 117.460 94.040 117.630 ;
        RECT 94.210 117.460 94.400 117.630 ;
        RECT 94.870 117.590 96.800 117.760 ;
        RECT 93.680 116.780 94.570 117.460 ;
        RECT 94.870 117.160 95.200 117.590 ;
        RECT 95.650 117.150 95.980 117.410 ;
        RECT 95.380 116.980 95.980 117.150 ;
        RECT 96.470 117.000 96.800 117.590 ;
        RECT 97.010 117.630 98.310 117.660 ;
        RECT 97.010 117.460 97.040 117.630 ;
        RECT 97.210 117.460 97.400 117.630 ;
        RECT 97.570 117.460 97.760 117.630 ;
        RECT 97.930 117.460 98.120 117.630 ;
        RECT 98.290 117.460 98.310 117.630 ;
        RECT 97.010 116.980 98.310 117.460 ;
        RECT 98.570 117.630 100.180 117.660 ;
        RECT 100.870 117.630 102.120 117.660 ;
        RECT 102.890 117.630 104.500 117.660 ;
        RECT 98.570 117.460 98.620 117.630 ;
        RECT 98.790 117.460 99.060 117.630 ;
        RECT 99.230 117.460 99.500 117.630 ;
        RECT 99.670 117.460 99.910 117.630 ;
        RECT 100.080 117.460 100.180 117.630 ;
        RECT 98.570 117.180 100.180 117.460 ;
        RECT 94.750 116.810 95.550 116.980 ;
        RECT 94.750 116.600 94.920 116.810 ;
      LAYER li1 ;
        RECT 96.160 116.800 96.830 116.820 ;
        RECT 95.730 116.630 98.000 116.800 ;
      LAYER li1 ;
        RECT 93.710 116.430 94.920 116.600 ;
      LAYER li1 ;
        RECT 95.100 116.460 95.900 116.630 ;
      LAYER li1 ;
        RECT 93.710 115.730 94.040 116.430 ;
      LAYER li1 ;
        RECT 95.100 116.250 95.270 116.460 ;
        RECT 97.670 116.450 98.000 116.630 ;
        RECT 94.540 115.970 95.270 116.250 ;
        RECT 95.450 115.910 95.880 116.280 ;
        RECT 96.080 115.910 96.370 116.450 ;
        RECT 96.610 116.120 97.320 116.450 ;
        RECT 97.590 116.280 98.000 116.450 ;
        RECT 97.670 116.010 98.000 116.280 ;
      LAYER li1 ;
        RECT 98.880 116.780 100.180 117.180 ;
        RECT 98.880 116.000 99.210 116.780 ;
        RECT 96.550 115.730 96.800 115.850 ;
        RECT 93.710 115.560 96.800 115.730 ;
        RECT 93.680 114.520 96.370 115.380 ;
        RECT 93.850 114.350 94.040 114.520 ;
        RECT 94.210 114.350 94.400 114.520 ;
        RECT 94.570 114.350 94.760 114.520 ;
        RECT 94.930 114.350 95.120 114.520 ;
        RECT 95.290 114.350 95.480 114.520 ;
        RECT 95.650 114.350 95.840 114.520 ;
        RECT 96.010 114.350 96.200 114.520 ;
        RECT 93.680 114.270 96.370 114.350 ;
        RECT 96.550 114.270 96.800 115.560 ;
        RECT 96.980 114.520 98.290 115.830 ;
        RECT 99.420 115.340 99.750 116.330 ;
      LAYER li1 ;
        RECT 100.440 115.850 100.690 117.530 ;
      LAYER li1 ;
        RECT 101.040 117.460 101.230 117.630 ;
        RECT 101.400 117.460 101.590 117.630 ;
        RECT 101.760 117.460 101.950 117.630 ;
        RECT 100.870 117.090 102.120 117.460 ;
        RECT 102.300 116.910 102.550 117.530 ;
        RECT 102.890 117.460 102.940 117.630 ;
        RECT 103.110 117.460 103.380 117.630 ;
        RECT 103.550 117.460 103.820 117.630 ;
        RECT 103.990 117.460 104.230 117.630 ;
        RECT 104.400 117.460 104.500 117.630 ;
        RECT 102.890 117.180 104.500 117.460 ;
        RECT 101.000 116.740 102.550 116.910 ;
        RECT 101.000 116.280 101.330 116.740 ;
        RECT 96.980 114.350 97.010 114.520 ;
        RECT 97.180 114.350 97.370 114.520 ;
        RECT 97.540 114.350 97.730 114.520 ;
        RECT 97.900 114.350 98.090 114.520 ;
        RECT 98.260 114.350 98.290 114.520 ;
        RECT 96.980 114.290 98.290 114.350 ;
        RECT 98.650 114.470 100.100 115.340 ;
        RECT 98.650 114.300 98.900 114.470 ;
        RECT 99.070 114.300 99.260 114.470 ;
        RECT 99.430 114.300 99.700 114.470 ;
        RECT 99.870 114.300 100.100 114.470 ;
        RECT 98.650 114.270 100.100 114.300 ;
      LAYER li1 ;
        RECT 100.440 114.270 100.870 115.850 ;
      LAYER li1 ;
        RECT 101.050 114.520 101.610 115.850 ;
      LAYER li1 ;
        RECT 101.790 114.770 102.120 116.560 ;
      LAYER li1 ;
        RECT 102.300 115.020 102.550 116.740 ;
        RECT 103.200 116.780 104.500 117.180 ;
        RECT 104.730 117.630 105.680 117.660 ;
        RECT 104.730 117.460 104.760 117.630 ;
        RECT 104.930 117.460 105.120 117.630 ;
        RECT 105.290 117.460 105.480 117.630 ;
        RECT 105.650 117.460 105.680 117.630 ;
        RECT 106.290 117.630 107.240 117.660 ;
        RECT 103.200 116.000 103.530 116.780 ;
        RECT 104.730 116.700 105.680 117.460 ;
      LAYER li1 ;
        RECT 105.860 116.820 106.110 117.530 ;
      LAYER li1 ;
        RECT 106.290 117.460 106.320 117.630 ;
        RECT 106.490 117.460 106.680 117.630 ;
        RECT 106.850 117.460 107.040 117.630 ;
        RECT 107.210 117.460 107.240 117.630 ;
        RECT 107.850 117.630 108.800 117.660 ;
        RECT 106.290 117.000 107.240 117.460 ;
      LAYER li1 ;
        RECT 107.420 116.820 107.670 117.530 ;
        RECT 105.860 116.650 107.670 116.820 ;
      LAYER li1 ;
        RECT 107.850 117.460 107.880 117.630 ;
        RECT 108.050 117.460 108.240 117.630 ;
        RECT 108.410 117.460 108.600 117.630 ;
        RECT 108.770 117.460 108.800 117.630 ;
        RECT 109.610 117.630 111.220 117.660 ;
        RECT 111.910 117.630 113.160 117.660 ;
        RECT 113.930 117.630 115.540 117.660 ;
        RECT 117.670 117.630 118.920 117.660 ;
        RECT 119.690 117.630 121.300 117.660 ;
        RECT 107.850 116.780 108.800 117.460 ;
      LAYER li1 ;
        RECT 105.860 116.480 106.030 116.650 ;
      LAYER li1 ;
        RECT 108.980 116.600 109.310 117.530 ;
        RECT 109.610 117.460 109.660 117.630 ;
        RECT 109.830 117.460 110.100 117.630 ;
        RECT 110.270 117.460 110.540 117.630 ;
        RECT 110.710 117.460 110.950 117.630 ;
        RECT 111.120 117.460 111.220 117.630 ;
        RECT 109.610 117.180 111.220 117.460 ;
        RECT 103.740 115.340 104.070 116.330 ;
      LAYER li1 ;
        RECT 104.770 116.250 106.030 116.480 ;
      LAYER li1 ;
        RECT 108.070 116.470 109.310 116.600 ;
        RECT 106.210 116.430 109.310 116.470 ;
        RECT 106.210 116.300 108.240 116.430 ;
      LAYER li1 ;
        RECT 105.860 116.120 106.030 116.250 ;
        RECT 105.860 115.950 107.750 116.120 ;
      LAYER li1 ;
        RECT 101.050 114.350 101.060 114.520 ;
        RECT 101.230 114.350 101.420 114.520 ;
        RECT 101.590 114.350 101.610 114.520 ;
        RECT 101.050 114.270 101.610 114.350 ;
        RECT 102.970 114.470 104.420 115.340 ;
        RECT 102.970 114.300 103.220 114.470 ;
        RECT 103.390 114.300 103.580 114.470 ;
        RECT 103.750 114.300 104.020 114.470 ;
        RECT 104.190 114.300 104.420 114.470 ;
        RECT 102.970 114.270 104.420 114.300 ;
        RECT 104.730 114.520 105.680 115.850 ;
        RECT 104.730 114.350 104.760 114.520 ;
        RECT 104.930 114.350 105.120 114.520 ;
        RECT 105.290 114.350 105.480 114.520 ;
        RECT 105.650 114.350 105.680 114.520 ;
        RECT 104.730 114.270 105.680 114.350 ;
      LAYER li1 ;
        RECT 105.860 114.270 106.110 115.950 ;
      LAYER li1 ;
        RECT 106.290 114.520 107.240 115.770 ;
        RECT 106.290 114.350 106.320 114.520 ;
        RECT 106.490 114.350 106.680 114.520 ;
        RECT 106.850 114.350 107.040 114.520 ;
        RECT 107.210 114.350 107.240 114.520 ;
        RECT 106.290 114.270 107.240 114.350 ;
      LAYER li1 ;
        RECT 107.420 114.270 107.750 115.950 ;
        RECT 108.530 115.910 108.860 116.250 ;
      LAYER li1 ;
        RECT 107.930 114.520 108.880 115.730 ;
        RECT 107.930 114.350 107.960 114.520 ;
        RECT 108.130 114.350 108.320 114.520 ;
        RECT 108.490 114.350 108.680 114.520 ;
        RECT 108.850 114.350 108.880 114.520 ;
        RECT 107.930 114.270 108.880 114.350 ;
        RECT 109.060 114.270 109.310 116.430 ;
        RECT 109.920 116.780 111.220 117.180 ;
        RECT 109.920 116.000 110.250 116.780 ;
        RECT 110.460 115.340 110.790 116.330 ;
      LAYER li1 ;
        RECT 111.480 115.850 111.730 117.530 ;
      LAYER li1 ;
        RECT 112.080 117.460 112.270 117.630 ;
        RECT 112.440 117.460 112.630 117.630 ;
        RECT 112.800 117.460 112.990 117.630 ;
        RECT 111.910 117.090 113.160 117.460 ;
        RECT 113.340 116.910 113.590 117.530 ;
        RECT 113.930 117.460 113.980 117.630 ;
        RECT 114.150 117.460 114.420 117.630 ;
        RECT 114.590 117.460 114.860 117.630 ;
        RECT 115.030 117.460 115.270 117.630 ;
        RECT 115.440 117.460 115.540 117.630 ;
        RECT 113.930 117.180 115.540 117.460 ;
        RECT 112.040 116.740 113.590 116.910 ;
        RECT 112.040 116.280 112.370 116.740 ;
        RECT 109.690 114.470 111.140 115.340 ;
        RECT 109.690 114.300 109.940 114.470 ;
        RECT 110.110 114.300 110.300 114.470 ;
        RECT 110.470 114.300 110.740 114.470 ;
        RECT 110.910 114.300 111.140 114.470 ;
        RECT 109.690 114.270 111.140 114.300 ;
      LAYER li1 ;
        RECT 111.480 114.270 111.910 115.850 ;
      LAYER li1 ;
        RECT 112.090 114.520 112.650 115.850 ;
      LAYER li1 ;
        RECT 112.830 114.770 113.160 116.560 ;
      LAYER li1 ;
        RECT 113.340 115.020 113.590 116.740 ;
        RECT 114.240 116.780 115.540 117.180 ;
        RECT 114.240 116.000 114.570 116.780 ;
        RECT 114.780 115.340 115.110 116.330 ;
      LAYER li1 ;
        RECT 117.240 115.850 117.490 117.530 ;
      LAYER li1 ;
        RECT 117.840 117.460 118.030 117.630 ;
        RECT 118.200 117.460 118.390 117.630 ;
        RECT 118.560 117.460 118.750 117.630 ;
        RECT 117.670 117.090 118.920 117.460 ;
        RECT 119.100 116.910 119.350 117.530 ;
        RECT 119.690 117.460 119.740 117.630 ;
        RECT 119.910 117.460 120.180 117.630 ;
        RECT 120.350 117.460 120.620 117.630 ;
        RECT 120.790 117.460 121.030 117.630 ;
        RECT 121.200 117.460 121.300 117.630 ;
        RECT 119.690 117.180 121.300 117.460 ;
        RECT 117.800 116.740 119.350 116.910 ;
        RECT 117.800 116.280 118.130 116.740 ;
        RECT 112.090 114.350 112.100 114.520 ;
        RECT 112.270 114.350 112.460 114.520 ;
        RECT 112.630 114.350 112.650 114.520 ;
        RECT 112.090 114.270 112.650 114.350 ;
        RECT 114.010 114.470 115.460 115.340 ;
        RECT 114.010 114.300 114.260 114.470 ;
        RECT 114.430 114.300 114.620 114.470 ;
        RECT 114.790 114.300 115.060 114.470 ;
        RECT 115.230 114.300 115.460 114.470 ;
        RECT 114.010 114.270 115.460 114.300 ;
      LAYER li1 ;
        RECT 117.240 114.270 117.670 115.850 ;
      LAYER li1 ;
        RECT 117.850 114.520 118.410 115.850 ;
      LAYER li1 ;
        RECT 118.590 114.770 118.920 116.560 ;
      LAYER li1 ;
        RECT 119.100 115.020 119.350 116.740 ;
        RECT 120.000 116.780 121.300 117.180 ;
        RECT 121.530 117.630 122.120 117.660 ;
        RECT 121.530 117.460 121.560 117.630 ;
        RECT 121.730 117.460 121.920 117.630 ;
        RECT 122.090 117.460 122.120 117.630 ;
        RECT 123.460 117.640 126.190 117.670 ;
        RECT 120.000 116.000 120.330 116.780 ;
        RECT 121.530 116.700 122.120 117.460 ;
        RECT 120.540 115.340 120.870 116.330 ;
      LAYER li1 ;
        RECT 121.570 116.090 122.280 116.480 ;
        RECT 122.460 115.850 122.790 117.530 ;
      LAYER li1 ;
        RECT 123.460 117.470 123.630 117.640 ;
        RECT 123.800 117.470 124.070 117.640 ;
        RECT 124.240 117.470 124.480 117.640 ;
        RECT 124.650 117.470 124.910 117.640 ;
        RECT 125.080 117.470 125.350 117.640 ;
        RECT 125.520 117.470 125.760 117.640 ;
        RECT 125.930 117.470 126.190 117.640 ;
        RECT 123.460 116.670 126.190 117.470 ;
        RECT 127.300 117.640 130.030 117.670 ;
        RECT 127.300 117.470 127.470 117.640 ;
        RECT 127.640 117.470 127.910 117.640 ;
        RECT 128.080 117.470 128.320 117.640 ;
        RECT 128.490 117.470 128.750 117.640 ;
        RECT 128.920 117.470 129.190 117.640 ;
        RECT 129.360 117.470 129.600 117.640 ;
        RECT 129.770 117.470 130.030 117.640 ;
        RECT 127.300 116.670 130.030 117.470 ;
        RECT 131.140 117.640 133.870 117.670 ;
        RECT 131.140 117.470 131.310 117.640 ;
        RECT 131.480 117.470 131.750 117.640 ;
        RECT 131.920 117.470 132.160 117.640 ;
        RECT 132.330 117.470 132.590 117.640 ;
        RECT 132.760 117.470 133.030 117.640 ;
        RECT 133.200 117.470 133.440 117.640 ;
        RECT 133.610 117.470 133.870 117.640 ;
        RECT 131.140 116.670 133.870 117.470 ;
        RECT 134.980 117.640 137.710 117.670 ;
        RECT 134.980 117.470 135.150 117.640 ;
        RECT 135.320 117.470 135.590 117.640 ;
        RECT 135.760 117.470 136.000 117.640 ;
        RECT 136.170 117.470 136.430 117.640 ;
        RECT 136.600 117.470 136.870 117.640 ;
        RECT 137.040 117.470 137.280 117.640 ;
        RECT 137.450 117.470 137.710 117.640 ;
        RECT 134.980 116.670 137.710 117.470 ;
        RECT 138.820 117.640 141.550 117.670 ;
        RECT 138.820 117.470 138.990 117.640 ;
        RECT 139.160 117.470 139.430 117.640 ;
        RECT 139.600 117.470 139.840 117.640 ;
        RECT 140.010 117.470 140.270 117.640 ;
        RECT 140.440 117.470 140.710 117.640 ;
        RECT 140.880 117.470 141.120 117.640 ;
        RECT 141.290 117.470 141.550 117.640 ;
        RECT 138.820 116.670 141.550 117.470 ;
        RECT 123.620 116.000 123.950 116.670 ;
        RECT 117.850 114.350 117.860 114.520 ;
        RECT 118.030 114.350 118.220 114.520 ;
        RECT 118.390 114.350 118.410 114.520 ;
        RECT 117.850 114.270 118.410 114.350 ;
        RECT 119.770 114.470 121.220 115.340 ;
        RECT 119.770 114.300 120.020 114.470 ;
        RECT 120.190 114.300 120.380 114.470 ;
        RECT 120.550 114.300 120.820 114.470 ;
        RECT 120.990 114.300 121.220 114.470 ;
        RECT 119.770 114.270 121.220 114.300 ;
        RECT 121.530 114.520 122.120 115.850 ;
        RECT 121.530 114.350 121.560 114.520 ;
        RECT 121.730 114.350 121.920 114.520 ;
        RECT 122.090 114.350 122.120 114.520 ;
        RECT 121.530 114.270 122.120 114.350 ;
      LAYER li1 ;
        RECT 122.400 114.270 122.790 115.850 ;
      LAYER li1 ;
        RECT 124.350 115.350 124.680 116.330 ;
        RECT 124.900 116.000 125.230 116.670 ;
        RECT 125.630 115.350 125.960 116.330 ;
        RECT 127.460 116.000 127.790 116.670 ;
        RECT 128.190 115.350 128.520 116.330 ;
        RECT 128.740 116.000 129.070 116.670 ;
        RECT 129.470 115.350 129.800 116.330 ;
        RECT 131.300 116.000 131.630 116.670 ;
        RECT 132.030 115.350 132.360 116.330 ;
        RECT 132.580 116.000 132.910 116.670 ;
        RECT 133.310 115.350 133.640 116.330 ;
        RECT 135.140 116.000 135.470 116.670 ;
        RECT 135.870 115.350 136.200 116.330 ;
        RECT 136.420 116.000 136.750 116.670 ;
        RECT 137.150 115.350 137.480 116.330 ;
        RECT 138.980 116.000 139.310 116.670 ;
        RECT 139.710 115.350 140.040 116.330 ;
        RECT 140.260 116.000 140.590 116.670 ;
        RECT 140.990 115.350 141.320 116.330 ;
        RECT 123.380 114.470 126.120 115.350 ;
        RECT 123.380 114.300 123.590 114.470 ;
        RECT 123.760 114.300 124.030 114.470 ;
        RECT 124.200 114.300 124.440 114.470 ;
        RECT 124.610 114.300 124.870 114.470 ;
        RECT 125.040 114.300 125.310 114.470 ;
        RECT 125.480 114.300 125.720 114.470 ;
        RECT 125.890 114.300 126.120 114.470 ;
        RECT 123.380 114.280 126.120 114.300 ;
        RECT 127.220 114.470 129.960 115.350 ;
        RECT 127.220 114.300 127.430 114.470 ;
        RECT 127.600 114.300 127.870 114.470 ;
        RECT 128.040 114.300 128.280 114.470 ;
        RECT 128.450 114.300 128.710 114.470 ;
        RECT 128.880 114.300 129.150 114.470 ;
        RECT 129.320 114.300 129.560 114.470 ;
        RECT 129.730 114.300 129.960 114.470 ;
        RECT 127.220 114.280 129.960 114.300 ;
        RECT 131.060 114.470 133.800 115.350 ;
        RECT 131.060 114.300 131.270 114.470 ;
        RECT 131.440 114.300 131.710 114.470 ;
        RECT 131.880 114.300 132.120 114.470 ;
        RECT 132.290 114.300 132.550 114.470 ;
        RECT 132.720 114.300 132.990 114.470 ;
        RECT 133.160 114.300 133.400 114.470 ;
        RECT 133.570 114.300 133.800 114.470 ;
        RECT 131.060 114.280 133.800 114.300 ;
        RECT 134.900 114.470 137.640 115.350 ;
        RECT 134.900 114.300 135.110 114.470 ;
        RECT 135.280 114.300 135.550 114.470 ;
        RECT 135.720 114.300 135.960 114.470 ;
        RECT 136.130 114.300 136.390 114.470 ;
        RECT 136.560 114.300 136.830 114.470 ;
        RECT 137.000 114.300 137.240 114.470 ;
        RECT 137.410 114.300 137.640 114.470 ;
        RECT 134.900 114.280 137.640 114.300 ;
        RECT 138.740 114.470 141.480 115.350 ;
        RECT 138.740 114.300 138.950 114.470 ;
        RECT 139.120 114.300 139.390 114.470 ;
        RECT 139.560 114.300 139.800 114.470 ;
        RECT 139.970 114.300 140.230 114.470 ;
        RECT 140.400 114.300 140.670 114.470 ;
        RECT 140.840 114.300 141.080 114.470 ;
        RECT 141.250 114.300 141.480 114.470 ;
        RECT 138.740 114.280 141.480 114.300 ;
        RECT 5.760 113.870 5.920 114.050 ;
        RECT 6.090 113.870 6.400 114.050 ;
        RECT 6.570 113.870 6.880 114.050 ;
        RECT 7.050 113.870 7.360 114.050 ;
        RECT 7.530 113.870 7.840 114.050 ;
        RECT 8.010 113.870 8.320 114.050 ;
        RECT 8.490 113.870 8.800 114.050 ;
        RECT 8.970 113.870 9.280 114.050 ;
        RECT 9.450 113.870 9.760 114.050 ;
        RECT 9.930 113.870 10.240 114.050 ;
        RECT 10.410 113.870 10.720 114.050 ;
        RECT 10.890 113.870 11.200 114.050 ;
        RECT 11.370 113.870 11.680 114.050 ;
        RECT 11.850 113.870 12.160 114.050 ;
        RECT 12.330 113.870 12.640 114.050 ;
        RECT 12.810 113.870 13.120 114.050 ;
        RECT 13.290 114.040 13.600 114.050 ;
        RECT 13.770 114.040 14.080 114.050 ;
        RECT 13.290 113.870 13.440 114.040 ;
        RECT 13.920 113.870 14.080 114.040 ;
        RECT 14.250 113.870 14.560 114.050 ;
        RECT 14.730 113.870 15.040 114.050 ;
        RECT 15.210 113.870 15.520 114.050 ;
        RECT 15.690 113.870 16.000 114.050 ;
        RECT 16.170 113.870 16.480 114.050 ;
        RECT 16.650 113.870 16.960 114.050 ;
        RECT 17.130 113.870 17.440 114.050 ;
        RECT 17.610 113.870 17.920 114.050 ;
        RECT 18.090 113.870 18.400 114.050 ;
        RECT 18.570 113.870 18.880 114.050 ;
        RECT 19.050 113.870 19.360 114.050 ;
        RECT 19.530 113.870 19.840 114.050 ;
        RECT 20.010 113.870 20.320 114.050 ;
        RECT 20.490 113.870 20.800 114.050 ;
        RECT 20.970 113.870 21.280 114.050 ;
        RECT 21.450 113.870 21.760 114.050 ;
        RECT 21.930 113.870 22.240 114.050 ;
        RECT 22.410 113.870 22.720 114.050 ;
        RECT 22.890 113.870 23.200 114.050 ;
        RECT 23.370 113.870 23.680 114.050 ;
        RECT 23.850 114.040 24.000 114.050 ;
        RECT 24.480 114.040 24.640 114.050 ;
        RECT 23.850 113.870 24.160 114.040 ;
        RECT 24.330 113.870 24.640 114.040 ;
        RECT 24.810 113.870 25.120 114.050 ;
        RECT 25.290 113.870 25.600 114.050 ;
        RECT 25.770 113.870 26.080 114.050 ;
        RECT 26.250 113.870 26.560 114.050 ;
        RECT 26.730 113.870 27.040 114.050 ;
        RECT 27.210 113.870 27.520 114.050 ;
        RECT 27.690 113.870 28.000 114.050 ;
        RECT 28.170 113.870 28.480 114.050 ;
        RECT 28.650 113.870 28.960 114.050 ;
        RECT 29.130 113.870 29.440 114.050 ;
        RECT 29.610 113.870 29.920 114.050 ;
        RECT 30.090 113.870 30.400 114.050 ;
        RECT 30.570 113.870 30.880 114.050 ;
        RECT 31.050 113.870 31.360 114.050 ;
        RECT 31.530 113.870 31.840 114.050 ;
        RECT 32.010 113.870 32.320 114.050 ;
        RECT 32.490 113.870 32.800 114.050 ;
        RECT 32.970 113.870 33.280 114.050 ;
        RECT 33.450 113.870 33.760 114.050 ;
        RECT 33.930 113.870 34.240 114.050 ;
        RECT 34.410 113.870 34.720 114.050 ;
        RECT 34.890 113.870 35.200 114.050 ;
        RECT 35.370 113.870 35.680 114.050 ;
        RECT 35.850 113.870 36.160 114.050 ;
        RECT 36.330 113.870 36.640 114.050 ;
        RECT 36.810 114.040 36.960 114.050 ;
        RECT 37.440 114.040 37.600 114.050 ;
        RECT 36.810 113.870 37.120 114.040 ;
        RECT 37.290 113.870 37.600 114.040 ;
        RECT 37.770 113.870 38.080 114.050 ;
        RECT 38.250 113.870 38.560 114.050 ;
        RECT 38.730 113.870 39.040 114.050 ;
        RECT 39.210 113.870 39.520 114.050 ;
        RECT 39.690 113.870 40.000 114.050 ;
        RECT 40.170 113.870 40.480 114.050 ;
        RECT 40.650 113.870 40.960 114.050 ;
        RECT 41.130 113.870 41.440 114.050 ;
        RECT 41.610 113.870 41.920 114.050 ;
        RECT 42.090 113.870 42.400 114.050 ;
        RECT 42.570 113.870 42.880 114.050 ;
        RECT 43.050 113.870 43.360 114.050 ;
        RECT 43.530 113.870 43.840 114.050 ;
        RECT 44.010 113.870 44.320 114.050 ;
        RECT 44.490 113.870 44.800 114.050 ;
        RECT 44.970 113.870 45.280 114.050 ;
        RECT 45.450 113.870 45.760 114.050 ;
        RECT 45.930 113.870 46.240 114.050 ;
        RECT 46.410 113.870 46.720 114.050 ;
        RECT 46.890 113.870 47.200 114.050 ;
        RECT 47.370 113.870 47.680 114.050 ;
        RECT 47.850 113.870 48.160 114.050 ;
        RECT 48.330 113.870 48.640 114.050 ;
        RECT 48.810 113.870 49.120 114.050 ;
        RECT 49.290 113.870 49.600 114.050 ;
        RECT 49.770 113.870 50.080 114.050 ;
        RECT 50.250 113.870 50.560 114.050 ;
        RECT 50.730 113.870 51.040 114.050 ;
        RECT 51.210 113.870 51.520 114.050 ;
        RECT 51.690 113.870 52.000 114.050 ;
        RECT 52.170 113.870 52.480 114.050 ;
        RECT 52.650 113.870 52.960 114.050 ;
        RECT 53.130 113.870 53.440 114.050 ;
        RECT 53.610 113.870 53.920 114.050 ;
        RECT 54.090 113.870 54.400 114.050 ;
        RECT 54.570 113.870 54.880 114.050 ;
        RECT 55.050 113.870 55.360 114.050 ;
        RECT 55.530 113.870 55.840 114.050 ;
        RECT 56.010 113.870 56.320 114.050 ;
        RECT 56.490 113.870 56.800 114.050 ;
        RECT 56.970 113.870 57.280 114.050 ;
        RECT 57.450 113.870 57.760 114.050 ;
        RECT 57.930 113.870 58.240 114.050 ;
        RECT 58.410 113.870 58.720 114.050 ;
        RECT 58.890 113.870 59.200 114.050 ;
        RECT 59.370 113.870 59.680 114.050 ;
        RECT 59.850 113.870 60.160 114.050 ;
        RECT 60.330 113.870 60.640 114.050 ;
        RECT 60.810 113.870 61.120 114.050 ;
        RECT 61.290 113.870 61.600 114.050 ;
        RECT 61.770 113.870 62.080 114.050 ;
        RECT 62.250 113.870 62.560 114.050 ;
        RECT 62.730 113.870 63.040 114.050 ;
        RECT 63.210 113.870 63.520 114.050 ;
        RECT 63.690 113.870 64.000 114.050 ;
        RECT 64.170 113.870 64.480 114.050 ;
        RECT 64.650 113.870 64.960 114.050 ;
        RECT 65.130 113.870 65.440 114.050 ;
        RECT 65.610 113.870 65.920 114.050 ;
        RECT 66.090 113.870 66.400 114.050 ;
        RECT 66.570 113.870 66.880 114.050 ;
        RECT 67.050 113.870 67.360 114.050 ;
        RECT 67.530 113.870 67.840 114.050 ;
        RECT 68.010 113.870 68.320 114.050 ;
        RECT 68.490 113.870 68.800 114.050 ;
        RECT 68.970 113.870 69.280 114.050 ;
        RECT 69.450 113.870 69.760 114.050 ;
        RECT 69.930 113.870 70.240 114.050 ;
        RECT 70.410 113.870 70.720 114.050 ;
        RECT 70.890 113.870 71.200 114.050 ;
        RECT 71.370 114.040 71.520 114.050 ;
        RECT 72.000 114.040 72.160 114.050 ;
        RECT 71.370 113.870 71.680 114.040 ;
        RECT 71.850 113.870 72.160 114.040 ;
        RECT 72.330 113.870 72.640 114.050 ;
        RECT 72.810 113.870 73.120 114.050 ;
        RECT 73.290 113.870 73.600 114.050 ;
        RECT 73.770 113.870 74.080 114.050 ;
        RECT 74.250 113.870 74.560 114.050 ;
        RECT 74.730 113.870 75.040 114.050 ;
        RECT 75.210 113.870 75.520 114.050 ;
        RECT 75.690 113.870 76.000 114.050 ;
        RECT 76.170 113.870 76.480 114.050 ;
        RECT 76.650 113.870 76.960 114.050 ;
        RECT 77.130 113.870 77.440 114.050 ;
        RECT 77.610 113.870 77.920 114.050 ;
        RECT 78.090 113.870 78.400 114.050 ;
        RECT 78.570 113.870 78.880 114.050 ;
        RECT 79.050 113.870 79.360 114.050 ;
        RECT 79.530 113.870 79.840 114.050 ;
        RECT 80.010 113.870 80.320 114.050 ;
        RECT 80.490 113.870 80.800 114.050 ;
        RECT 80.970 113.870 81.280 114.050 ;
        RECT 81.450 113.870 81.760 114.050 ;
        RECT 81.930 113.870 82.240 114.050 ;
        RECT 82.410 113.870 82.720 114.050 ;
        RECT 82.890 113.870 83.200 114.050 ;
        RECT 83.370 113.870 83.680 114.050 ;
        RECT 83.850 113.870 84.160 114.050 ;
        RECT 84.330 113.870 84.640 114.050 ;
        RECT 84.810 113.870 85.120 114.050 ;
        RECT 85.290 113.870 85.600 114.050 ;
        RECT 85.770 113.870 86.080 114.050 ;
        RECT 86.250 113.870 86.560 114.050 ;
        RECT 86.730 113.870 87.040 114.050 ;
        RECT 87.210 113.870 87.520 114.050 ;
        RECT 87.690 113.870 88.000 114.050 ;
        RECT 88.170 114.040 88.480 114.050 ;
        RECT 88.650 114.040 88.960 114.050 ;
        RECT 88.170 113.870 88.320 114.040 ;
        RECT 88.800 113.870 88.960 114.040 ;
        RECT 89.130 113.870 89.440 114.050 ;
        RECT 89.610 113.870 89.920 114.050 ;
        RECT 90.090 113.870 90.400 114.050 ;
        RECT 90.570 113.870 90.880 114.050 ;
        RECT 91.050 113.870 91.360 114.050 ;
        RECT 91.530 113.870 91.840 114.050 ;
        RECT 92.010 113.870 92.320 114.050 ;
        RECT 92.490 113.870 92.800 114.050 ;
        RECT 92.970 113.870 93.280 114.050 ;
        RECT 93.450 113.870 93.760 114.050 ;
        RECT 93.930 113.870 94.240 114.050 ;
        RECT 94.410 113.870 94.720 114.050 ;
        RECT 94.890 113.870 95.200 114.050 ;
        RECT 95.370 113.870 95.680 114.050 ;
        RECT 95.850 113.870 96.160 114.050 ;
        RECT 96.330 113.870 96.640 114.050 ;
        RECT 96.810 113.870 97.120 114.050 ;
        RECT 97.290 113.870 97.600 114.050 ;
        RECT 97.770 113.870 98.080 114.050 ;
        RECT 98.250 113.870 98.560 114.050 ;
        RECT 98.730 113.870 99.040 114.050 ;
        RECT 99.210 113.870 99.520 114.050 ;
        RECT 99.690 113.870 100.000 114.050 ;
        RECT 100.170 113.870 100.480 114.050 ;
        RECT 100.650 113.870 100.960 114.050 ;
        RECT 101.130 113.870 101.440 114.050 ;
        RECT 101.610 113.870 101.920 114.050 ;
        RECT 102.090 113.870 102.400 114.050 ;
        RECT 102.570 113.870 102.880 114.050 ;
        RECT 103.050 113.870 103.360 114.050 ;
        RECT 103.530 113.870 103.840 114.050 ;
        RECT 104.010 113.870 104.320 114.050 ;
        RECT 104.490 113.870 104.800 114.050 ;
        RECT 104.970 113.870 105.280 114.050 ;
        RECT 105.450 113.870 105.760 114.050 ;
        RECT 105.930 113.870 106.240 114.050 ;
        RECT 106.410 113.870 106.720 114.050 ;
        RECT 106.890 113.870 107.200 114.050 ;
        RECT 107.370 113.870 107.680 114.050 ;
        RECT 107.850 113.870 108.160 114.050 ;
        RECT 108.330 113.870 108.640 114.050 ;
        RECT 108.810 113.870 109.120 114.050 ;
        RECT 109.290 113.870 109.600 114.050 ;
        RECT 109.770 113.870 110.080 114.050 ;
        RECT 110.250 113.870 110.560 114.050 ;
        RECT 110.730 113.870 111.040 114.050 ;
        RECT 111.210 113.870 111.520 114.050 ;
        RECT 111.690 113.870 112.000 114.050 ;
        RECT 112.170 113.870 112.480 114.050 ;
        RECT 112.650 113.870 112.960 114.050 ;
        RECT 113.130 113.870 113.440 114.050 ;
        RECT 113.610 113.870 113.920 114.050 ;
        RECT 114.090 113.870 114.400 114.050 ;
        RECT 114.570 113.870 114.880 114.050 ;
        RECT 115.050 113.870 115.360 114.050 ;
        RECT 115.530 113.870 115.840 114.050 ;
        RECT 116.010 113.870 116.320 114.050 ;
        RECT 116.490 114.040 116.800 114.050 ;
        RECT 116.970 114.040 117.280 114.050 ;
        RECT 116.490 113.870 116.640 114.040 ;
        RECT 117.120 113.870 117.280 114.040 ;
        RECT 117.450 113.870 117.760 114.050 ;
        RECT 117.930 113.870 118.240 114.050 ;
        RECT 118.410 113.870 118.720 114.050 ;
        RECT 118.890 113.870 119.200 114.050 ;
        RECT 119.370 113.870 119.680 114.050 ;
        RECT 119.850 113.870 120.160 114.050 ;
        RECT 120.330 113.870 120.640 114.050 ;
        RECT 120.810 113.870 121.120 114.050 ;
        RECT 121.290 113.870 121.600 114.050 ;
        RECT 121.770 113.870 122.080 114.050 ;
        RECT 122.250 113.870 122.560 114.050 ;
        RECT 122.730 113.870 123.040 114.050 ;
        RECT 123.210 113.870 123.520 114.050 ;
        RECT 123.690 113.870 124.000 114.050 ;
        RECT 124.170 113.870 124.480 114.050 ;
        RECT 124.650 113.870 124.960 114.050 ;
        RECT 125.130 113.870 125.440 114.050 ;
        RECT 125.610 113.870 125.920 114.050 ;
        RECT 126.090 113.870 126.400 114.050 ;
        RECT 126.570 113.870 126.880 114.050 ;
        RECT 127.050 113.870 127.360 114.050 ;
        RECT 127.530 113.870 127.840 114.050 ;
        RECT 128.010 113.870 128.320 114.050 ;
        RECT 128.490 113.870 128.800 114.050 ;
        RECT 128.970 113.870 129.280 114.050 ;
        RECT 129.450 113.870 129.760 114.050 ;
        RECT 129.930 113.870 130.240 114.050 ;
        RECT 130.410 113.870 130.720 114.050 ;
        RECT 130.890 113.870 131.200 114.050 ;
        RECT 131.370 113.870 131.680 114.050 ;
        RECT 131.850 113.870 132.160 114.050 ;
        RECT 132.330 113.870 132.640 114.050 ;
        RECT 132.810 113.870 133.120 114.050 ;
        RECT 133.290 113.870 133.600 114.050 ;
        RECT 133.770 113.870 134.080 114.050 ;
        RECT 134.250 113.870 134.560 114.050 ;
        RECT 134.730 113.870 135.040 114.050 ;
        RECT 135.210 113.870 135.520 114.050 ;
        RECT 135.690 113.870 136.000 114.050 ;
        RECT 136.170 113.870 136.480 114.050 ;
        RECT 136.650 113.870 136.960 114.050 ;
        RECT 137.130 113.870 137.440 114.050 ;
        RECT 137.610 113.870 137.920 114.050 ;
        RECT 138.090 113.870 138.400 114.050 ;
        RECT 138.570 113.870 138.880 114.050 ;
        RECT 139.050 113.870 139.360 114.050 ;
        RECT 139.530 113.870 139.840 114.050 ;
        RECT 140.010 113.870 140.320 114.050 ;
        RECT 140.490 113.870 140.800 114.050 ;
        RECT 140.970 113.870 141.280 114.050 ;
        RECT 141.450 113.870 141.760 114.050 ;
        RECT 141.930 113.870 142.080 114.050 ;
        RECT 6.390 113.570 6.980 113.600 ;
        RECT 6.390 113.400 6.420 113.570 ;
        RECT 6.590 113.400 6.780 113.570 ;
        RECT 6.950 113.400 6.980 113.570 ;
        RECT 5.870 112.420 6.200 113.350 ;
        RECT 6.390 112.620 6.980 113.400 ;
        RECT 7.160 113.530 8.600 113.700 ;
        RECT 7.160 112.420 7.330 113.530 ;
        RECT 5.870 112.250 7.330 112.420 ;
        RECT 5.870 110.390 6.140 112.250 ;
        RECT 7.000 111.750 7.330 112.250 ;
        RECT 7.510 112.040 7.760 113.350 ;
        RECT 8.000 112.730 8.250 113.350 ;
        RECT 8.430 113.080 8.600 113.530 ;
        RECT 8.780 113.570 9.110 113.600 ;
        RECT 8.780 113.400 8.810 113.570 ;
        RECT 8.980 113.400 9.110 113.570 ;
        RECT 8.780 113.260 9.110 113.400 ;
        RECT 9.290 113.530 11.030 113.700 ;
        RECT 9.290 113.080 9.460 113.530 ;
        RECT 8.430 112.910 9.460 113.080 ;
        RECT 9.640 112.730 9.810 113.350 ;
        RECT 10.340 113.090 10.670 113.350 ;
        RECT 8.000 112.560 9.810 112.730 ;
        RECT 9.990 112.560 10.210 112.890 ;
        RECT 9.640 112.380 9.810 112.560 ;
        RECT 7.510 111.810 8.040 112.040 ;
        RECT 7.510 110.890 7.780 111.810 ;
      LAYER li1 ;
        RECT 8.460 111.510 9.000 112.380 ;
      LAYER li1 ;
        RECT 9.640 112.210 9.860 112.380 ;
        RECT 6.320 110.260 7.270 110.890 ;
        RECT 7.450 110.390 7.780 110.890 ;
        RECT 7.960 110.260 8.550 111.140 ;
      LAYER li1 ;
        RECT 8.830 110.520 9.000 111.510 ;
        RECT 9.180 110.700 9.510 112.000 ;
      LAYER li1 ;
        RECT 9.690 111.220 9.860 112.210 ;
        RECT 10.040 112.040 10.210 112.560 ;
        RECT 10.390 112.390 10.560 113.090 ;
        RECT 10.860 112.940 11.030 113.530 ;
        RECT 11.210 113.570 12.160 113.600 ;
        RECT 11.210 113.400 11.240 113.570 ;
        RECT 11.410 113.400 11.600 113.570 ;
        RECT 11.770 113.400 11.960 113.570 ;
        RECT 12.130 113.400 12.160 113.570 ;
        RECT 11.210 113.120 12.160 113.400 ;
        RECT 12.340 113.530 13.370 113.700 ;
        RECT 12.340 112.940 12.510 113.530 ;
        RECT 10.860 112.890 12.510 112.940 ;
        RECT 10.740 112.770 12.510 112.890 ;
        RECT 10.740 112.570 11.070 112.770 ;
        RECT 12.690 112.590 13.020 113.350 ;
        RECT 13.200 113.170 13.370 113.530 ;
        RECT 13.550 113.570 14.500 113.650 ;
        RECT 13.550 113.400 13.580 113.570 ;
        RECT 13.750 113.400 13.940 113.570 ;
        RECT 14.110 113.400 14.300 113.570 ;
        RECT 14.470 113.400 14.500 113.570 ;
        RECT 13.550 113.350 14.500 113.400 ;
        RECT 13.200 113.000 15.010 113.170 ;
        RECT 11.250 112.420 13.020 112.590 ;
        RECT 11.250 112.390 11.420 112.420 ;
        RECT 10.390 112.220 11.420 112.390 ;
        RECT 14.330 112.240 14.660 112.820 ;
        RECT 10.040 111.810 11.070 112.040 ;
        RECT 10.740 111.320 11.070 111.810 ;
        RECT 11.250 111.540 11.420 112.220 ;
        RECT 11.600 112.070 14.660 112.240 ;
        RECT 11.600 111.720 11.930 112.070 ;
      LAYER li1 ;
        RECT 12.370 111.720 14.220 111.890 ;
      LAYER li1 ;
        RECT 11.250 111.370 13.870 111.540 ;
        RECT 9.690 110.720 9.960 111.220 ;
        RECT 11.250 111.140 11.420 111.370 ;
      LAYER li1 ;
        RECT 14.050 111.190 14.220 111.720 ;
      LAYER li1 ;
        RECT 10.410 110.970 11.420 111.140 ;
      LAYER li1 ;
        RECT 11.600 111.020 14.220 111.190 ;
      LAYER li1 ;
        RECT 10.410 110.720 10.740 110.970 ;
      LAYER li1 ;
        RECT 11.600 110.520 11.770 111.020 ;
        RECT 8.830 110.350 11.770 110.520 ;
      LAYER li1 ;
        RECT 12.920 110.260 13.870 110.840 ;
      LAYER li1 ;
        RECT 14.050 110.330 14.220 111.020 ;
      LAYER li1 ;
        RECT 14.400 111.220 14.660 112.070 ;
        RECT 14.840 111.650 15.010 113.000 ;
        RECT 15.190 112.740 15.440 113.650 ;
        RECT 16.250 113.570 17.200 113.600 ;
        RECT 18.030 113.570 18.930 113.600 ;
        RECT 16.250 113.400 16.280 113.570 ;
        RECT 16.450 113.400 16.640 113.570 ;
        RECT 16.810 113.400 17.000 113.570 ;
        RECT 17.170 113.400 17.200 113.570 ;
        RECT 18.200 113.400 18.390 113.570 ;
        RECT 18.560 113.400 18.750 113.570 ;
        RECT 18.920 113.400 18.930 113.570 ;
        RECT 15.190 112.570 16.070 112.740 ;
        RECT 16.250 112.570 17.200 113.400 ;
        RECT 17.600 112.600 17.850 113.070 ;
        RECT 18.030 112.780 18.930 113.400 ;
        RECT 19.540 113.570 20.480 113.630 ;
        RECT 19.540 113.400 19.560 113.570 ;
        RECT 19.730 113.400 19.920 113.570 ;
        RECT 20.090 113.400 20.280 113.570 ;
        RECT 20.450 113.400 20.480 113.570 ;
        RECT 15.390 111.830 15.720 112.330 ;
        RECT 15.900 112.250 16.070 112.570 ;
        RECT 17.600 112.430 18.610 112.600 ;
        RECT 15.900 112.080 18.260 112.250 ;
        RECT 14.840 111.480 16.010 111.650 ;
        RECT 14.400 110.510 14.730 111.220 ;
        RECT 15.190 110.680 15.520 111.220 ;
        RECT 15.730 110.980 16.010 111.480 ;
        RECT 16.190 110.680 16.360 112.080 ;
        RECT 18.440 111.900 18.610 112.430 ;
        RECT 16.570 111.730 18.610 111.900 ;
        RECT 16.570 111.340 16.900 111.730 ;
      LAYER li1 ;
        RECT 17.220 111.160 17.550 111.550 ;
      LAYER li1 ;
        RECT 15.190 110.510 16.360 110.680 ;
      LAYER li1 ;
        RECT 16.540 110.990 17.550 111.160 ;
        RECT 16.540 110.330 16.710 110.990 ;
      LAYER li1 ;
        RECT 18.380 110.890 18.610 111.730 ;
        RECT 19.110 111.900 19.360 112.900 ;
        RECT 19.540 112.090 20.480 113.400 ;
        RECT 19.110 111.570 20.480 111.900 ;
        RECT 19.110 111.390 19.320 111.570 ;
        RECT 18.990 110.890 19.320 111.390 ;
      LAYER li1 ;
        RECT 14.050 110.160 16.710 110.330 ;
      LAYER li1 ;
        RECT 16.890 110.260 17.840 110.810 ;
        RECT 18.380 110.390 18.710 110.890 ;
        RECT 19.500 110.260 20.450 111.390 ;
      LAYER li1 ;
        RECT 20.660 110.560 21.000 113.630 ;
      LAYER li1 ;
        RECT 21.370 113.620 22.820 113.650 ;
        RECT 21.370 113.450 21.620 113.620 ;
        RECT 21.790 113.450 21.980 113.620 ;
        RECT 22.150 113.450 22.420 113.620 ;
        RECT 22.590 113.450 22.820 113.620 ;
        RECT 21.370 112.580 22.820 113.450 ;
        RECT 24.570 113.570 25.830 113.650 ;
        RECT 24.570 113.400 24.580 113.570 ;
        RECT 24.750 113.400 24.940 113.570 ;
        RECT 25.110 113.400 25.300 113.570 ;
        RECT 25.470 113.400 25.660 113.570 ;
        RECT 21.600 111.140 21.930 111.920 ;
        RECT 22.140 111.590 22.470 112.580 ;
        RECT 24.570 112.170 25.830 113.400 ;
      LAYER li1 ;
        RECT 26.360 113.150 26.530 113.650 ;
        RECT 26.010 112.070 26.530 113.150 ;
      LAYER li1 ;
        RECT 26.790 113.570 28.100 113.650 ;
        RECT 26.790 113.400 26.820 113.570 ;
        RECT 26.990 113.400 27.180 113.570 ;
        RECT 27.350 113.400 27.540 113.570 ;
        RECT 27.710 113.400 27.900 113.570 ;
        RECT 28.070 113.400 28.100 113.570 ;
        RECT 26.790 112.190 28.100 113.400 ;
        RECT 28.820 113.620 31.560 113.640 ;
        RECT 28.820 113.450 29.030 113.620 ;
        RECT 29.200 113.450 29.470 113.620 ;
        RECT 29.640 113.450 29.880 113.620 ;
        RECT 30.050 113.450 30.310 113.620 ;
        RECT 30.480 113.450 30.750 113.620 ;
        RECT 30.920 113.450 31.160 113.620 ;
        RECT 31.330 113.450 31.560 113.620 ;
        RECT 28.820 112.570 31.560 113.450 ;
        RECT 32.660 113.620 35.400 113.640 ;
        RECT 32.660 113.450 32.870 113.620 ;
        RECT 33.040 113.450 33.310 113.620 ;
        RECT 33.480 113.450 33.720 113.620 ;
        RECT 33.890 113.450 34.150 113.620 ;
        RECT 34.320 113.450 34.590 113.620 ;
        RECT 34.760 113.450 35.000 113.620 ;
        RECT 35.170 113.450 35.400 113.620 ;
        RECT 32.660 112.570 35.400 113.450 ;
      LAYER li1 ;
        RECT 26.010 111.990 26.280 112.070 ;
        RECT 25.220 111.820 26.280 111.990 ;
        RECT 24.610 111.430 25.030 111.760 ;
        RECT 25.220 111.250 25.390 111.820 ;
        RECT 26.730 111.700 27.240 112.010 ;
        RECT 27.490 111.700 28.200 112.010 ;
        RECT 25.570 111.430 26.080 111.640 ;
      LAYER li1 ;
        RECT 26.280 111.350 28.150 111.520 ;
        RECT 21.600 110.740 22.900 111.140 ;
        RECT 21.290 110.260 22.900 110.740 ;
        RECT 24.640 110.330 24.970 111.250 ;
      LAYER li1 ;
        RECT 25.220 110.900 25.750 111.250 ;
        RECT 25.220 110.730 25.760 110.900 ;
        RECT 25.220 110.510 25.750 110.730 ;
      LAYER li1 ;
        RECT 26.280 110.330 26.450 111.350 ;
        RECT 24.640 110.160 26.450 110.330 ;
        RECT 26.630 110.260 27.730 111.170 ;
        RECT 27.900 110.420 28.150 111.350 ;
        RECT 29.060 111.250 29.390 111.920 ;
        RECT 29.790 111.590 30.120 112.570 ;
        RECT 30.340 111.250 30.670 111.920 ;
        RECT 31.070 111.590 31.400 112.570 ;
        RECT 32.900 111.250 33.230 111.920 ;
        RECT 33.630 111.590 33.960 112.570 ;
        RECT 34.180 111.250 34.510 111.920 ;
        RECT 34.910 111.590 35.240 112.570 ;
      LAYER li1 ;
        RECT 37.560 112.070 37.990 113.650 ;
      LAYER li1 ;
        RECT 38.170 113.570 38.730 113.650 ;
        RECT 38.170 113.400 38.180 113.570 ;
        RECT 38.350 113.400 38.540 113.570 ;
        RECT 38.710 113.400 38.730 113.570 ;
        RECT 38.170 112.070 38.730 113.400 ;
        RECT 40.090 113.620 41.540 113.650 ;
        RECT 40.090 113.450 40.340 113.620 ;
        RECT 40.510 113.450 40.700 113.620 ;
        RECT 40.870 113.450 41.140 113.620 ;
        RECT 41.310 113.450 41.540 113.620 ;
        RECT 28.900 110.250 31.630 111.250 ;
        RECT 32.740 110.250 35.470 111.250 ;
      LAYER li1 ;
        RECT 37.560 110.390 37.810 112.070 ;
      LAYER li1 ;
        RECT 38.120 111.180 38.450 111.640 ;
      LAYER li1 ;
        RECT 38.910 111.360 39.240 113.150 ;
      LAYER li1 ;
        RECT 39.420 111.180 39.670 112.900 ;
        RECT 40.090 112.580 41.540 113.450 ;
        RECT 41.850 113.570 42.800 113.650 ;
        RECT 41.850 113.400 41.880 113.570 ;
        RECT 42.050 113.400 42.240 113.570 ;
        RECT 42.410 113.400 42.600 113.570 ;
        RECT 42.770 113.400 42.800 113.570 ;
        RECT 38.120 111.010 39.670 111.180 ;
        RECT 37.990 110.260 39.240 110.830 ;
        RECT 39.420 110.390 39.670 111.010 ;
        RECT 40.320 111.140 40.650 111.920 ;
        RECT 40.860 111.590 41.190 112.580 ;
        RECT 41.850 112.070 42.800 113.400 ;
      LAYER li1 ;
        RECT 42.980 111.970 43.230 113.650 ;
      LAYER li1 ;
        RECT 43.410 113.570 44.360 113.650 ;
        RECT 43.410 113.400 43.440 113.570 ;
        RECT 43.610 113.400 43.800 113.570 ;
        RECT 43.970 113.400 44.160 113.570 ;
        RECT 44.330 113.400 44.360 113.570 ;
        RECT 43.410 112.150 44.360 113.400 ;
      LAYER li1 ;
        RECT 44.540 111.970 44.870 113.650 ;
      LAYER li1 ;
        RECT 45.050 113.570 46.000 113.650 ;
        RECT 45.050 113.400 45.080 113.570 ;
        RECT 45.250 113.400 45.440 113.570 ;
        RECT 45.610 113.400 45.800 113.570 ;
        RECT 45.970 113.400 46.000 113.570 ;
        RECT 45.050 112.190 46.000 113.400 ;
      LAYER li1 ;
        RECT 42.980 111.800 44.870 111.970 ;
        RECT 42.980 111.670 43.150 111.800 ;
        RECT 45.650 111.670 45.980 112.010 ;
        RECT 41.890 111.440 43.150 111.670 ;
      LAYER li1 ;
        RECT 43.330 111.490 45.360 111.620 ;
        RECT 46.180 111.490 46.430 113.650 ;
        RECT 46.810 113.620 48.260 113.650 ;
        RECT 46.810 113.450 47.060 113.620 ;
        RECT 47.230 113.450 47.420 113.620 ;
        RECT 47.590 113.450 47.860 113.620 ;
        RECT 48.030 113.450 48.260 113.620 ;
        RECT 46.810 112.580 48.260 113.450 ;
        RECT 48.570 113.570 49.520 113.650 ;
        RECT 48.570 113.400 48.600 113.570 ;
        RECT 48.770 113.400 48.960 113.570 ;
        RECT 49.130 113.400 49.320 113.570 ;
        RECT 49.490 113.400 49.520 113.570 ;
        RECT 43.330 111.450 46.430 111.490 ;
      LAYER li1 ;
        RECT 42.980 111.270 43.150 111.440 ;
      LAYER li1 ;
        RECT 45.190 111.320 46.430 111.450 ;
        RECT 40.320 110.740 41.620 111.140 ;
        RECT 40.010 110.260 41.620 110.740 ;
        RECT 41.850 110.260 42.800 111.220 ;
      LAYER li1 ;
        RECT 42.980 111.100 44.790 111.270 ;
        RECT 42.980 110.390 43.230 111.100 ;
      LAYER li1 ;
        RECT 43.410 110.260 44.360 110.920 ;
      LAYER li1 ;
        RECT 44.540 110.390 44.790 111.100 ;
      LAYER li1 ;
        RECT 44.970 110.260 45.920 111.140 ;
        RECT 46.100 110.390 46.430 111.320 ;
        RECT 47.040 111.140 47.370 111.920 ;
        RECT 47.580 111.590 47.910 112.580 ;
        RECT 48.570 112.070 49.520 113.400 ;
      LAYER li1 ;
        RECT 49.700 111.970 49.950 113.650 ;
      LAYER li1 ;
        RECT 50.130 113.570 51.080 113.650 ;
        RECT 50.130 113.400 50.160 113.570 ;
        RECT 50.330 113.400 50.520 113.570 ;
        RECT 50.690 113.400 50.880 113.570 ;
        RECT 51.050 113.400 51.080 113.570 ;
        RECT 50.130 112.150 51.080 113.400 ;
      LAYER li1 ;
        RECT 51.260 111.970 51.590 113.650 ;
      LAYER li1 ;
        RECT 51.770 113.570 52.720 113.650 ;
        RECT 51.770 113.400 51.800 113.570 ;
        RECT 51.970 113.400 52.160 113.570 ;
        RECT 52.330 113.400 52.520 113.570 ;
        RECT 52.690 113.400 52.720 113.570 ;
        RECT 51.770 112.190 52.720 113.400 ;
      LAYER li1 ;
        RECT 49.700 111.800 51.590 111.970 ;
        RECT 49.700 111.670 49.870 111.800 ;
        RECT 52.370 111.670 52.700 112.010 ;
        RECT 48.610 111.440 49.870 111.670 ;
      LAYER li1 ;
        RECT 50.050 111.490 52.080 111.620 ;
        RECT 52.900 111.490 53.150 113.650 ;
        RECT 53.530 113.620 54.980 113.650 ;
        RECT 53.530 113.450 53.780 113.620 ;
        RECT 53.950 113.450 54.140 113.620 ;
        RECT 54.310 113.450 54.580 113.620 ;
        RECT 54.750 113.450 54.980 113.620 ;
        RECT 53.530 112.580 54.980 113.450 ;
        RECT 55.290 113.570 56.240 113.650 ;
        RECT 55.290 113.400 55.320 113.570 ;
        RECT 55.490 113.400 55.680 113.570 ;
        RECT 55.850 113.400 56.040 113.570 ;
        RECT 56.210 113.400 56.240 113.570 ;
        RECT 50.050 111.450 53.150 111.490 ;
      LAYER li1 ;
        RECT 49.700 111.270 49.870 111.440 ;
      LAYER li1 ;
        RECT 51.910 111.320 53.150 111.450 ;
        RECT 47.040 110.740 48.340 111.140 ;
        RECT 46.730 110.260 48.340 110.740 ;
        RECT 48.570 110.260 49.520 111.220 ;
      LAYER li1 ;
        RECT 49.700 111.100 51.510 111.270 ;
        RECT 49.700 110.390 49.950 111.100 ;
      LAYER li1 ;
        RECT 50.130 110.260 51.080 110.920 ;
      LAYER li1 ;
        RECT 51.260 110.390 51.510 111.100 ;
      LAYER li1 ;
        RECT 51.690 110.260 52.640 111.140 ;
        RECT 52.820 110.390 53.150 111.320 ;
        RECT 53.760 111.140 54.090 111.920 ;
        RECT 54.300 111.590 54.630 112.580 ;
        RECT 55.290 112.070 56.240 113.400 ;
      LAYER li1 ;
        RECT 56.420 111.970 56.670 113.650 ;
      LAYER li1 ;
        RECT 56.850 113.570 57.800 113.650 ;
        RECT 56.850 113.400 56.880 113.570 ;
        RECT 57.050 113.400 57.240 113.570 ;
        RECT 57.410 113.400 57.600 113.570 ;
        RECT 57.770 113.400 57.800 113.570 ;
        RECT 56.850 112.150 57.800 113.400 ;
      LAYER li1 ;
        RECT 57.980 111.970 58.310 113.650 ;
      LAYER li1 ;
        RECT 58.490 113.570 59.440 113.650 ;
        RECT 58.490 113.400 58.520 113.570 ;
        RECT 58.690 113.400 58.880 113.570 ;
        RECT 59.050 113.400 59.240 113.570 ;
        RECT 59.410 113.400 59.440 113.570 ;
        RECT 58.490 112.190 59.440 113.400 ;
      LAYER li1 ;
        RECT 56.420 111.800 58.310 111.970 ;
        RECT 56.420 111.670 56.590 111.800 ;
        RECT 59.090 111.670 59.420 112.010 ;
        RECT 55.330 111.440 56.590 111.670 ;
      LAYER li1 ;
        RECT 56.770 111.490 58.800 111.620 ;
        RECT 59.620 111.490 59.870 113.650 ;
        RECT 60.250 113.620 61.700 113.650 ;
        RECT 60.250 113.450 60.500 113.620 ;
        RECT 60.670 113.450 60.860 113.620 ;
        RECT 61.030 113.450 61.300 113.620 ;
        RECT 61.470 113.450 61.700 113.620 ;
        RECT 60.250 112.580 61.700 113.450 ;
        RECT 62.970 113.570 63.920 113.650 ;
        RECT 62.970 113.400 63.000 113.570 ;
        RECT 63.170 113.400 63.360 113.570 ;
        RECT 63.530 113.400 63.720 113.570 ;
        RECT 63.890 113.400 63.920 113.570 ;
        RECT 56.770 111.450 59.870 111.490 ;
      LAYER li1 ;
        RECT 56.420 111.270 56.590 111.440 ;
      LAYER li1 ;
        RECT 58.630 111.320 59.870 111.450 ;
        RECT 53.760 110.740 55.060 111.140 ;
        RECT 53.450 110.260 55.060 110.740 ;
        RECT 55.290 110.260 56.240 111.220 ;
      LAYER li1 ;
        RECT 56.420 111.100 58.230 111.270 ;
        RECT 56.420 110.390 56.670 111.100 ;
      LAYER li1 ;
        RECT 56.850 110.260 57.800 110.920 ;
      LAYER li1 ;
        RECT 57.980 110.390 58.230 111.100 ;
      LAYER li1 ;
        RECT 58.410 110.260 59.360 111.140 ;
        RECT 59.540 110.390 59.870 111.320 ;
        RECT 60.480 111.140 60.810 111.920 ;
        RECT 61.020 111.590 61.350 112.580 ;
        RECT 62.970 112.070 63.920 113.400 ;
      LAYER li1 ;
        RECT 64.100 111.970 64.350 113.650 ;
      LAYER li1 ;
        RECT 64.530 113.570 65.480 113.650 ;
        RECT 64.530 113.400 64.560 113.570 ;
        RECT 64.730 113.400 64.920 113.570 ;
        RECT 65.090 113.400 65.280 113.570 ;
        RECT 65.450 113.400 65.480 113.570 ;
        RECT 64.530 112.150 65.480 113.400 ;
      LAYER li1 ;
        RECT 65.660 111.970 65.990 113.650 ;
      LAYER li1 ;
        RECT 66.170 113.570 67.120 113.650 ;
        RECT 66.170 113.400 66.200 113.570 ;
        RECT 66.370 113.400 66.560 113.570 ;
        RECT 66.730 113.400 66.920 113.570 ;
        RECT 67.090 113.400 67.120 113.570 ;
        RECT 66.170 112.190 67.120 113.400 ;
      LAYER li1 ;
        RECT 64.100 111.800 65.990 111.970 ;
        RECT 64.100 111.670 64.270 111.800 ;
        RECT 66.770 111.670 67.100 112.010 ;
        RECT 63.010 111.440 64.270 111.670 ;
      LAYER li1 ;
        RECT 64.450 111.490 66.480 111.620 ;
        RECT 67.300 111.490 67.550 113.650 ;
        RECT 68.180 113.620 70.920 113.640 ;
        RECT 68.180 113.450 68.390 113.620 ;
        RECT 68.560 113.450 68.830 113.620 ;
        RECT 69.000 113.450 69.240 113.620 ;
        RECT 69.410 113.450 69.670 113.620 ;
        RECT 69.840 113.450 70.110 113.620 ;
        RECT 70.280 113.450 70.520 113.620 ;
        RECT 70.690 113.450 70.920 113.620 ;
        RECT 68.180 112.570 70.920 113.450 ;
        RECT 64.450 111.450 67.550 111.490 ;
      LAYER li1 ;
        RECT 64.100 111.270 64.270 111.440 ;
      LAYER li1 ;
        RECT 66.310 111.320 67.550 111.450 ;
        RECT 60.480 110.740 61.780 111.140 ;
        RECT 60.170 110.260 61.780 110.740 ;
        RECT 62.970 110.260 63.920 111.220 ;
      LAYER li1 ;
        RECT 64.100 111.100 65.910 111.270 ;
        RECT 64.100 110.390 64.350 111.100 ;
      LAYER li1 ;
        RECT 64.530 110.260 65.480 110.920 ;
      LAYER li1 ;
        RECT 65.660 110.390 65.910 111.100 ;
      LAYER li1 ;
        RECT 66.090 110.260 67.040 111.140 ;
        RECT 67.220 110.390 67.550 111.320 ;
        RECT 68.420 111.250 68.750 111.920 ;
        RECT 69.150 111.590 69.480 112.570 ;
        RECT 69.700 111.250 70.030 111.920 ;
        RECT 70.430 111.590 70.760 112.570 ;
      LAYER li1 ;
        RECT 72.120 112.070 72.550 113.650 ;
      LAYER li1 ;
        RECT 72.730 113.570 73.290 113.650 ;
        RECT 72.730 113.400 72.740 113.570 ;
        RECT 72.910 113.400 73.100 113.570 ;
        RECT 73.270 113.400 73.290 113.570 ;
        RECT 72.730 112.070 73.290 113.400 ;
        RECT 74.650 113.620 76.100 113.650 ;
        RECT 74.650 113.450 74.900 113.620 ;
        RECT 75.070 113.450 75.260 113.620 ;
        RECT 75.430 113.450 75.700 113.620 ;
        RECT 75.870 113.450 76.100 113.620 ;
        RECT 68.260 110.250 70.990 111.250 ;
      LAYER li1 ;
        RECT 72.120 110.390 72.370 112.070 ;
      LAYER li1 ;
        RECT 72.680 111.180 73.010 111.640 ;
      LAYER li1 ;
        RECT 73.470 111.360 73.800 113.150 ;
      LAYER li1 ;
        RECT 73.980 111.180 74.230 112.900 ;
        RECT 74.650 112.580 76.100 113.450 ;
        RECT 77.370 113.570 78.320 113.650 ;
        RECT 77.370 113.400 77.400 113.570 ;
        RECT 77.570 113.400 77.760 113.570 ;
        RECT 77.930 113.400 78.120 113.570 ;
        RECT 78.290 113.400 78.320 113.570 ;
        RECT 72.680 111.010 74.230 111.180 ;
        RECT 72.550 110.260 73.800 110.830 ;
        RECT 73.980 110.390 74.230 111.010 ;
        RECT 74.880 111.140 75.210 111.920 ;
        RECT 75.420 111.590 75.750 112.580 ;
        RECT 77.370 112.070 78.320 113.400 ;
      LAYER li1 ;
        RECT 78.850 112.000 79.320 113.650 ;
      LAYER li1 ;
        RECT 79.500 113.570 80.450 113.650 ;
        RECT 79.500 113.400 79.530 113.570 ;
        RECT 79.700 113.400 79.890 113.570 ;
        RECT 80.060 113.400 80.250 113.570 ;
        RECT 80.420 113.400 80.450 113.570 ;
        RECT 79.500 112.190 80.450 113.400 ;
        RECT 80.890 113.620 82.340 113.650 ;
        RECT 80.890 113.450 81.140 113.620 ;
        RECT 81.310 113.450 81.500 113.620 ;
        RECT 81.670 113.450 81.940 113.620 ;
        RECT 82.110 113.450 82.340 113.620 ;
        RECT 80.890 112.580 82.340 113.450 ;
      LAYER li1 ;
        RECT 78.850 111.830 79.430 112.000 ;
        RECT 78.350 111.400 79.080 111.650 ;
        RECT 79.260 111.520 79.430 111.830 ;
        RECT 79.610 111.700 80.520 112.010 ;
        RECT 79.260 111.350 80.100 111.520 ;
      LAYER li1 ;
        RECT 77.410 111.170 77.740 111.220 ;
        RECT 74.880 110.740 76.180 111.140 ;
        RECT 74.570 110.260 76.180 110.740 ;
        RECT 77.410 111.000 79.320 111.170 ;
        RECT 77.410 110.390 77.740 111.000 ;
        RECT 77.920 110.260 78.810 110.820 ;
        RECT 78.990 110.390 79.320 111.000 ;
      LAYER li1 ;
        RECT 79.770 110.390 80.100 111.350 ;
      LAYER li1 ;
        RECT 81.120 111.140 81.450 111.920 ;
        RECT 81.660 111.590 81.990 112.580 ;
        RECT 81.120 110.740 82.420 111.140 ;
        RECT 80.810 110.260 82.420 110.740 ;
      LAYER li1 ;
        RECT 82.690 110.390 82.940 113.650 ;
      LAYER li1 ;
        RECT 83.120 113.570 85.810 113.650 ;
        RECT 83.290 113.400 83.480 113.570 ;
        RECT 83.650 113.400 83.840 113.570 ;
        RECT 84.010 113.400 84.200 113.570 ;
        RECT 84.370 113.400 84.560 113.570 ;
        RECT 84.730 113.400 84.920 113.570 ;
        RECT 85.090 113.400 85.280 113.570 ;
        RECT 85.450 113.400 85.640 113.570 ;
        RECT 83.120 112.540 85.810 113.400 ;
        RECT 85.990 112.360 86.240 113.650 ;
        RECT 83.150 112.190 86.240 112.360 ;
        RECT 83.150 111.490 83.480 112.190 ;
        RECT 85.990 112.070 86.240 112.190 ;
        RECT 86.420 113.570 87.730 113.630 ;
        RECT 86.420 113.400 86.450 113.570 ;
        RECT 86.620 113.400 86.810 113.570 ;
        RECT 86.980 113.400 87.170 113.570 ;
        RECT 87.340 113.400 87.530 113.570 ;
        RECT 87.700 113.400 87.730 113.570 ;
        RECT 86.420 112.090 87.730 113.400 ;
        RECT 88.090 113.620 89.540 113.650 ;
        RECT 88.090 113.450 88.340 113.620 ;
        RECT 88.510 113.450 88.700 113.620 ;
        RECT 88.870 113.450 89.140 113.620 ;
        RECT 89.310 113.450 89.540 113.620 ;
        RECT 88.090 112.580 89.540 113.450 ;
      LAYER li1 ;
        RECT 83.980 111.670 84.710 111.950 ;
      LAYER li1 ;
        RECT 83.150 111.320 84.360 111.490 ;
        RECT 83.120 110.260 84.010 111.140 ;
        RECT 84.190 111.110 84.360 111.320 ;
      LAYER li1 ;
        RECT 84.540 111.460 84.710 111.670 ;
        RECT 84.890 111.640 85.320 112.010 ;
        RECT 85.520 111.470 85.810 112.010 ;
        RECT 86.050 111.470 86.760 111.800 ;
        RECT 87.110 111.640 87.440 111.910 ;
        RECT 87.030 111.470 87.440 111.640 ;
        RECT 84.540 111.290 85.340 111.460 ;
        RECT 87.110 111.290 87.440 111.470 ;
        RECT 85.170 111.120 87.440 111.290 ;
      LAYER li1 ;
        RECT 88.320 111.140 88.650 111.920 ;
        RECT 88.860 111.590 89.190 112.580 ;
      LAYER li1 ;
        RECT 89.870 111.220 90.120 113.630 ;
      LAYER li1 ;
        RECT 90.300 113.570 91.200 113.650 ;
        RECT 90.300 113.400 90.310 113.570 ;
        RECT 90.480 113.400 90.670 113.570 ;
        RECT 90.840 113.400 91.030 113.570 ;
        RECT 90.300 112.170 91.200 113.400 ;
        RECT 91.380 111.990 91.630 113.650 ;
        RECT 92.080 112.340 92.410 113.650 ;
        RECT 92.590 113.570 93.540 113.650 ;
        RECT 92.590 113.400 92.620 113.570 ;
        RECT 92.790 113.400 92.980 113.570 ;
        RECT 93.150 113.400 93.340 113.570 ;
        RECT 93.510 113.400 93.540 113.570 ;
        RECT 92.590 112.520 93.540 113.400 ;
        RECT 93.720 112.340 93.970 113.630 ;
        RECT 94.330 113.620 95.780 113.650 ;
        RECT 94.330 113.450 94.580 113.620 ;
        RECT 94.750 113.450 94.940 113.620 ;
        RECT 95.110 113.450 95.380 113.620 ;
        RECT 95.550 113.450 95.780 113.620 ;
        RECT 94.330 112.580 95.780 113.450 ;
        RECT 96.090 113.570 97.040 113.650 ;
        RECT 96.090 113.400 96.120 113.570 ;
        RECT 96.290 113.400 96.480 113.570 ;
        RECT 96.650 113.400 96.840 113.570 ;
        RECT 97.010 113.400 97.040 113.570 ;
        RECT 92.080 112.170 93.970 112.340 ;
        RECT 93.720 112.090 93.970 112.170 ;
        RECT 90.330 111.820 92.390 111.990 ;
        RECT 90.330 111.620 90.660 111.820 ;
      LAYER li1 ;
        RECT 90.850 111.400 92.040 111.640 ;
      LAYER li1 ;
        RECT 92.220 111.220 92.390 111.820 ;
      LAYER li1 ;
        RECT 93.660 111.400 93.960 111.730 ;
      LAYER li1 ;
        RECT 84.190 110.940 84.990 111.110 ;
      LAYER li1 ;
        RECT 85.600 111.100 86.270 111.120 ;
      LAYER li1 ;
        RECT 84.820 110.770 85.420 110.940 ;
        RECT 84.310 110.330 84.640 110.760 ;
        RECT 85.090 110.510 85.420 110.770 ;
        RECT 85.910 110.330 86.240 110.920 ;
        RECT 84.310 110.160 86.240 110.330 ;
        RECT 86.450 110.260 87.750 110.940 ;
        RECT 88.320 110.740 89.620 111.140 ;
        RECT 88.010 110.260 89.620 110.740 ;
      LAYER li1 ;
        RECT 89.870 110.390 90.220 111.220 ;
      LAYER li1 ;
        RECT 90.400 110.260 92.010 111.220 ;
        RECT 92.190 110.390 92.440 111.220 ;
        RECT 92.620 110.260 93.930 111.220 ;
        RECT 94.560 111.140 94.890 111.920 ;
        RECT 95.100 111.590 95.430 112.580 ;
        RECT 96.090 112.070 97.040 113.400 ;
      LAYER li1 ;
        RECT 97.220 111.970 97.470 113.650 ;
      LAYER li1 ;
        RECT 97.650 113.570 98.600 113.650 ;
        RECT 97.650 113.400 97.680 113.570 ;
        RECT 97.850 113.400 98.040 113.570 ;
        RECT 98.210 113.400 98.400 113.570 ;
        RECT 98.570 113.400 98.600 113.570 ;
        RECT 97.650 112.150 98.600 113.400 ;
      LAYER li1 ;
        RECT 98.780 111.970 99.110 113.650 ;
      LAYER li1 ;
        RECT 99.290 113.570 100.240 113.650 ;
        RECT 99.290 113.400 99.320 113.570 ;
        RECT 99.490 113.400 99.680 113.570 ;
        RECT 99.850 113.400 100.040 113.570 ;
        RECT 100.210 113.400 100.240 113.570 ;
        RECT 99.290 112.190 100.240 113.400 ;
      LAYER li1 ;
        RECT 97.220 111.800 99.110 111.970 ;
        RECT 97.220 111.670 97.390 111.800 ;
        RECT 99.890 111.670 100.220 112.010 ;
        RECT 96.130 111.440 97.390 111.670 ;
      LAYER li1 ;
        RECT 97.570 111.490 99.600 111.620 ;
        RECT 100.420 111.490 100.670 113.650 ;
        RECT 101.050 113.620 102.500 113.650 ;
        RECT 101.050 113.450 101.300 113.620 ;
        RECT 101.470 113.450 101.660 113.620 ;
        RECT 101.830 113.450 102.100 113.620 ;
        RECT 102.270 113.450 102.500 113.620 ;
        RECT 101.050 112.580 102.500 113.450 ;
        RECT 102.810 113.570 103.760 113.650 ;
        RECT 102.810 113.400 102.840 113.570 ;
        RECT 103.010 113.400 103.200 113.570 ;
        RECT 103.370 113.400 103.560 113.570 ;
        RECT 103.730 113.400 103.760 113.570 ;
        RECT 97.570 111.450 100.670 111.490 ;
      LAYER li1 ;
        RECT 97.220 111.270 97.390 111.440 ;
      LAYER li1 ;
        RECT 99.430 111.320 100.670 111.450 ;
        RECT 94.560 110.740 95.860 111.140 ;
        RECT 94.250 110.260 95.860 110.740 ;
        RECT 96.090 110.260 97.040 111.220 ;
      LAYER li1 ;
        RECT 97.220 111.100 99.030 111.270 ;
        RECT 97.220 110.390 97.470 111.100 ;
      LAYER li1 ;
        RECT 97.650 110.260 98.600 110.920 ;
      LAYER li1 ;
        RECT 98.780 110.390 99.030 111.100 ;
      LAYER li1 ;
        RECT 99.210 110.260 100.160 111.140 ;
        RECT 100.340 110.390 100.670 111.320 ;
        RECT 101.280 111.140 101.610 111.920 ;
        RECT 101.820 111.590 102.150 112.580 ;
        RECT 102.810 112.070 103.760 113.400 ;
      LAYER li1 ;
        RECT 103.940 111.970 104.190 113.650 ;
      LAYER li1 ;
        RECT 104.370 113.570 105.320 113.650 ;
        RECT 104.370 113.400 104.400 113.570 ;
        RECT 104.570 113.400 104.760 113.570 ;
        RECT 104.930 113.400 105.120 113.570 ;
        RECT 105.290 113.400 105.320 113.570 ;
        RECT 104.370 112.150 105.320 113.400 ;
      LAYER li1 ;
        RECT 105.500 111.970 105.830 113.650 ;
      LAYER li1 ;
        RECT 106.010 113.570 106.960 113.650 ;
        RECT 106.010 113.400 106.040 113.570 ;
        RECT 106.210 113.400 106.400 113.570 ;
        RECT 106.570 113.400 106.760 113.570 ;
        RECT 106.930 113.400 106.960 113.570 ;
        RECT 106.010 112.190 106.960 113.400 ;
      LAYER li1 ;
        RECT 103.940 111.800 105.830 111.970 ;
        RECT 103.940 111.670 104.110 111.800 ;
        RECT 106.610 111.670 106.940 112.010 ;
        RECT 102.850 111.440 104.110 111.670 ;
      LAYER li1 ;
        RECT 104.290 111.490 106.320 111.620 ;
        RECT 107.140 111.490 107.390 113.650 ;
        RECT 107.770 113.620 109.220 113.650 ;
        RECT 107.770 113.450 108.020 113.620 ;
        RECT 108.190 113.450 108.380 113.620 ;
        RECT 108.550 113.450 108.820 113.620 ;
        RECT 108.990 113.450 109.220 113.620 ;
        RECT 107.770 112.580 109.220 113.450 ;
        RECT 110.070 113.570 110.660 113.600 ;
        RECT 110.070 113.400 110.100 113.570 ;
        RECT 110.270 113.400 110.460 113.570 ;
        RECT 110.630 113.400 110.660 113.570 ;
        RECT 104.290 111.450 107.390 111.490 ;
      LAYER li1 ;
        RECT 103.940 111.270 104.110 111.440 ;
      LAYER li1 ;
        RECT 106.150 111.320 107.390 111.450 ;
        RECT 101.280 110.740 102.580 111.140 ;
        RECT 100.970 110.260 102.580 110.740 ;
        RECT 102.810 110.260 103.760 111.220 ;
      LAYER li1 ;
        RECT 103.940 111.100 105.750 111.270 ;
        RECT 103.940 110.390 104.190 111.100 ;
      LAYER li1 ;
        RECT 104.370 110.260 105.320 110.920 ;
      LAYER li1 ;
        RECT 105.500 110.390 105.750 111.100 ;
      LAYER li1 ;
        RECT 105.930 110.260 106.880 111.140 ;
        RECT 107.060 110.390 107.390 111.320 ;
        RECT 108.000 111.140 108.330 111.920 ;
        RECT 108.540 111.590 108.870 112.580 ;
        RECT 109.550 112.420 109.880 113.350 ;
        RECT 110.070 112.620 110.660 113.400 ;
        RECT 110.840 113.530 112.280 113.700 ;
        RECT 110.840 112.420 111.010 113.530 ;
        RECT 109.550 112.250 111.010 112.420 ;
        RECT 108.000 110.740 109.300 111.140 ;
        RECT 107.690 110.260 109.300 110.740 ;
        RECT 109.550 110.390 109.820 112.250 ;
      LAYER li1 ;
        RECT 110.000 111.070 110.330 112.040 ;
      LAYER li1 ;
        RECT 110.680 111.750 111.010 112.250 ;
        RECT 111.190 112.040 111.440 113.350 ;
        RECT 111.680 112.730 111.930 113.350 ;
        RECT 112.110 113.080 112.280 113.530 ;
        RECT 112.460 113.570 112.790 113.600 ;
        RECT 112.460 113.400 112.490 113.570 ;
        RECT 112.660 113.400 112.790 113.570 ;
        RECT 112.460 113.260 112.790 113.400 ;
        RECT 112.970 113.530 114.710 113.700 ;
        RECT 112.970 113.080 113.140 113.530 ;
        RECT 112.110 112.910 113.140 113.080 ;
        RECT 113.320 112.730 113.490 113.350 ;
        RECT 114.020 113.090 114.350 113.350 ;
        RECT 111.680 112.560 113.490 112.730 ;
        RECT 113.670 112.560 113.890 112.890 ;
        RECT 113.320 112.380 113.490 112.560 ;
        RECT 111.190 111.810 111.720 112.040 ;
        RECT 111.190 110.890 111.460 111.810 ;
      LAYER li1 ;
        RECT 112.140 111.510 112.680 112.380 ;
      LAYER li1 ;
        RECT 113.320 112.210 113.540 112.380 ;
        RECT 110.000 110.260 110.950 110.890 ;
        RECT 111.130 110.390 111.460 110.890 ;
        RECT 111.640 110.260 112.230 111.140 ;
      LAYER li1 ;
        RECT 112.510 110.520 112.680 111.510 ;
        RECT 112.860 110.700 113.190 112.000 ;
      LAYER li1 ;
        RECT 113.370 111.220 113.540 112.210 ;
        RECT 113.720 112.040 113.890 112.560 ;
        RECT 114.070 112.390 114.240 113.090 ;
        RECT 114.540 112.940 114.710 113.530 ;
        RECT 114.890 113.570 115.840 113.600 ;
        RECT 114.890 113.400 114.920 113.570 ;
        RECT 115.090 113.400 115.280 113.570 ;
        RECT 115.450 113.400 115.640 113.570 ;
        RECT 115.810 113.400 115.840 113.570 ;
        RECT 114.890 113.120 115.840 113.400 ;
        RECT 116.020 113.530 117.050 113.700 ;
        RECT 116.020 112.940 116.190 113.530 ;
        RECT 114.540 112.890 116.190 112.940 ;
        RECT 114.420 112.770 116.190 112.890 ;
        RECT 114.420 112.570 114.750 112.770 ;
        RECT 116.370 112.590 116.700 113.350 ;
        RECT 116.880 113.170 117.050 113.530 ;
        RECT 117.230 113.570 118.180 113.650 ;
        RECT 117.230 113.400 117.260 113.570 ;
        RECT 117.430 113.400 117.620 113.570 ;
        RECT 117.790 113.400 117.980 113.570 ;
        RECT 118.150 113.400 118.180 113.570 ;
        RECT 117.230 113.350 118.180 113.400 ;
        RECT 116.880 113.000 118.690 113.170 ;
        RECT 114.930 112.420 116.700 112.590 ;
        RECT 114.930 112.390 115.100 112.420 ;
        RECT 114.070 112.220 115.100 112.390 ;
        RECT 118.010 112.240 118.340 112.820 ;
        RECT 113.720 111.810 114.750 112.040 ;
        RECT 114.420 111.320 114.750 111.810 ;
        RECT 114.930 111.540 115.100 112.220 ;
        RECT 115.280 112.070 118.340 112.240 ;
        RECT 115.280 111.720 115.610 112.070 ;
      LAYER li1 ;
        RECT 116.050 111.720 117.900 111.890 ;
      LAYER li1 ;
        RECT 114.930 111.370 117.550 111.540 ;
        RECT 113.370 110.720 113.640 111.220 ;
        RECT 114.930 111.140 115.100 111.370 ;
      LAYER li1 ;
        RECT 117.730 111.190 117.900 111.720 ;
      LAYER li1 ;
        RECT 114.090 110.970 115.100 111.140 ;
      LAYER li1 ;
        RECT 115.280 111.020 117.900 111.190 ;
      LAYER li1 ;
        RECT 114.090 110.720 114.420 110.970 ;
      LAYER li1 ;
        RECT 115.280 110.520 115.450 111.020 ;
        RECT 112.510 110.350 115.450 110.520 ;
      LAYER li1 ;
        RECT 116.600 110.260 117.550 110.840 ;
      LAYER li1 ;
        RECT 117.730 110.330 117.900 111.020 ;
      LAYER li1 ;
        RECT 118.080 111.220 118.340 112.070 ;
        RECT 118.520 111.650 118.690 113.000 ;
        RECT 118.870 112.740 119.120 113.650 ;
        RECT 119.930 113.570 120.880 113.600 ;
        RECT 121.710 113.570 122.610 113.600 ;
        RECT 119.930 113.400 119.960 113.570 ;
        RECT 120.130 113.400 120.320 113.570 ;
        RECT 120.490 113.400 120.680 113.570 ;
        RECT 120.850 113.400 120.880 113.570 ;
        RECT 121.880 113.400 122.070 113.570 ;
        RECT 122.240 113.400 122.430 113.570 ;
        RECT 122.600 113.400 122.610 113.570 ;
        RECT 118.870 112.570 119.750 112.740 ;
        RECT 119.930 112.570 120.880 113.400 ;
        RECT 121.280 112.600 121.530 113.070 ;
        RECT 121.710 112.780 122.610 113.400 ;
        RECT 123.220 113.570 124.160 113.630 ;
        RECT 123.220 113.400 123.240 113.570 ;
        RECT 123.410 113.400 123.600 113.570 ;
        RECT 123.770 113.400 123.960 113.570 ;
        RECT 124.130 113.400 124.160 113.570 ;
        RECT 119.070 111.830 119.400 112.330 ;
        RECT 119.580 112.250 119.750 112.570 ;
        RECT 121.280 112.430 122.290 112.600 ;
        RECT 119.580 112.080 121.940 112.250 ;
        RECT 118.520 111.480 119.690 111.650 ;
        RECT 118.080 110.510 118.410 111.220 ;
        RECT 118.870 110.680 119.200 111.220 ;
        RECT 119.410 110.980 119.690 111.480 ;
        RECT 119.870 110.680 120.040 112.080 ;
        RECT 122.120 111.900 122.290 112.430 ;
        RECT 120.250 111.730 122.290 111.900 ;
        RECT 120.250 111.340 120.580 111.730 ;
      LAYER li1 ;
        RECT 120.900 111.270 121.230 111.550 ;
        RECT 120.900 111.160 121.280 111.270 ;
      LAYER li1 ;
        RECT 118.870 110.510 120.040 110.680 ;
      LAYER li1 ;
        RECT 120.220 111.100 121.280 111.160 ;
        RECT 120.220 110.990 121.230 111.100 ;
        RECT 120.220 110.330 120.390 110.990 ;
      LAYER li1 ;
        RECT 122.060 110.890 122.290 111.730 ;
        RECT 122.790 111.900 123.040 112.900 ;
        RECT 123.220 112.090 124.160 113.400 ;
        RECT 122.790 111.570 124.160 111.900 ;
        RECT 122.790 111.390 123.000 111.570 ;
        RECT 122.670 110.890 123.000 111.390 ;
      LAYER li1 ;
        RECT 117.730 110.160 120.390 110.330 ;
      LAYER li1 ;
        RECT 120.570 110.260 121.520 110.810 ;
        RECT 122.060 110.390 122.390 110.890 ;
        RECT 123.180 110.260 124.130 111.390 ;
      LAYER li1 ;
        RECT 124.340 110.560 124.680 113.630 ;
      LAYER li1 ;
        RECT 125.300 113.620 128.040 113.640 ;
        RECT 125.300 113.450 125.510 113.620 ;
        RECT 125.680 113.450 125.950 113.620 ;
        RECT 126.120 113.450 126.360 113.620 ;
        RECT 126.530 113.450 126.790 113.620 ;
        RECT 126.960 113.450 127.230 113.620 ;
        RECT 127.400 113.450 127.640 113.620 ;
        RECT 127.810 113.450 128.040 113.620 ;
        RECT 125.300 112.570 128.040 113.450 ;
        RECT 129.140 113.620 131.880 113.640 ;
        RECT 129.140 113.450 129.350 113.620 ;
        RECT 129.520 113.450 129.790 113.620 ;
        RECT 129.960 113.450 130.200 113.620 ;
        RECT 130.370 113.450 130.630 113.620 ;
        RECT 130.800 113.450 131.070 113.620 ;
        RECT 131.240 113.450 131.480 113.620 ;
        RECT 131.650 113.450 131.880 113.620 ;
        RECT 129.140 112.570 131.880 113.450 ;
        RECT 132.980 113.620 135.720 113.640 ;
        RECT 132.980 113.450 133.190 113.620 ;
        RECT 133.360 113.450 133.630 113.620 ;
        RECT 133.800 113.450 134.040 113.620 ;
        RECT 134.210 113.450 134.470 113.620 ;
        RECT 134.640 113.450 134.910 113.620 ;
        RECT 135.080 113.450 135.320 113.620 ;
        RECT 135.490 113.450 135.720 113.620 ;
        RECT 132.980 112.570 135.720 113.450 ;
        RECT 136.820 113.620 139.560 113.640 ;
        RECT 136.820 113.450 137.030 113.620 ;
        RECT 137.200 113.450 137.470 113.620 ;
        RECT 137.640 113.450 137.880 113.620 ;
        RECT 138.050 113.450 138.310 113.620 ;
        RECT 138.480 113.450 138.750 113.620 ;
        RECT 138.920 113.450 139.160 113.620 ;
        RECT 139.330 113.450 139.560 113.620 ;
        RECT 136.820 112.570 139.560 113.450 ;
        RECT 140.410 113.620 141.860 113.650 ;
        RECT 140.410 113.450 140.660 113.620 ;
        RECT 140.830 113.450 141.020 113.620 ;
        RECT 141.190 113.450 141.460 113.620 ;
        RECT 141.630 113.450 141.860 113.620 ;
        RECT 140.410 112.580 141.860 113.450 ;
        RECT 125.540 111.250 125.870 111.920 ;
        RECT 126.270 111.590 126.600 112.570 ;
        RECT 126.820 111.250 127.150 111.920 ;
        RECT 127.550 111.590 127.880 112.570 ;
        RECT 129.380 111.250 129.710 111.920 ;
        RECT 130.110 111.590 130.440 112.570 ;
        RECT 130.660 111.250 130.990 111.920 ;
        RECT 131.390 111.590 131.720 112.570 ;
        RECT 133.220 111.250 133.550 111.920 ;
        RECT 133.950 111.590 134.280 112.570 ;
        RECT 134.500 111.250 134.830 111.920 ;
        RECT 135.230 111.590 135.560 112.570 ;
        RECT 137.060 111.250 137.390 111.920 ;
        RECT 137.790 111.590 138.120 112.570 ;
        RECT 138.340 111.250 138.670 111.920 ;
        RECT 139.070 111.590 139.400 112.570 ;
        RECT 125.380 110.250 128.110 111.250 ;
        RECT 129.220 110.250 131.950 111.250 ;
        RECT 133.060 110.250 135.790 111.250 ;
        RECT 136.900 110.250 139.630 111.250 ;
        RECT 140.640 111.140 140.970 111.920 ;
        RECT 141.180 111.590 141.510 112.580 ;
        RECT 140.640 110.740 141.940 111.140 ;
        RECT 140.330 110.260 141.940 110.740 ;
        RECT 5.760 109.800 5.920 109.980 ;
        RECT 6.090 109.800 6.400 109.980 ;
        RECT 6.570 109.800 6.880 109.980 ;
        RECT 7.050 109.800 7.360 109.980 ;
        RECT 7.530 109.800 7.840 109.980 ;
        RECT 8.010 109.800 8.320 109.980 ;
        RECT 8.490 109.800 8.800 109.980 ;
        RECT 8.970 109.800 9.280 109.980 ;
        RECT 9.450 109.800 9.760 109.980 ;
        RECT 9.930 109.800 10.240 109.980 ;
        RECT 10.410 109.800 10.720 109.980 ;
        RECT 10.890 109.800 11.200 109.980 ;
        RECT 11.370 109.800 11.680 109.980 ;
        RECT 11.850 109.800 12.160 109.980 ;
        RECT 12.330 109.800 12.640 109.980 ;
        RECT 12.810 109.800 13.120 109.980 ;
        RECT 13.290 109.800 13.600 109.980 ;
        RECT 13.770 109.800 14.080 109.980 ;
        RECT 14.250 109.800 14.560 109.980 ;
        RECT 14.730 109.800 15.040 109.980 ;
        RECT 15.210 109.800 15.520 109.980 ;
        RECT 15.690 109.800 16.000 109.980 ;
        RECT 16.170 109.800 16.480 109.980 ;
        RECT 16.650 109.800 16.960 109.980 ;
        RECT 17.130 109.800 17.440 109.980 ;
        RECT 17.610 109.800 17.920 109.980 ;
        RECT 18.090 109.800 18.400 109.980 ;
        RECT 18.570 109.800 18.880 109.980 ;
        RECT 19.050 109.800 19.360 109.980 ;
        RECT 19.530 109.800 19.840 109.980 ;
        RECT 20.010 109.800 20.320 109.980 ;
        RECT 20.490 109.800 20.800 109.980 ;
        RECT 20.970 109.800 21.280 109.980 ;
        RECT 21.450 109.800 21.760 109.980 ;
        RECT 21.930 109.800 22.240 109.980 ;
        RECT 22.410 109.800 22.720 109.980 ;
        RECT 22.890 109.800 23.200 109.980 ;
        RECT 23.370 109.800 23.680 109.980 ;
        RECT 23.850 109.800 24.000 109.980 ;
        RECT 24.480 109.800 24.640 109.980 ;
        RECT 24.810 109.800 25.120 109.980 ;
        RECT 25.290 109.800 25.600 109.980 ;
        RECT 25.770 109.800 26.080 109.980 ;
        RECT 26.250 109.800 26.560 109.980 ;
        RECT 26.730 109.800 27.040 109.980 ;
        RECT 27.210 109.800 27.520 109.980 ;
        RECT 27.690 109.800 28.000 109.980 ;
        RECT 28.170 109.800 28.480 109.980 ;
        RECT 28.650 109.800 28.960 109.980 ;
        RECT 29.130 109.800 29.440 109.980 ;
        RECT 29.610 109.800 29.920 109.980 ;
        RECT 30.090 109.800 30.400 109.980 ;
        RECT 30.570 109.800 30.880 109.980 ;
        RECT 31.050 109.800 31.360 109.980 ;
        RECT 31.530 109.800 31.840 109.980 ;
        RECT 32.010 109.800 32.320 109.980 ;
        RECT 32.490 109.800 32.800 109.980 ;
        RECT 32.970 109.800 33.280 109.980 ;
        RECT 33.450 109.800 33.760 109.980 ;
        RECT 33.930 109.800 34.240 109.980 ;
        RECT 34.410 109.800 34.720 109.980 ;
        RECT 34.890 109.800 35.200 109.980 ;
        RECT 35.370 109.800 35.680 109.980 ;
        RECT 35.850 109.800 36.160 109.980 ;
        RECT 36.330 109.800 36.640 109.980 ;
        RECT 36.810 109.800 36.960 109.980 ;
        RECT 37.440 109.800 37.600 109.980 ;
        RECT 37.770 109.800 38.080 109.980 ;
        RECT 38.250 109.800 38.560 109.980 ;
        RECT 38.730 109.800 39.040 109.980 ;
        RECT 39.210 109.800 39.520 109.980 ;
        RECT 39.690 109.800 40.000 109.980 ;
        RECT 40.170 109.800 40.480 109.980 ;
        RECT 40.650 109.800 40.960 109.980 ;
        RECT 41.130 109.800 41.440 109.980 ;
        RECT 41.610 109.800 41.920 109.980 ;
        RECT 42.090 109.800 42.400 109.980 ;
        RECT 42.570 109.800 42.880 109.980 ;
        RECT 43.050 109.800 43.360 109.980 ;
        RECT 43.530 109.800 43.840 109.980 ;
        RECT 44.010 109.800 44.320 109.980 ;
        RECT 44.490 109.800 44.800 109.980 ;
        RECT 44.970 109.800 45.280 109.980 ;
        RECT 45.450 109.800 45.760 109.980 ;
        RECT 45.930 109.800 46.240 109.980 ;
        RECT 46.410 109.800 46.720 109.980 ;
        RECT 46.890 109.800 47.200 109.980 ;
        RECT 47.370 109.800 47.680 109.980 ;
        RECT 47.850 109.800 48.160 109.980 ;
        RECT 48.330 109.800 48.640 109.980 ;
        RECT 48.810 109.800 49.120 109.980 ;
        RECT 49.290 109.800 49.600 109.980 ;
        RECT 49.770 109.800 50.080 109.980 ;
        RECT 50.250 109.800 50.560 109.980 ;
        RECT 50.730 109.800 51.040 109.980 ;
        RECT 51.210 109.800 51.520 109.980 ;
        RECT 51.690 109.800 52.000 109.980 ;
        RECT 52.170 109.800 52.480 109.980 ;
        RECT 52.650 109.800 52.960 109.980 ;
        RECT 53.130 109.800 53.440 109.980 ;
        RECT 53.610 109.800 53.920 109.980 ;
        RECT 54.090 109.800 54.400 109.980 ;
        RECT 54.570 109.800 54.880 109.980 ;
        RECT 55.050 109.800 55.360 109.980 ;
        RECT 55.530 109.800 55.840 109.980 ;
        RECT 56.010 109.800 56.320 109.980 ;
        RECT 56.490 109.800 56.800 109.980 ;
        RECT 56.970 109.800 57.280 109.980 ;
        RECT 57.450 109.800 57.760 109.980 ;
        RECT 57.930 109.800 58.240 109.980 ;
        RECT 58.410 109.800 58.720 109.980 ;
        RECT 58.890 109.800 59.200 109.980 ;
        RECT 59.370 109.800 59.680 109.980 ;
        RECT 59.850 109.800 60.160 109.980 ;
        RECT 60.330 109.800 60.640 109.980 ;
        RECT 60.810 109.800 61.120 109.980 ;
        RECT 61.290 109.800 61.600 109.980 ;
        RECT 61.770 109.800 62.080 109.980 ;
        RECT 62.250 109.800 62.560 109.980 ;
        RECT 62.730 109.800 63.040 109.980 ;
        RECT 63.210 109.800 63.520 109.980 ;
        RECT 63.690 109.800 64.000 109.980 ;
        RECT 64.170 109.800 64.480 109.980 ;
        RECT 64.650 109.800 64.960 109.980 ;
        RECT 65.130 109.800 65.440 109.980 ;
        RECT 65.610 109.800 65.920 109.980 ;
        RECT 66.090 109.800 66.400 109.980 ;
        RECT 66.570 109.800 66.880 109.980 ;
        RECT 67.050 109.800 67.360 109.980 ;
        RECT 67.530 109.800 67.840 109.980 ;
        RECT 68.010 109.800 68.320 109.980 ;
        RECT 68.490 109.800 68.800 109.980 ;
        RECT 68.970 109.800 69.280 109.980 ;
        RECT 69.450 109.800 69.760 109.980 ;
        RECT 69.930 109.800 70.240 109.980 ;
        RECT 70.410 109.800 70.720 109.980 ;
        RECT 70.890 109.800 71.200 109.980 ;
        RECT 71.370 109.800 71.520 109.980 ;
        RECT 72.000 109.800 72.160 109.980 ;
        RECT 72.330 109.800 72.640 109.980 ;
        RECT 72.810 109.800 73.120 109.980 ;
        RECT 73.290 109.800 73.600 109.980 ;
        RECT 73.770 109.800 74.080 109.980 ;
        RECT 74.250 109.800 74.560 109.980 ;
        RECT 74.730 109.800 75.040 109.980 ;
        RECT 75.210 109.800 75.520 109.980 ;
        RECT 75.690 109.800 76.000 109.980 ;
        RECT 76.170 109.800 76.480 109.980 ;
        RECT 76.650 109.800 76.960 109.980 ;
        RECT 77.130 109.800 77.440 109.980 ;
        RECT 77.610 109.800 77.920 109.980 ;
        RECT 78.090 109.800 78.400 109.980 ;
        RECT 78.570 109.800 78.880 109.980 ;
        RECT 79.050 109.800 79.360 109.980 ;
        RECT 79.530 109.800 79.840 109.980 ;
        RECT 80.010 109.800 80.320 109.980 ;
        RECT 80.490 109.800 80.800 109.980 ;
        RECT 80.970 109.800 81.280 109.980 ;
        RECT 81.450 109.800 81.760 109.980 ;
        RECT 81.930 109.800 82.240 109.980 ;
        RECT 82.410 109.800 82.720 109.980 ;
        RECT 82.890 109.800 83.200 109.980 ;
        RECT 83.370 109.800 83.680 109.980 ;
        RECT 83.850 109.800 84.160 109.980 ;
        RECT 84.330 109.800 84.640 109.980 ;
        RECT 84.810 109.800 85.120 109.980 ;
        RECT 85.290 109.800 85.600 109.980 ;
        RECT 85.770 109.800 86.080 109.980 ;
        RECT 86.250 109.800 86.560 109.980 ;
        RECT 86.730 109.800 87.040 109.980 ;
        RECT 87.210 109.800 87.520 109.980 ;
        RECT 87.690 109.800 88.000 109.980 ;
        RECT 88.170 109.800 88.480 109.980 ;
        RECT 88.650 109.800 88.960 109.980 ;
        RECT 89.130 109.800 89.440 109.980 ;
        RECT 89.610 109.800 89.920 109.980 ;
        RECT 90.090 109.800 90.400 109.980 ;
        RECT 90.570 109.800 90.880 109.980 ;
        RECT 91.050 109.800 91.360 109.980 ;
        RECT 91.530 109.800 91.840 109.980 ;
        RECT 92.010 109.800 92.320 109.980 ;
        RECT 92.490 109.800 92.800 109.980 ;
        RECT 92.970 109.800 93.280 109.980 ;
        RECT 93.450 109.800 93.760 109.980 ;
        RECT 93.930 109.800 94.240 109.980 ;
        RECT 94.410 109.800 94.720 109.980 ;
        RECT 94.890 109.800 95.200 109.980 ;
        RECT 95.370 109.800 95.680 109.980 ;
        RECT 95.850 109.800 96.160 109.980 ;
        RECT 96.330 109.800 96.640 109.980 ;
        RECT 96.810 109.800 97.120 109.980 ;
        RECT 97.290 109.800 97.600 109.980 ;
        RECT 97.770 109.800 98.080 109.980 ;
        RECT 98.250 109.800 98.560 109.980 ;
        RECT 98.730 109.800 99.040 109.980 ;
        RECT 99.210 109.800 99.520 109.980 ;
        RECT 99.690 109.800 100.000 109.980 ;
        RECT 100.170 109.800 100.480 109.980 ;
        RECT 100.650 109.800 100.960 109.980 ;
        RECT 101.130 109.800 101.440 109.980 ;
        RECT 101.610 109.800 101.920 109.980 ;
        RECT 102.090 109.800 102.400 109.980 ;
        RECT 102.570 109.800 102.880 109.980 ;
        RECT 103.050 109.800 103.360 109.980 ;
        RECT 103.530 109.800 103.840 109.980 ;
        RECT 104.010 109.800 104.320 109.980 ;
        RECT 104.490 109.800 104.800 109.980 ;
        RECT 104.970 109.800 105.280 109.980 ;
        RECT 105.450 109.800 105.760 109.980 ;
        RECT 105.930 109.800 106.240 109.980 ;
        RECT 106.410 109.800 106.720 109.980 ;
        RECT 106.890 109.800 107.200 109.980 ;
        RECT 107.370 109.800 107.680 109.980 ;
        RECT 107.850 109.800 108.160 109.980 ;
        RECT 108.330 109.800 108.640 109.980 ;
        RECT 108.810 109.800 109.120 109.980 ;
        RECT 109.290 109.800 109.600 109.980 ;
        RECT 109.770 109.800 110.080 109.980 ;
        RECT 110.250 109.800 110.560 109.980 ;
        RECT 110.730 109.800 111.040 109.980 ;
        RECT 111.210 109.800 111.520 109.980 ;
        RECT 111.690 109.800 112.000 109.980 ;
        RECT 112.170 109.800 112.480 109.980 ;
        RECT 112.650 109.800 112.960 109.980 ;
        RECT 113.130 109.800 113.440 109.980 ;
        RECT 113.610 109.800 113.920 109.980 ;
        RECT 114.090 109.800 114.400 109.980 ;
        RECT 114.570 109.800 114.880 109.980 ;
        RECT 115.050 109.800 115.360 109.980 ;
        RECT 115.530 109.800 115.840 109.980 ;
        RECT 116.010 109.800 116.320 109.980 ;
        RECT 116.490 109.800 116.800 109.980 ;
        RECT 116.970 109.800 117.280 109.980 ;
        RECT 117.450 109.800 117.760 109.980 ;
        RECT 117.930 109.800 118.240 109.980 ;
        RECT 118.410 109.800 118.720 109.980 ;
        RECT 118.890 109.800 119.200 109.980 ;
        RECT 119.370 109.800 119.680 109.980 ;
        RECT 119.850 109.800 120.160 109.980 ;
        RECT 120.330 109.800 120.640 109.980 ;
        RECT 120.810 109.800 121.120 109.980 ;
        RECT 121.290 109.800 121.600 109.980 ;
        RECT 121.770 109.800 122.080 109.980 ;
        RECT 122.250 109.800 122.560 109.980 ;
        RECT 122.730 109.800 123.040 109.980 ;
        RECT 123.210 109.800 123.520 109.980 ;
        RECT 123.690 109.800 124.000 109.980 ;
        RECT 124.170 109.800 124.480 109.980 ;
        RECT 124.650 109.800 124.960 109.980 ;
        RECT 125.130 109.800 125.440 109.980 ;
        RECT 125.610 109.800 125.920 109.980 ;
        RECT 126.090 109.800 126.400 109.980 ;
        RECT 126.570 109.800 126.880 109.980 ;
        RECT 127.050 109.800 127.360 109.980 ;
        RECT 127.530 109.800 127.840 109.980 ;
        RECT 128.010 109.800 128.320 109.980 ;
        RECT 128.490 109.800 128.800 109.980 ;
        RECT 128.970 109.800 129.280 109.980 ;
        RECT 129.450 109.800 129.760 109.980 ;
        RECT 129.930 109.800 130.240 109.980 ;
        RECT 130.410 109.800 130.720 109.980 ;
        RECT 130.890 109.800 131.200 109.980 ;
        RECT 131.370 109.800 131.680 109.980 ;
        RECT 131.850 109.800 132.160 109.980 ;
        RECT 132.330 109.800 132.640 109.980 ;
        RECT 132.810 109.800 133.120 109.980 ;
        RECT 133.290 109.800 133.600 109.980 ;
        RECT 133.770 109.800 134.080 109.980 ;
        RECT 134.250 109.800 134.560 109.980 ;
        RECT 134.730 109.800 135.040 109.980 ;
        RECT 135.210 109.800 135.520 109.980 ;
        RECT 135.690 109.800 136.000 109.980 ;
        RECT 136.170 109.800 136.480 109.980 ;
        RECT 136.650 109.800 136.960 109.980 ;
        RECT 137.130 109.800 137.440 109.980 ;
        RECT 137.610 109.800 137.920 109.980 ;
        RECT 138.090 109.800 138.400 109.980 ;
        RECT 138.570 109.800 138.880 109.980 ;
        RECT 139.050 109.800 139.360 109.980 ;
        RECT 139.530 109.800 139.840 109.980 ;
        RECT 140.010 109.800 140.320 109.980 ;
        RECT 140.490 109.800 140.800 109.980 ;
        RECT 140.970 109.800 141.280 109.980 ;
        RECT 141.450 109.800 141.760 109.980 ;
        RECT 141.930 109.800 142.080 109.980 ;
        RECT 6.340 109.500 9.070 109.530 ;
        RECT 6.340 109.330 6.510 109.500 ;
        RECT 6.680 109.330 6.950 109.500 ;
        RECT 7.120 109.330 7.360 109.500 ;
        RECT 7.530 109.330 7.790 109.500 ;
        RECT 7.960 109.330 8.230 109.500 ;
        RECT 8.400 109.330 8.640 109.500 ;
        RECT 8.810 109.330 9.070 109.500 ;
        RECT 6.340 108.530 9.070 109.330 ;
        RECT 10.180 109.500 12.910 109.530 ;
        RECT 10.180 109.330 10.350 109.500 ;
        RECT 10.520 109.330 10.790 109.500 ;
        RECT 10.960 109.330 11.200 109.500 ;
        RECT 11.370 109.330 11.630 109.500 ;
        RECT 11.800 109.330 12.070 109.500 ;
        RECT 12.240 109.330 12.480 109.500 ;
        RECT 12.650 109.330 12.910 109.500 ;
        RECT 10.180 108.530 12.910 109.330 ;
        RECT 14.020 109.500 16.750 109.530 ;
        RECT 14.020 109.330 14.190 109.500 ;
        RECT 14.360 109.330 14.630 109.500 ;
        RECT 14.800 109.330 15.040 109.500 ;
        RECT 15.210 109.330 15.470 109.500 ;
        RECT 15.640 109.330 15.910 109.500 ;
        RECT 16.080 109.330 16.320 109.500 ;
        RECT 16.490 109.330 16.750 109.500 ;
        RECT 14.020 108.530 16.750 109.330 ;
        RECT 17.860 109.500 20.590 109.530 ;
        RECT 17.860 109.330 18.030 109.500 ;
        RECT 18.200 109.330 18.470 109.500 ;
        RECT 18.640 109.330 18.880 109.500 ;
        RECT 19.050 109.330 19.310 109.500 ;
        RECT 19.480 109.330 19.750 109.500 ;
        RECT 19.920 109.330 20.160 109.500 ;
        RECT 20.330 109.330 20.590 109.500 ;
        RECT 17.860 108.530 20.590 109.330 ;
        RECT 21.290 109.490 22.900 109.520 ;
        RECT 21.290 109.320 21.340 109.490 ;
        RECT 21.510 109.320 21.780 109.490 ;
        RECT 21.950 109.320 22.220 109.490 ;
        RECT 22.390 109.320 22.630 109.490 ;
        RECT 22.800 109.320 22.900 109.490 ;
        RECT 21.290 109.040 22.900 109.320 ;
        RECT 21.600 108.640 22.900 109.040 ;
        RECT 23.200 109.450 25.010 109.620 ;
        RECT 6.500 107.860 6.830 108.530 ;
        RECT 7.230 107.210 7.560 108.190 ;
        RECT 7.780 107.860 8.110 108.530 ;
        RECT 8.510 107.210 8.840 108.190 ;
        RECT 10.340 107.860 10.670 108.530 ;
        RECT 11.070 107.210 11.400 108.190 ;
        RECT 11.620 107.860 11.950 108.530 ;
        RECT 12.350 107.210 12.680 108.190 ;
        RECT 14.180 107.860 14.510 108.530 ;
        RECT 14.910 107.210 15.240 108.190 ;
        RECT 15.460 107.860 15.790 108.530 ;
        RECT 16.190 107.210 16.520 108.190 ;
        RECT 18.020 107.860 18.350 108.530 ;
        RECT 18.750 107.210 19.080 108.190 ;
        RECT 19.300 107.860 19.630 108.530 ;
        RECT 20.030 107.210 20.360 108.190 ;
        RECT 21.600 107.860 21.930 108.640 ;
        RECT 23.200 108.530 23.530 109.450 ;
      LAYER li1 ;
        RECT 23.780 108.530 24.310 109.270 ;
      LAYER li1 ;
        RECT 6.260 106.330 9.000 107.210 ;
        RECT 6.260 106.160 6.470 106.330 ;
        RECT 6.640 106.160 6.910 106.330 ;
        RECT 7.080 106.160 7.320 106.330 ;
        RECT 7.490 106.160 7.750 106.330 ;
        RECT 7.920 106.160 8.190 106.330 ;
        RECT 8.360 106.160 8.600 106.330 ;
        RECT 8.770 106.160 9.000 106.330 ;
        RECT 6.260 106.140 9.000 106.160 ;
        RECT 10.100 106.330 12.840 107.210 ;
        RECT 10.100 106.160 10.310 106.330 ;
        RECT 10.480 106.160 10.750 106.330 ;
        RECT 10.920 106.160 11.160 106.330 ;
        RECT 11.330 106.160 11.590 106.330 ;
        RECT 11.760 106.160 12.030 106.330 ;
        RECT 12.200 106.160 12.440 106.330 ;
        RECT 12.610 106.160 12.840 106.330 ;
        RECT 10.100 106.140 12.840 106.160 ;
        RECT 13.940 106.330 16.680 107.210 ;
        RECT 13.940 106.160 14.150 106.330 ;
        RECT 14.320 106.160 14.590 106.330 ;
        RECT 14.760 106.160 15.000 106.330 ;
        RECT 15.170 106.160 15.430 106.330 ;
        RECT 15.600 106.160 15.870 106.330 ;
        RECT 16.040 106.160 16.280 106.330 ;
        RECT 16.450 106.160 16.680 106.330 ;
        RECT 13.940 106.140 16.680 106.160 ;
        RECT 17.780 106.330 20.520 107.210 ;
        RECT 22.140 107.200 22.470 108.190 ;
      LAYER li1 ;
        RECT 23.170 108.020 23.590 108.350 ;
        RECT 23.780 107.960 23.950 108.530 ;
      LAYER li1 ;
        RECT 24.840 108.430 25.010 109.450 ;
        RECT 25.190 109.490 26.290 109.520 ;
        RECT 25.190 109.320 25.240 109.490 ;
        RECT 25.410 109.320 25.600 109.490 ;
        RECT 25.770 109.320 25.960 109.490 ;
        RECT 26.130 109.320 26.290 109.490 ;
        RECT 27.050 109.490 28.660 109.520 ;
        RECT 25.190 108.610 26.290 109.320 ;
        RECT 26.460 108.430 26.710 109.360 ;
        RECT 27.050 109.320 27.100 109.490 ;
        RECT 27.270 109.320 27.540 109.490 ;
        RECT 27.710 109.320 27.980 109.490 ;
        RECT 28.150 109.320 28.390 109.490 ;
        RECT 28.560 109.320 28.660 109.490 ;
        RECT 29.360 109.490 30.310 109.520 ;
        RECT 27.050 109.040 28.660 109.320 ;
      LAYER li1 ;
        RECT 24.130 108.140 24.640 108.350 ;
      LAYER li1 ;
        RECT 24.840 108.260 26.710 108.430 ;
        RECT 27.360 108.640 28.660 109.040 ;
      LAYER li1 ;
        RECT 23.780 107.790 24.840 107.960 ;
        RECT 24.570 107.710 24.840 107.790 ;
        RECT 25.290 107.770 25.800 108.080 ;
        RECT 26.050 107.770 26.760 108.080 ;
      LAYER li1 ;
        RECT 27.360 107.860 27.690 108.640 ;
        RECT 17.780 106.160 17.990 106.330 ;
        RECT 18.160 106.160 18.430 106.330 ;
        RECT 18.600 106.160 18.840 106.330 ;
        RECT 19.010 106.160 19.270 106.330 ;
        RECT 19.440 106.160 19.710 106.330 ;
        RECT 19.880 106.160 20.120 106.330 ;
        RECT 20.290 106.160 20.520 106.330 ;
        RECT 17.780 106.140 20.520 106.160 ;
        RECT 21.370 106.330 22.820 107.200 ;
        RECT 21.370 106.160 21.620 106.330 ;
        RECT 21.790 106.160 21.980 106.330 ;
        RECT 22.150 106.160 22.420 106.330 ;
        RECT 22.590 106.160 22.820 106.330 ;
        RECT 21.370 106.130 22.820 106.160 ;
        RECT 23.130 106.380 24.390 107.610 ;
      LAYER li1 ;
        RECT 24.570 106.630 25.090 107.710 ;
      LAYER li1 ;
        RECT 23.130 106.210 23.140 106.380 ;
        RECT 23.310 106.210 23.500 106.380 ;
        RECT 23.670 106.210 23.860 106.380 ;
        RECT 24.030 106.210 24.220 106.380 ;
        RECT 23.130 106.130 24.390 106.210 ;
      LAYER li1 ;
        RECT 24.920 106.130 25.090 106.630 ;
      LAYER li1 ;
        RECT 25.350 106.380 26.660 107.590 ;
        RECT 27.900 107.200 28.230 108.190 ;
        RECT 28.910 107.530 29.180 109.390 ;
        RECT 29.360 109.320 29.390 109.490 ;
        RECT 29.560 109.320 29.750 109.490 ;
        RECT 29.920 109.320 30.110 109.490 ;
        RECT 30.280 109.320 30.310 109.490 ;
        RECT 31.000 109.490 31.590 109.520 ;
        RECT 29.360 108.890 30.310 109.320 ;
        RECT 30.490 108.890 30.820 109.390 ;
        RECT 30.040 107.530 30.370 108.030 ;
        RECT 28.910 107.360 30.370 107.530 ;
        RECT 25.350 106.210 25.380 106.380 ;
        RECT 25.550 106.210 25.740 106.380 ;
        RECT 25.910 106.210 26.100 106.380 ;
        RECT 26.270 106.210 26.460 106.380 ;
        RECT 26.630 106.210 26.660 106.380 ;
        RECT 25.350 106.130 26.660 106.210 ;
        RECT 27.130 106.330 28.580 107.200 ;
        RECT 28.910 106.430 29.240 107.360 ;
        RECT 27.130 106.160 27.380 106.330 ;
        RECT 27.550 106.160 27.740 106.330 ;
        RECT 27.910 106.160 28.180 106.330 ;
        RECT 28.350 106.160 28.580 106.330 ;
        RECT 29.430 106.380 30.020 107.160 ;
        RECT 29.430 106.210 29.460 106.380 ;
        RECT 29.630 106.210 29.820 106.380 ;
        RECT 29.990 106.210 30.020 106.380 ;
        RECT 29.430 106.180 30.020 106.210 ;
        RECT 30.200 106.250 30.370 107.360 ;
        RECT 30.550 107.970 30.820 108.890 ;
        RECT 31.000 109.320 31.030 109.490 ;
        RECT 31.200 109.320 31.390 109.490 ;
        RECT 31.560 109.320 31.590 109.490 ;
        RECT 35.960 109.490 36.910 109.520 ;
        RECT 31.000 108.640 31.590 109.320 ;
      LAYER li1 ;
        RECT 31.870 109.260 34.810 109.430 ;
        RECT 31.870 108.310 32.040 109.260 ;
        RECT 31.830 108.270 32.040 108.310 ;
      LAYER li1 ;
        RECT 30.550 107.740 31.080 107.970 ;
        RECT 30.550 106.430 30.800 107.740 ;
      LAYER li1 ;
        RECT 31.500 107.400 32.040 108.270 ;
        RECT 32.220 107.780 32.550 109.080 ;
      LAYER li1 ;
        RECT 32.730 108.560 33.000 109.060 ;
        RECT 33.450 108.810 33.780 109.060 ;
        RECT 33.450 108.640 34.460 108.810 ;
        RECT 32.730 107.570 32.900 108.560 ;
        RECT 33.780 107.970 34.110 108.460 ;
        RECT 32.680 107.400 32.900 107.570 ;
        RECT 33.080 107.740 34.110 107.970 ;
        RECT 34.290 108.410 34.460 108.640 ;
      LAYER li1 ;
        RECT 34.640 108.760 34.810 109.260 ;
      LAYER li1 ;
        RECT 35.960 109.320 35.990 109.490 ;
        RECT 36.160 109.320 36.350 109.490 ;
        RECT 36.520 109.320 36.710 109.490 ;
        RECT 36.880 109.320 36.910 109.490 ;
        RECT 35.960 108.940 36.910 109.320 ;
      LAYER li1 ;
        RECT 37.090 109.450 39.750 109.620 ;
        RECT 37.090 108.760 37.260 109.450 ;
        RECT 34.640 108.590 37.260 108.760 ;
      LAYER li1 ;
        RECT 34.290 108.240 36.910 108.410 ;
        RECT 32.680 107.220 32.850 107.400 ;
        RECT 33.080 107.220 33.250 107.740 ;
        RECT 34.290 107.560 34.460 108.240 ;
      LAYER li1 ;
        RECT 37.090 108.060 37.260 108.590 ;
      LAYER li1 ;
        RECT 31.040 107.050 32.850 107.220 ;
        RECT 31.040 106.430 31.290 107.050 ;
        RECT 31.470 106.700 32.500 106.870 ;
        RECT 31.470 106.250 31.640 106.700 ;
        RECT 27.130 106.130 28.580 106.160 ;
        RECT 30.200 106.080 31.640 106.250 ;
        RECT 31.820 106.380 32.150 106.520 ;
        RECT 31.820 106.210 31.850 106.380 ;
        RECT 32.020 106.210 32.150 106.380 ;
        RECT 31.820 106.180 32.150 106.210 ;
        RECT 32.330 106.250 32.500 106.700 ;
        RECT 32.680 106.430 32.850 107.050 ;
        RECT 33.030 106.890 33.250 107.220 ;
        RECT 33.430 107.390 34.460 107.560 ;
        RECT 34.640 107.710 34.970 108.060 ;
      LAYER li1 ;
        RECT 35.410 107.890 37.260 108.060 ;
      LAYER li1 ;
        RECT 37.440 108.560 37.770 109.270 ;
        RECT 38.230 109.100 39.400 109.270 ;
        RECT 38.230 108.560 38.560 109.100 ;
        RECT 37.440 107.710 37.700 108.560 ;
        RECT 38.770 108.300 39.050 108.800 ;
        RECT 34.640 107.540 37.700 107.710 ;
        RECT 33.430 106.690 33.600 107.390 ;
        RECT 34.290 107.360 34.460 107.390 ;
        RECT 33.780 107.010 34.110 107.210 ;
        RECT 34.290 107.190 36.060 107.360 ;
        RECT 33.780 106.890 35.550 107.010 ;
        RECT 33.900 106.840 35.550 106.890 ;
        RECT 33.380 106.430 33.710 106.690 ;
        RECT 33.900 106.250 34.070 106.840 ;
        RECT 32.330 106.080 34.070 106.250 ;
        RECT 34.250 106.380 35.200 106.660 ;
        RECT 34.250 106.210 34.280 106.380 ;
        RECT 34.450 106.210 34.640 106.380 ;
        RECT 34.810 106.210 35.000 106.380 ;
        RECT 35.170 106.210 35.200 106.380 ;
        RECT 34.250 106.180 35.200 106.210 ;
        RECT 35.380 106.250 35.550 106.840 ;
        RECT 35.730 106.430 36.060 107.190 ;
        RECT 37.370 106.960 37.700 107.540 ;
        RECT 37.880 108.130 39.050 108.300 ;
        RECT 37.880 106.780 38.050 108.130 ;
        RECT 38.430 107.450 38.760 107.950 ;
        RECT 39.230 107.700 39.400 109.100 ;
      LAYER li1 ;
        RECT 39.580 108.790 39.750 109.450 ;
      LAYER li1 ;
        RECT 39.930 109.490 40.880 109.520 ;
        RECT 39.930 109.320 39.960 109.490 ;
        RECT 40.130 109.320 40.320 109.490 ;
        RECT 40.490 109.320 40.680 109.490 ;
        RECT 40.850 109.320 40.880 109.490 ;
        RECT 42.540 109.490 43.490 109.520 ;
        RECT 39.930 108.970 40.880 109.320 ;
        RECT 41.420 108.890 41.750 109.390 ;
        RECT 42.540 109.320 42.570 109.490 ;
        RECT 42.740 109.320 42.930 109.490 ;
        RECT 43.100 109.320 43.290 109.490 ;
        RECT 43.460 109.320 43.490 109.490 ;
      LAYER li1 ;
        RECT 39.580 108.620 40.590 108.790 ;
      LAYER li1 ;
        RECT 39.610 108.050 39.940 108.440 ;
      LAYER li1 ;
        RECT 40.260 108.230 40.590 108.620 ;
      LAYER li1 ;
        RECT 41.420 108.050 41.650 108.890 ;
        RECT 42.030 108.390 42.360 108.890 ;
        RECT 42.540 108.390 43.490 109.320 ;
        RECT 44.330 109.490 45.940 109.520 ;
        RECT 44.330 109.320 44.380 109.490 ;
        RECT 44.550 109.320 44.820 109.490 ;
        RECT 44.990 109.320 45.260 109.490 ;
        RECT 45.430 109.320 45.670 109.490 ;
        RECT 45.840 109.320 45.940 109.490 ;
        RECT 44.330 109.040 45.940 109.320 ;
        RECT 44.640 108.640 45.940 109.040 ;
        RECT 46.170 109.490 46.760 109.520 ;
        RECT 46.170 109.320 46.200 109.490 ;
        RECT 46.370 109.320 46.560 109.490 ;
        RECT 46.730 109.320 46.760 109.490 ;
        RECT 47.690 109.490 49.300 109.520 ;
        RECT 39.610 107.880 41.650 108.050 ;
        RECT 38.940 107.530 41.300 107.700 ;
        RECT 38.940 107.210 39.110 107.530 ;
        RECT 41.480 107.350 41.650 107.880 ;
        RECT 36.240 106.610 38.050 106.780 ;
        RECT 38.230 107.040 39.110 107.210 ;
        RECT 36.240 106.250 36.410 106.610 ;
        RECT 35.380 106.080 36.410 106.250 ;
        RECT 36.590 106.380 37.540 106.430 ;
        RECT 36.590 106.210 36.620 106.380 ;
        RECT 36.790 106.210 36.980 106.380 ;
        RECT 37.150 106.210 37.340 106.380 ;
        RECT 37.510 106.210 37.540 106.380 ;
        RECT 36.590 106.130 37.540 106.210 ;
        RECT 38.230 106.130 38.480 107.040 ;
        RECT 39.290 106.380 40.240 107.210 ;
        RECT 40.640 107.180 41.650 107.350 ;
        RECT 42.150 108.210 42.360 108.390 ;
        RECT 42.150 107.880 43.520 108.210 ;
        RECT 40.640 106.710 40.890 107.180 ;
        RECT 41.070 106.380 41.970 107.000 ;
        RECT 42.150 106.880 42.400 107.880 ;
        RECT 44.640 107.860 44.970 108.640 ;
        RECT 46.170 108.560 46.760 109.320 ;
        RECT 39.290 106.210 39.320 106.380 ;
        RECT 39.490 106.210 39.680 106.380 ;
        RECT 39.850 106.210 40.040 106.380 ;
        RECT 40.210 106.210 40.240 106.380 ;
        RECT 41.240 106.210 41.430 106.380 ;
        RECT 41.600 106.210 41.790 106.380 ;
        RECT 41.960 106.210 41.970 106.380 ;
        RECT 39.290 106.180 40.240 106.210 ;
        RECT 41.070 106.180 41.970 106.210 ;
        RECT 42.580 106.380 43.520 107.690 ;
        RECT 45.180 107.200 45.510 108.190 ;
      LAYER li1 ;
        RECT 47.100 107.710 47.430 109.390 ;
      LAYER li1 ;
        RECT 47.690 109.320 47.740 109.490 ;
        RECT 47.910 109.320 48.180 109.490 ;
        RECT 48.350 109.320 48.620 109.490 ;
        RECT 48.790 109.320 49.030 109.490 ;
        RECT 49.200 109.320 49.300 109.490 ;
        RECT 50.000 109.490 50.950 109.520 ;
        RECT 47.690 109.040 49.300 109.320 ;
        RECT 48.000 108.640 49.300 109.040 ;
        RECT 48.000 107.860 48.330 108.640 ;
        RECT 42.580 106.210 42.600 106.380 ;
        RECT 42.770 106.210 42.960 106.380 ;
        RECT 43.130 106.210 43.320 106.380 ;
        RECT 43.490 106.210 43.520 106.380 ;
        RECT 42.580 106.150 43.520 106.210 ;
        RECT 44.410 106.330 45.860 107.200 ;
        RECT 44.410 106.160 44.660 106.330 ;
        RECT 44.830 106.160 45.020 106.330 ;
        RECT 45.190 106.160 45.460 106.330 ;
        RECT 45.630 106.160 45.860 106.330 ;
        RECT 44.410 106.130 45.860 106.160 ;
        RECT 46.170 106.380 46.760 107.710 ;
        RECT 46.170 106.210 46.200 106.380 ;
        RECT 46.370 106.210 46.560 106.380 ;
        RECT 46.730 106.210 46.760 106.380 ;
        RECT 46.170 106.130 46.760 106.210 ;
      LAYER li1 ;
        RECT 47.040 106.130 47.430 107.710 ;
      LAYER li1 ;
        RECT 48.540 107.200 48.870 108.190 ;
        RECT 49.550 107.530 49.820 109.390 ;
        RECT 50.000 109.320 50.030 109.490 ;
        RECT 50.200 109.320 50.390 109.490 ;
        RECT 50.560 109.320 50.750 109.490 ;
        RECT 50.920 109.320 50.950 109.490 ;
        RECT 51.640 109.490 52.230 109.520 ;
        RECT 50.000 108.890 50.950 109.320 ;
        RECT 51.130 108.890 51.460 109.390 ;
        RECT 50.680 107.530 51.010 108.030 ;
        RECT 49.550 107.360 51.010 107.530 ;
        RECT 47.770 106.330 49.220 107.200 ;
        RECT 49.550 106.430 49.880 107.360 ;
        RECT 47.770 106.160 48.020 106.330 ;
        RECT 48.190 106.160 48.380 106.330 ;
        RECT 48.550 106.160 48.820 106.330 ;
        RECT 48.990 106.160 49.220 106.330 ;
        RECT 50.070 106.380 50.660 107.160 ;
        RECT 50.070 106.210 50.100 106.380 ;
        RECT 50.270 106.210 50.460 106.380 ;
        RECT 50.630 106.210 50.660 106.380 ;
        RECT 50.070 106.180 50.660 106.210 ;
        RECT 50.840 106.250 51.010 107.360 ;
        RECT 51.190 107.970 51.460 108.890 ;
        RECT 51.640 109.320 51.670 109.490 ;
        RECT 51.840 109.320 52.030 109.490 ;
        RECT 52.200 109.320 52.230 109.490 ;
        RECT 56.600 109.490 57.550 109.520 ;
        RECT 51.640 108.640 52.230 109.320 ;
      LAYER li1 ;
        RECT 52.510 109.260 55.450 109.430 ;
        RECT 52.510 108.270 52.680 109.260 ;
      LAYER li1 ;
        RECT 51.190 107.740 51.720 107.970 ;
        RECT 51.190 106.430 51.440 107.740 ;
      LAYER li1 ;
        RECT 52.140 107.400 52.680 108.270 ;
        RECT 52.860 107.780 53.190 109.080 ;
      LAYER li1 ;
        RECT 53.370 108.560 53.640 109.060 ;
        RECT 54.090 108.810 54.420 109.060 ;
        RECT 54.090 108.640 55.100 108.810 ;
        RECT 53.370 107.570 53.540 108.560 ;
        RECT 54.420 107.970 54.750 108.460 ;
        RECT 53.320 107.400 53.540 107.570 ;
        RECT 53.720 107.740 54.750 107.970 ;
        RECT 54.930 108.410 55.100 108.640 ;
      LAYER li1 ;
        RECT 55.280 108.760 55.450 109.260 ;
      LAYER li1 ;
        RECT 56.600 109.320 56.630 109.490 ;
        RECT 56.800 109.320 56.990 109.490 ;
        RECT 57.160 109.320 57.350 109.490 ;
        RECT 57.520 109.320 57.550 109.490 ;
        RECT 56.600 108.940 57.550 109.320 ;
      LAYER li1 ;
        RECT 57.730 109.450 60.390 109.620 ;
        RECT 57.730 108.760 57.900 109.450 ;
        RECT 55.280 108.590 57.900 108.760 ;
      LAYER li1 ;
        RECT 54.930 108.240 57.550 108.410 ;
        RECT 53.320 107.220 53.490 107.400 ;
        RECT 53.720 107.220 53.890 107.740 ;
        RECT 54.930 107.560 55.100 108.240 ;
      LAYER li1 ;
        RECT 57.730 108.060 57.900 108.590 ;
      LAYER li1 ;
        RECT 51.680 107.050 53.490 107.220 ;
        RECT 51.680 106.430 51.930 107.050 ;
        RECT 52.110 106.700 53.140 106.870 ;
        RECT 52.110 106.250 52.280 106.700 ;
        RECT 47.770 106.130 49.220 106.160 ;
        RECT 50.840 106.080 52.280 106.250 ;
        RECT 52.460 106.380 52.790 106.520 ;
        RECT 52.460 106.210 52.490 106.380 ;
        RECT 52.660 106.210 52.790 106.380 ;
        RECT 52.460 106.180 52.790 106.210 ;
        RECT 52.970 106.250 53.140 106.700 ;
        RECT 53.320 106.430 53.490 107.050 ;
        RECT 53.670 106.890 53.890 107.220 ;
        RECT 54.070 107.390 55.100 107.560 ;
        RECT 55.280 107.710 55.610 108.060 ;
      LAYER li1 ;
        RECT 56.050 107.890 57.900 108.060 ;
      LAYER li1 ;
        RECT 58.080 108.560 58.410 109.270 ;
        RECT 58.870 109.100 60.040 109.270 ;
        RECT 58.870 108.560 59.200 109.100 ;
        RECT 58.080 107.710 58.340 108.560 ;
        RECT 59.410 108.300 59.690 108.800 ;
        RECT 55.280 107.540 58.340 107.710 ;
        RECT 54.070 106.690 54.240 107.390 ;
        RECT 54.930 107.360 55.100 107.390 ;
        RECT 54.420 107.010 54.750 107.210 ;
        RECT 54.930 107.190 56.700 107.360 ;
        RECT 54.420 106.890 56.190 107.010 ;
        RECT 54.540 106.840 56.190 106.890 ;
        RECT 54.020 106.430 54.350 106.690 ;
        RECT 54.540 106.250 54.710 106.840 ;
        RECT 52.970 106.080 54.710 106.250 ;
        RECT 54.890 106.380 55.840 106.660 ;
        RECT 54.890 106.210 54.920 106.380 ;
        RECT 55.090 106.210 55.280 106.380 ;
        RECT 55.450 106.210 55.640 106.380 ;
        RECT 55.810 106.210 55.840 106.380 ;
        RECT 54.890 106.180 55.840 106.210 ;
        RECT 56.020 106.250 56.190 106.840 ;
        RECT 56.370 106.430 56.700 107.190 ;
        RECT 58.010 106.960 58.340 107.540 ;
        RECT 58.520 108.130 59.690 108.300 ;
        RECT 58.520 106.780 58.690 108.130 ;
        RECT 59.070 107.450 59.400 107.950 ;
        RECT 59.870 107.700 60.040 109.100 ;
      LAYER li1 ;
        RECT 60.220 108.790 60.390 109.450 ;
      LAYER li1 ;
        RECT 60.570 109.490 61.520 109.520 ;
        RECT 60.570 109.320 60.600 109.490 ;
        RECT 60.770 109.320 60.960 109.490 ;
        RECT 61.130 109.320 61.320 109.490 ;
        RECT 61.490 109.320 61.520 109.490 ;
        RECT 63.180 109.490 64.130 109.520 ;
        RECT 60.570 108.970 61.520 109.320 ;
        RECT 62.060 108.890 62.390 109.390 ;
        RECT 63.180 109.320 63.210 109.490 ;
        RECT 63.380 109.320 63.570 109.490 ;
        RECT 63.740 109.320 63.930 109.490 ;
        RECT 64.100 109.320 64.130 109.490 ;
      LAYER li1 ;
        RECT 60.220 108.680 61.230 108.790 ;
        RECT 60.220 108.620 61.280 108.680 ;
        RECT 60.900 108.510 61.280 108.620 ;
      LAYER li1 ;
        RECT 60.250 108.050 60.580 108.440 ;
      LAYER li1 ;
        RECT 60.900 108.230 61.230 108.510 ;
      LAYER li1 ;
        RECT 62.060 108.050 62.290 108.890 ;
        RECT 62.670 108.390 63.000 108.890 ;
        RECT 63.180 108.390 64.130 109.320 ;
        RECT 64.970 109.490 66.580 109.520 ;
        RECT 64.970 109.320 65.020 109.490 ;
        RECT 65.190 109.320 65.460 109.490 ;
        RECT 65.630 109.320 65.900 109.490 ;
        RECT 66.070 109.320 66.310 109.490 ;
        RECT 66.480 109.320 66.580 109.490 ;
        RECT 64.970 109.040 66.580 109.320 ;
        RECT 65.280 108.640 66.580 109.040 ;
        RECT 66.810 109.490 67.760 109.520 ;
        RECT 66.810 109.320 66.840 109.490 ;
        RECT 67.010 109.320 67.200 109.490 ;
        RECT 67.370 109.320 67.560 109.490 ;
        RECT 67.730 109.320 67.760 109.490 ;
        RECT 68.370 109.490 69.320 109.520 ;
        RECT 60.250 107.880 62.290 108.050 ;
        RECT 59.580 107.530 61.940 107.700 ;
        RECT 59.580 107.210 59.750 107.530 ;
        RECT 62.120 107.350 62.290 107.880 ;
        RECT 56.880 106.610 58.690 106.780 ;
        RECT 58.870 107.040 59.750 107.210 ;
        RECT 56.880 106.250 57.050 106.610 ;
        RECT 56.020 106.080 57.050 106.250 ;
        RECT 57.230 106.380 58.180 106.430 ;
        RECT 57.230 106.210 57.260 106.380 ;
        RECT 57.430 106.210 57.620 106.380 ;
        RECT 57.790 106.210 57.980 106.380 ;
        RECT 58.150 106.210 58.180 106.380 ;
        RECT 57.230 106.130 58.180 106.210 ;
        RECT 58.870 106.130 59.120 107.040 ;
        RECT 59.930 106.380 60.880 107.210 ;
        RECT 61.280 107.180 62.290 107.350 ;
        RECT 62.790 108.210 63.000 108.390 ;
        RECT 62.790 107.880 64.160 108.210 ;
        RECT 61.280 106.710 61.530 107.180 ;
        RECT 61.710 106.380 62.610 107.000 ;
        RECT 62.790 106.880 63.040 107.880 ;
        RECT 65.280 107.860 65.610 108.640 ;
        RECT 66.810 108.560 67.760 109.320 ;
      LAYER li1 ;
        RECT 67.940 108.680 68.190 109.390 ;
      LAYER li1 ;
        RECT 68.370 109.320 68.400 109.490 ;
        RECT 68.570 109.320 68.760 109.490 ;
        RECT 68.930 109.320 69.120 109.490 ;
        RECT 69.290 109.320 69.320 109.490 ;
        RECT 69.930 109.490 70.880 109.520 ;
        RECT 68.370 108.860 69.320 109.320 ;
      LAYER li1 ;
        RECT 69.500 108.680 69.750 109.390 ;
        RECT 67.940 108.510 69.750 108.680 ;
      LAYER li1 ;
        RECT 69.930 109.320 69.960 109.490 ;
        RECT 70.130 109.320 70.320 109.490 ;
        RECT 70.490 109.320 70.680 109.490 ;
        RECT 70.850 109.320 70.880 109.490 ;
        RECT 71.690 109.490 73.300 109.520 ;
        RECT 69.930 108.640 70.880 109.320 ;
      LAYER li1 ;
        RECT 67.940 108.340 68.110 108.510 ;
      LAYER li1 ;
        RECT 71.060 108.460 71.390 109.390 ;
        RECT 71.690 109.320 71.740 109.490 ;
        RECT 71.910 109.320 72.180 109.490 ;
        RECT 72.350 109.320 72.620 109.490 ;
        RECT 72.790 109.320 73.030 109.490 ;
        RECT 73.200 109.320 73.300 109.490 ;
        RECT 71.690 109.040 73.300 109.320 ;
        RECT 59.930 106.210 59.960 106.380 ;
        RECT 60.130 106.210 60.320 106.380 ;
        RECT 60.490 106.210 60.680 106.380 ;
        RECT 60.850 106.210 60.880 106.380 ;
        RECT 61.880 106.210 62.070 106.380 ;
        RECT 62.240 106.210 62.430 106.380 ;
        RECT 62.600 106.210 62.610 106.380 ;
        RECT 59.930 106.180 60.880 106.210 ;
        RECT 61.710 106.180 62.610 106.210 ;
        RECT 63.220 106.380 64.160 107.690 ;
        RECT 65.820 107.200 66.150 108.190 ;
      LAYER li1 ;
        RECT 66.850 108.110 68.110 108.340 ;
      LAYER li1 ;
        RECT 70.150 108.330 71.390 108.460 ;
        RECT 68.290 108.290 71.390 108.330 ;
        RECT 68.290 108.160 70.320 108.290 ;
      LAYER li1 ;
        RECT 67.940 107.980 68.110 108.110 ;
        RECT 67.940 107.810 69.830 107.980 ;
      LAYER li1 ;
        RECT 63.220 106.210 63.240 106.380 ;
        RECT 63.410 106.210 63.600 106.380 ;
        RECT 63.770 106.210 63.960 106.380 ;
        RECT 64.130 106.210 64.160 106.380 ;
        RECT 63.220 106.150 64.160 106.210 ;
        RECT 65.050 106.330 66.500 107.200 ;
        RECT 65.050 106.160 65.300 106.330 ;
        RECT 65.470 106.160 65.660 106.330 ;
        RECT 65.830 106.160 66.100 106.330 ;
        RECT 66.270 106.160 66.500 106.330 ;
        RECT 65.050 106.130 66.500 106.160 ;
        RECT 66.810 106.380 67.760 107.710 ;
        RECT 66.810 106.210 66.840 106.380 ;
        RECT 67.010 106.210 67.200 106.380 ;
        RECT 67.370 106.210 67.560 106.380 ;
        RECT 67.730 106.210 67.760 106.380 ;
        RECT 66.810 106.130 67.760 106.210 ;
      LAYER li1 ;
        RECT 67.940 106.130 68.190 107.810 ;
      LAYER li1 ;
        RECT 68.370 106.380 69.320 107.630 ;
        RECT 68.370 106.210 68.400 106.380 ;
        RECT 68.570 106.210 68.760 106.380 ;
        RECT 68.930 106.210 69.120 106.380 ;
        RECT 69.290 106.210 69.320 106.380 ;
        RECT 68.370 106.130 69.320 106.210 ;
      LAYER li1 ;
        RECT 69.500 106.130 69.830 107.810 ;
        RECT 70.610 107.770 70.940 108.110 ;
      LAYER li1 ;
        RECT 70.010 106.380 70.960 107.590 ;
        RECT 70.010 106.210 70.040 106.380 ;
        RECT 70.210 106.210 70.400 106.380 ;
        RECT 70.570 106.210 70.760 106.380 ;
        RECT 70.930 106.210 70.960 106.380 ;
        RECT 70.010 106.130 70.960 106.210 ;
        RECT 71.140 106.130 71.390 108.290 ;
        RECT 72.000 108.640 73.300 109.040 ;
        RECT 74.010 109.490 74.940 109.520 ;
        RECT 74.010 109.320 74.030 109.490 ;
        RECT 74.200 109.320 74.390 109.490 ;
        RECT 74.560 109.320 74.750 109.490 ;
        RECT 74.920 109.320 74.940 109.490 ;
        RECT 75.640 109.490 76.230 109.520 ;
        RECT 72.000 107.860 72.330 108.640 ;
        RECT 74.010 108.560 74.940 109.320 ;
      LAYER li1 ;
        RECT 75.120 108.460 75.450 109.390 ;
      LAYER li1 ;
        RECT 75.640 109.320 75.670 109.490 ;
        RECT 75.840 109.320 76.030 109.490 ;
        RECT 76.200 109.320 76.230 109.490 ;
        RECT 75.640 108.640 76.230 109.320 ;
        RECT 76.490 109.490 78.100 109.520 ;
        RECT 76.490 109.320 76.540 109.490 ;
        RECT 76.710 109.320 76.980 109.490 ;
        RECT 77.150 109.320 77.420 109.490 ;
        RECT 77.590 109.320 77.830 109.490 ;
        RECT 78.000 109.320 78.100 109.490 ;
        RECT 76.490 109.040 78.100 109.320 ;
        RECT 76.800 108.640 78.100 109.040 ;
        RECT 78.400 109.450 80.210 109.620 ;
      LAYER li1 ;
        RECT 75.120 108.290 76.200 108.460 ;
      LAYER li1 ;
        RECT 72.540 107.200 72.870 108.190 ;
      LAYER li1 ;
        RECT 74.050 107.770 75.240 108.110 ;
        RECT 75.420 107.770 75.750 108.110 ;
      LAYER li1 ;
        RECT 71.770 106.330 73.220 107.200 ;
        RECT 71.770 106.160 72.020 106.330 ;
        RECT 72.190 106.160 72.380 106.330 ;
        RECT 72.550 106.160 72.820 106.330 ;
        RECT 72.990 106.160 73.220 106.330 ;
        RECT 71.770 106.130 73.220 106.160 ;
        RECT 74.010 106.380 75.680 107.590 ;
        RECT 74.010 106.210 74.040 106.380 ;
        RECT 74.210 106.210 74.400 106.380 ;
        RECT 74.570 106.210 74.760 106.380 ;
        RECT 74.930 106.210 75.120 106.380 ;
        RECT 75.290 106.210 75.480 106.380 ;
        RECT 75.650 106.210 75.680 106.380 ;
        RECT 74.010 106.130 75.680 106.210 ;
      LAYER li1 ;
        RECT 75.940 106.130 76.200 108.290 ;
      LAYER li1 ;
        RECT 76.800 107.860 77.130 108.640 ;
        RECT 78.400 108.530 78.730 109.450 ;
      LAYER li1 ;
        RECT 78.980 108.530 79.510 109.270 ;
      LAYER li1 ;
        RECT 77.340 107.200 77.670 108.190 ;
      LAYER li1 ;
        RECT 78.370 108.020 78.790 108.350 ;
        RECT 78.980 107.960 79.150 108.530 ;
      LAYER li1 ;
        RECT 80.040 108.430 80.210 109.450 ;
        RECT 80.390 109.490 81.490 109.520 ;
        RECT 80.390 109.320 80.440 109.490 ;
        RECT 80.610 109.320 80.800 109.490 ;
        RECT 80.970 109.320 81.160 109.490 ;
        RECT 81.330 109.320 81.490 109.490 ;
        RECT 82.250 109.490 83.860 109.520 ;
        RECT 84.560 109.490 85.450 109.520 ;
        RECT 80.390 108.610 81.490 109.320 ;
        RECT 81.660 108.430 81.910 109.360 ;
        RECT 82.250 109.320 82.300 109.490 ;
        RECT 82.470 109.320 82.740 109.490 ;
        RECT 82.910 109.320 83.180 109.490 ;
        RECT 83.350 109.320 83.590 109.490 ;
        RECT 83.760 109.320 83.860 109.490 ;
        RECT 82.250 109.040 83.860 109.320 ;
      LAYER li1 ;
        RECT 79.330 108.140 79.840 108.350 ;
      LAYER li1 ;
        RECT 80.040 108.260 81.910 108.430 ;
        RECT 82.560 108.640 83.860 109.040 ;
      LAYER li1 ;
        RECT 78.980 107.790 80.040 107.960 ;
        RECT 79.770 107.710 80.040 107.790 ;
        RECT 80.490 107.770 81.000 108.080 ;
        RECT 81.250 107.770 81.960 108.080 ;
      LAYER li1 ;
        RECT 82.560 107.860 82.890 108.640 ;
        RECT 76.570 106.330 78.020 107.200 ;
        RECT 76.570 106.160 76.820 106.330 ;
        RECT 76.990 106.160 77.180 106.330 ;
        RECT 77.350 106.160 77.620 106.330 ;
        RECT 77.790 106.160 78.020 106.330 ;
        RECT 76.570 106.130 78.020 106.160 ;
        RECT 78.330 106.380 79.590 107.610 ;
      LAYER li1 ;
        RECT 79.770 106.630 80.290 107.710 ;
      LAYER li1 ;
        RECT 78.330 106.210 78.340 106.380 ;
        RECT 78.510 106.210 78.700 106.380 ;
        RECT 78.870 106.210 79.060 106.380 ;
        RECT 79.230 106.210 79.420 106.380 ;
        RECT 78.330 106.130 79.590 106.210 ;
      LAYER li1 ;
        RECT 80.120 106.130 80.290 106.630 ;
      LAYER li1 ;
        RECT 80.550 106.380 81.860 107.590 ;
        RECT 83.100 107.200 83.430 108.190 ;
        RECT 80.550 106.210 80.580 106.380 ;
        RECT 80.750 106.210 80.940 106.380 ;
        RECT 81.110 106.210 81.300 106.380 ;
        RECT 81.470 106.210 81.660 106.380 ;
        RECT 81.830 106.210 81.860 106.380 ;
        RECT 80.550 106.130 81.860 106.210 ;
        RECT 82.330 106.330 83.780 107.200 ;
        RECT 82.330 106.160 82.580 106.330 ;
        RECT 82.750 106.160 82.940 106.330 ;
        RECT 83.110 106.160 83.380 106.330 ;
        RECT 83.550 106.160 83.780 106.330 ;
        RECT 82.330 106.130 83.780 106.160 ;
      LAYER li1 ;
        RECT 84.130 106.130 84.380 109.390 ;
      LAYER li1 ;
        RECT 84.730 109.320 84.920 109.490 ;
        RECT 85.090 109.320 85.280 109.490 ;
        RECT 85.750 109.450 87.680 109.620 ;
        RECT 84.560 108.640 85.450 109.320 ;
        RECT 85.750 109.020 86.080 109.450 ;
        RECT 86.530 109.010 86.860 109.270 ;
        RECT 86.260 108.840 86.860 109.010 ;
        RECT 87.350 108.860 87.680 109.450 ;
        RECT 87.890 109.490 89.190 109.520 ;
        RECT 87.890 109.320 87.920 109.490 ;
        RECT 88.090 109.320 88.280 109.490 ;
        RECT 88.450 109.320 88.640 109.490 ;
        RECT 88.810 109.320 89.000 109.490 ;
        RECT 89.170 109.320 89.190 109.490 ;
        RECT 87.890 108.840 89.190 109.320 ;
        RECT 89.450 109.490 91.060 109.520 ;
        RECT 89.450 109.320 89.500 109.490 ;
        RECT 89.670 109.320 89.940 109.490 ;
        RECT 90.110 109.320 90.380 109.490 ;
        RECT 90.550 109.320 90.790 109.490 ;
        RECT 90.960 109.320 91.060 109.490 ;
        RECT 89.450 109.040 91.060 109.320 ;
        RECT 85.630 108.670 86.430 108.840 ;
        RECT 85.630 108.460 85.800 108.670 ;
      LAYER li1 ;
        RECT 87.040 108.660 87.710 108.680 ;
        RECT 86.610 108.490 88.880 108.660 ;
      LAYER li1 ;
        RECT 84.590 108.290 85.800 108.460 ;
      LAYER li1 ;
        RECT 85.980 108.320 86.780 108.490 ;
      LAYER li1 ;
        RECT 84.590 107.590 84.920 108.290 ;
      LAYER li1 ;
        RECT 85.980 108.110 86.150 108.320 ;
        RECT 85.420 107.830 86.150 108.110 ;
        RECT 85.590 107.770 85.760 107.830 ;
        RECT 86.330 107.770 86.760 108.140 ;
        RECT 86.960 107.770 87.250 108.310 ;
        RECT 87.490 107.980 88.200 108.310 ;
        RECT 88.550 107.870 88.880 108.490 ;
      LAYER li1 ;
        RECT 89.760 108.640 91.060 109.040 ;
        RECT 92.250 109.490 93.200 109.520 ;
        RECT 92.250 109.320 92.280 109.490 ;
        RECT 92.450 109.320 92.640 109.490 ;
        RECT 92.810 109.320 93.000 109.490 ;
        RECT 93.170 109.320 93.200 109.490 ;
        RECT 93.810 109.490 94.760 109.520 ;
        RECT 89.760 107.860 90.090 108.640 ;
        RECT 92.250 108.560 93.200 109.320 ;
      LAYER li1 ;
        RECT 93.380 108.680 93.630 109.390 ;
      LAYER li1 ;
        RECT 93.810 109.320 93.840 109.490 ;
        RECT 94.010 109.320 94.200 109.490 ;
        RECT 94.370 109.320 94.560 109.490 ;
        RECT 94.730 109.320 94.760 109.490 ;
        RECT 95.370 109.490 96.320 109.520 ;
        RECT 93.810 108.860 94.760 109.320 ;
      LAYER li1 ;
        RECT 94.940 108.680 95.190 109.390 ;
        RECT 93.380 108.510 95.190 108.680 ;
      LAYER li1 ;
        RECT 95.370 109.320 95.400 109.490 ;
        RECT 95.570 109.320 95.760 109.490 ;
        RECT 95.930 109.320 96.120 109.490 ;
        RECT 96.290 109.320 96.320 109.490 ;
        RECT 97.130 109.490 98.740 109.520 ;
        RECT 95.370 108.640 96.320 109.320 ;
      LAYER li1 ;
        RECT 93.380 108.340 93.550 108.510 ;
      LAYER li1 ;
        RECT 96.500 108.460 96.830 109.390 ;
        RECT 97.130 109.320 97.180 109.490 ;
        RECT 97.350 109.320 97.620 109.490 ;
        RECT 97.790 109.320 98.060 109.490 ;
        RECT 98.230 109.320 98.470 109.490 ;
        RECT 98.640 109.320 98.740 109.490 ;
        RECT 97.130 109.040 98.740 109.320 ;
        RECT 87.430 107.590 87.680 107.710 ;
        RECT 84.590 107.420 87.680 107.590 ;
        RECT 84.560 106.380 87.250 107.240 ;
        RECT 84.730 106.210 84.920 106.380 ;
        RECT 85.090 106.210 85.280 106.380 ;
        RECT 85.450 106.210 85.640 106.380 ;
        RECT 85.810 106.210 86.000 106.380 ;
        RECT 86.170 106.210 86.360 106.380 ;
        RECT 86.530 106.210 86.720 106.380 ;
        RECT 86.890 106.210 87.080 106.380 ;
        RECT 84.560 106.130 87.250 106.210 ;
        RECT 87.430 106.130 87.680 107.420 ;
        RECT 87.860 106.380 89.170 107.690 ;
        RECT 90.300 107.200 90.630 108.190 ;
      LAYER li1 ;
        RECT 92.290 108.110 93.550 108.340 ;
      LAYER li1 ;
        RECT 95.590 108.330 96.830 108.460 ;
        RECT 93.730 108.290 96.830 108.330 ;
        RECT 93.730 108.160 95.760 108.290 ;
      LAYER li1 ;
        RECT 93.380 107.980 93.550 108.110 ;
        RECT 93.380 107.810 95.270 107.980 ;
      LAYER li1 ;
        RECT 87.860 106.210 87.890 106.380 ;
        RECT 88.060 106.210 88.250 106.380 ;
        RECT 88.420 106.210 88.610 106.380 ;
        RECT 88.780 106.210 88.970 106.380 ;
        RECT 89.140 106.210 89.170 106.380 ;
        RECT 87.860 106.150 89.170 106.210 ;
        RECT 89.530 106.330 90.980 107.200 ;
        RECT 89.530 106.160 89.780 106.330 ;
        RECT 89.950 106.160 90.140 106.330 ;
        RECT 90.310 106.160 90.580 106.330 ;
        RECT 90.750 106.160 90.980 106.330 ;
        RECT 89.530 106.130 90.980 106.160 ;
        RECT 92.250 106.380 93.200 107.710 ;
        RECT 92.250 106.210 92.280 106.380 ;
        RECT 92.450 106.210 92.640 106.380 ;
        RECT 92.810 106.210 93.000 106.380 ;
        RECT 93.170 106.210 93.200 106.380 ;
        RECT 92.250 106.130 93.200 106.210 ;
      LAYER li1 ;
        RECT 93.380 106.130 93.630 107.810 ;
      LAYER li1 ;
        RECT 93.810 106.380 94.760 107.630 ;
        RECT 93.810 106.210 93.840 106.380 ;
        RECT 94.010 106.210 94.200 106.380 ;
        RECT 94.370 106.210 94.560 106.380 ;
        RECT 94.730 106.210 94.760 106.380 ;
        RECT 93.810 106.130 94.760 106.210 ;
      LAYER li1 ;
        RECT 94.940 106.130 95.270 107.810 ;
        RECT 96.050 107.770 96.380 108.110 ;
      LAYER li1 ;
        RECT 95.450 106.380 96.400 107.590 ;
        RECT 95.450 106.210 95.480 106.380 ;
        RECT 95.650 106.210 95.840 106.380 ;
        RECT 96.010 106.210 96.200 106.380 ;
        RECT 96.370 106.210 96.400 106.380 ;
        RECT 95.450 106.130 96.400 106.210 ;
        RECT 96.580 106.130 96.830 108.290 ;
        RECT 97.440 108.640 98.740 109.040 ;
        RECT 98.970 109.490 99.920 109.520 ;
        RECT 98.970 109.320 99.000 109.490 ;
        RECT 99.170 109.320 99.360 109.490 ;
        RECT 99.530 109.320 99.720 109.490 ;
        RECT 99.890 109.320 99.920 109.490 ;
        RECT 100.530 109.490 101.480 109.520 ;
        RECT 97.440 107.860 97.770 108.640 ;
        RECT 98.970 108.560 99.920 109.320 ;
      LAYER li1 ;
        RECT 100.100 108.680 100.350 109.390 ;
      LAYER li1 ;
        RECT 100.530 109.320 100.560 109.490 ;
        RECT 100.730 109.320 100.920 109.490 ;
        RECT 101.090 109.320 101.280 109.490 ;
        RECT 101.450 109.320 101.480 109.490 ;
        RECT 102.090 109.490 103.040 109.520 ;
        RECT 100.530 108.860 101.480 109.320 ;
      LAYER li1 ;
        RECT 101.660 108.680 101.910 109.390 ;
        RECT 100.100 108.510 101.910 108.680 ;
      LAYER li1 ;
        RECT 102.090 109.320 102.120 109.490 ;
        RECT 102.290 109.320 102.480 109.490 ;
        RECT 102.650 109.320 102.840 109.490 ;
        RECT 103.010 109.320 103.040 109.490 ;
        RECT 103.850 109.490 105.460 109.520 ;
        RECT 102.090 108.640 103.040 109.320 ;
      LAYER li1 ;
        RECT 100.100 108.340 100.270 108.510 ;
      LAYER li1 ;
        RECT 103.220 108.460 103.550 109.390 ;
        RECT 103.850 109.320 103.900 109.490 ;
        RECT 104.070 109.320 104.340 109.490 ;
        RECT 104.510 109.320 104.780 109.490 ;
        RECT 104.950 109.320 105.190 109.490 ;
        RECT 105.360 109.320 105.460 109.490 ;
        RECT 103.850 109.040 105.460 109.320 ;
        RECT 97.980 107.200 98.310 108.190 ;
      LAYER li1 ;
        RECT 99.010 108.110 100.270 108.340 ;
      LAYER li1 ;
        RECT 102.310 108.330 103.550 108.460 ;
        RECT 100.450 108.290 103.550 108.330 ;
        RECT 100.450 108.160 102.480 108.290 ;
      LAYER li1 ;
        RECT 100.100 107.980 100.270 108.110 ;
        RECT 100.100 107.810 101.990 107.980 ;
      LAYER li1 ;
        RECT 97.210 106.330 98.660 107.200 ;
        RECT 97.210 106.160 97.460 106.330 ;
        RECT 97.630 106.160 97.820 106.330 ;
        RECT 97.990 106.160 98.260 106.330 ;
        RECT 98.430 106.160 98.660 106.330 ;
        RECT 97.210 106.130 98.660 106.160 ;
        RECT 98.970 106.380 99.920 107.710 ;
        RECT 98.970 106.210 99.000 106.380 ;
        RECT 99.170 106.210 99.360 106.380 ;
        RECT 99.530 106.210 99.720 106.380 ;
        RECT 99.890 106.210 99.920 106.380 ;
        RECT 98.970 106.130 99.920 106.210 ;
      LAYER li1 ;
        RECT 100.100 106.130 100.350 107.810 ;
      LAYER li1 ;
        RECT 100.530 106.380 101.480 107.630 ;
        RECT 100.530 106.210 100.560 106.380 ;
        RECT 100.730 106.210 100.920 106.380 ;
        RECT 101.090 106.210 101.280 106.380 ;
        RECT 101.450 106.210 101.480 106.380 ;
        RECT 100.530 106.130 101.480 106.210 ;
      LAYER li1 ;
        RECT 101.660 106.130 101.990 107.810 ;
        RECT 102.770 107.770 103.100 108.110 ;
      LAYER li1 ;
        RECT 102.170 106.380 103.120 107.590 ;
        RECT 102.170 106.210 102.200 106.380 ;
        RECT 102.370 106.210 102.560 106.380 ;
        RECT 102.730 106.210 102.920 106.380 ;
        RECT 103.090 106.210 103.120 106.380 ;
        RECT 102.170 106.130 103.120 106.210 ;
        RECT 103.300 106.130 103.550 108.290 ;
        RECT 104.160 108.640 105.460 109.040 ;
        RECT 105.690 109.490 106.640 109.520 ;
        RECT 105.690 109.320 105.720 109.490 ;
        RECT 105.890 109.320 106.080 109.490 ;
        RECT 106.250 109.320 106.440 109.490 ;
        RECT 106.610 109.320 106.640 109.490 ;
        RECT 107.250 109.490 108.200 109.520 ;
        RECT 104.160 107.860 104.490 108.640 ;
        RECT 105.690 108.560 106.640 109.320 ;
      LAYER li1 ;
        RECT 106.820 108.680 107.070 109.390 ;
      LAYER li1 ;
        RECT 107.250 109.320 107.280 109.490 ;
        RECT 107.450 109.320 107.640 109.490 ;
        RECT 107.810 109.320 108.000 109.490 ;
        RECT 108.170 109.320 108.200 109.490 ;
        RECT 108.810 109.490 109.760 109.520 ;
        RECT 107.250 108.860 108.200 109.320 ;
      LAYER li1 ;
        RECT 108.380 108.680 108.630 109.390 ;
        RECT 106.820 108.510 108.630 108.680 ;
      LAYER li1 ;
        RECT 108.810 109.320 108.840 109.490 ;
        RECT 109.010 109.320 109.200 109.490 ;
        RECT 109.370 109.320 109.560 109.490 ;
        RECT 109.730 109.320 109.760 109.490 ;
        RECT 110.570 109.490 112.180 109.520 ;
        RECT 112.870 109.490 114.120 109.520 ;
        RECT 114.890 109.490 116.500 109.520 ;
        RECT 117.670 109.490 118.920 109.520 ;
        RECT 119.690 109.490 121.300 109.520 ;
        RECT 108.810 108.640 109.760 109.320 ;
      LAYER li1 ;
        RECT 106.820 108.340 106.990 108.510 ;
      LAYER li1 ;
        RECT 109.940 108.460 110.270 109.390 ;
        RECT 110.570 109.320 110.620 109.490 ;
        RECT 110.790 109.320 111.060 109.490 ;
        RECT 111.230 109.320 111.500 109.490 ;
        RECT 111.670 109.320 111.910 109.490 ;
        RECT 112.080 109.320 112.180 109.490 ;
        RECT 110.570 109.040 112.180 109.320 ;
        RECT 104.700 107.200 105.030 108.190 ;
      LAYER li1 ;
        RECT 105.730 108.110 106.990 108.340 ;
      LAYER li1 ;
        RECT 109.030 108.330 110.270 108.460 ;
        RECT 107.170 108.290 110.270 108.330 ;
        RECT 107.170 108.160 109.200 108.290 ;
      LAYER li1 ;
        RECT 106.820 107.980 106.990 108.110 ;
        RECT 106.820 107.810 108.710 107.980 ;
      LAYER li1 ;
        RECT 103.930 106.330 105.380 107.200 ;
        RECT 103.930 106.160 104.180 106.330 ;
        RECT 104.350 106.160 104.540 106.330 ;
        RECT 104.710 106.160 104.980 106.330 ;
        RECT 105.150 106.160 105.380 106.330 ;
        RECT 103.930 106.130 105.380 106.160 ;
        RECT 105.690 106.380 106.640 107.710 ;
        RECT 105.690 106.210 105.720 106.380 ;
        RECT 105.890 106.210 106.080 106.380 ;
        RECT 106.250 106.210 106.440 106.380 ;
        RECT 106.610 106.210 106.640 106.380 ;
        RECT 105.690 106.130 106.640 106.210 ;
      LAYER li1 ;
        RECT 106.820 106.130 107.070 107.810 ;
      LAYER li1 ;
        RECT 107.250 106.380 108.200 107.630 ;
        RECT 107.250 106.210 107.280 106.380 ;
        RECT 107.450 106.210 107.640 106.380 ;
        RECT 107.810 106.210 108.000 106.380 ;
        RECT 108.170 106.210 108.200 106.380 ;
        RECT 107.250 106.130 108.200 106.210 ;
      LAYER li1 ;
        RECT 108.380 106.130 108.710 107.810 ;
        RECT 109.490 107.770 109.820 108.110 ;
      LAYER li1 ;
        RECT 108.890 106.380 109.840 107.590 ;
        RECT 108.890 106.210 108.920 106.380 ;
        RECT 109.090 106.210 109.280 106.380 ;
        RECT 109.450 106.210 109.640 106.380 ;
        RECT 109.810 106.210 109.840 106.380 ;
        RECT 108.890 106.130 109.840 106.210 ;
        RECT 110.020 106.130 110.270 108.290 ;
        RECT 110.880 108.640 112.180 109.040 ;
        RECT 110.880 107.860 111.210 108.640 ;
        RECT 111.420 107.200 111.750 108.190 ;
      LAYER li1 ;
        RECT 112.440 107.710 112.690 109.390 ;
      LAYER li1 ;
        RECT 113.040 109.320 113.230 109.490 ;
        RECT 113.400 109.320 113.590 109.490 ;
        RECT 113.760 109.320 113.950 109.490 ;
        RECT 112.870 108.950 114.120 109.320 ;
        RECT 114.300 108.770 114.550 109.390 ;
        RECT 114.890 109.320 114.940 109.490 ;
        RECT 115.110 109.320 115.380 109.490 ;
        RECT 115.550 109.320 115.820 109.490 ;
        RECT 115.990 109.320 116.230 109.490 ;
        RECT 116.400 109.320 116.500 109.490 ;
        RECT 114.890 109.040 116.500 109.320 ;
        RECT 113.000 108.600 114.550 108.770 ;
        RECT 113.000 108.140 113.330 108.600 ;
        RECT 110.650 106.330 112.100 107.200 ;
        RECT 110.650 106.160 110.900 106.330 ;
        RECT 111.070 106.160 111.260 106.330 ;
        RECT 111.430 106.160 111.700 106.330 ;
        RECT 111.870 106.160 112.100 106.330 ;
        RECT 110.650 106.130 112.100 106.160 ;
      LAYER li1 ;
        RECT 112.440 106.130 112.870 107.710 ;
      LAYER li1 ;
        RECT 113.050 106.380 113.610 107.710 ;
      LAYER li1 ;
        RECT 113.790 106.630 114.120 108.420 ;
      LAYER li1 ;
        RECT 114.300 106.880 114.550 108.600 ;
        RECT 115.200 108.640 116.500 109.040 ;
        RECT 115.200 107.860 115.530 108.640 ;
        RECT 115.740 107.200 116.070 108.190 ;
      LAYER li1 ;
        RECT 117.240 107.710 117.490 109.390 ;
      LAYER li1 ;
        RECT 117.840 109.320 118.030 109.490 ;
        RECT 118.200 109.320 118.390 109.490 ;
        RECT 118.560 109.320 118.750 109.490 ;
        RECT 117.670 108.950 118.920 109.320 ;
        RECT 119.100 108.770 119.350 109.390 ;
        RECT 119.690 109.320 119.740 109.490 ;
        RECT 119.910 109.320 120.180 109.490 ;
        RECT 120.350 109.320 120.620 109.490 ;
        RECT 120.790 109.320 121.030 109.490 ;
        RECT 121.200 109.320 121.300 109.490 ;
        RECT 119.690 109.040 121.300 109.320 ;
        RECT 117.800 108.600 119.350 108.770 ;
        RECT 117.800 108.140 118.130 108.600 ;
        RECT 113.050 106.210 113.060 106.380 ;
        RECT 113.230 106.210 113.420 106.380 ;
        RECT 113.590 106.210 113.610 106.380 ;
        RECT 113.050 106.130 113.610 106.210 ;
        RECT 114.970 106.330 116.420 107.200 ;
        RECT 114.970 106.160 115.220 106.330 ;
        RECT 115.390 106.160 115.580 106.330 ;
        RECT 115.750 106.160 116.020 106.330 ;
        RECT 116.190 106.160 116.420 106.330 ;
        RECT 114.970 106.130 116.420 106.160 ;
      LAYER li1 ;
        RECT 117.240 106.130 117.670 107.710 ;
      LAYER li1 ;
        RECT 117.850 106.380 118.410 107.710 ;
      LAYER li1 ;
        RECT 118.590 106.630 118.920 108.420 ;
      LAYER li1 ;
        RECT 119.100 106.880 119.350 108.600 ;
        RECT 120.000 108.640 121.300 109.040 ;
        RECT 121.530 109.490 122.480 109.520 ;
        RECT 121.530 109.320 121.560 109.490 ;
        RECT 121.730 109.320 121.920 109.490 ;
        RECT 122.090 109.320 122.280 109.490 ;
        RECT 122.450 109.320 122.480 109.490 ;
        RECT 123.090 109.490 124.040 109.520 ;
        RECT 120.000 107.860 120.330 108.640 ;
        RECT 121.530 108.560 122.480 109.320 ;
      LAYER li1 ;
        RECT 122.660 108.680 122.910 109.390 ;
      LAYER li1 ;
        RECT 123.090 109.320 123.120 109.490 ;
        RECT 123.290 109.320 123.480 109.490 ;
        RECT 123.650 109.320 123.840 109.490 ;
        RECT 124.010 109.320 124.040 109.490 ;
        RECT 124.650 109.490 125.600 109.520 ;
        RECT 123.090 108.860 124.040 109.320 ;
      LAYER li1 ;
        RECT 124.220 108.680 124.470 109.390 ;
        RECT 122.660 108.510 124.470 108.680 ;
      LAYER li1 ;
        RECT 124.650 109.320 124.680 109.490 ;
        RECT 124.850 109.320 125.040 109.490 ;
        RECT 125.210 109.320 125.400 109.490 ;
        RECT 125.570 109.320 125.600 109.490 ;
        RECT 126.820 109.500 129.550 109.530 ;
        RECT 124.650 108.640 125.600 109.320 ;
      LAYER li1 ;
        RECT 122.660 108.340 122.830 108.510 ;
      LAYER li1 ;
        RECT 125.780 108.460 126.110 109.390 ;
        RECT 126.820 109.330 126.990 109.500 ;
        RECT 127.160 109.330 127.430 109.500 ;
        RECT 127.600 109.330 127.840 109.500 ;
        RECT 128.010 109.330 128.270 109.500 ;
        RECT 128.440 109.330 128.710 109.500 ;
        RECT 128.880 109.330 129.120 109.500 ;
        RECT 129.290 109.330 129.550 109.500 ;
        RECT 126.820 108.530 129.550 109.330 ;
        RECT 130.660 109.500 133.390 109.530 ;
        RECT 130.660 109.330 130.830 109.500 ;
        RECT 131.000 109.330 131.270 109.500 ;
        RECT 131.440 109.330 131.680 109.500 ;
        RECT 131.850 109.330 132.110 109.500 ;
        RECT 132.280 109.330 132.550 109.500 ;
        RECT 132.720 109.330 132.960 109.500 ;
        RECT 133.130 109.330 133.390 109.500 ;
        RECT 130.660 108.530 133.390 109.330 ;
        RECT 134.500 109.500 137.230 109.530 ;
        RECT 134.500 109.330 134.670 109.500 ;
        RECT 134.840 109.330 135.110 109.500 ;
        RECT 135.280 109.330 135.520 109.500 ;
        RECT 135.690 109.330 135.950 109.500 ;
        RECT 136.120 109.330 136.390 109.500 ;
        RECT 136.560 109.330 136.800 109.500 ;
        RECT 136.970 109.330 137.230 109.500 ;
        RECT 134.500 108.530 137.230 109.330 ;
        RECT 138.340 109.500 141.070 109.530 ;
        RECT 138.340 109.330 138.510 109.500 ;
        RECT 138.680 109.330 138.950 109.500 ;
        RECT 139.120 109.330 139.360 109.500 ;
        RECT 139.530 109.330 139.790 109.500 ;
        RECT 139.960 109.330 140.230 109.500 ;
        RECT 140.400 109.330 140.640 109.500 ;
        RECT 140.810 109.330 141.070 109.500 ;
        RECT 138.340 108.530 141.070 109.330 ;
        RECT 120.540 107.200 120.870 108.190 ;
      LAYER li1 ;
        RECT 121.570 108.110 122.830 108.340 ;
      LAYER li1 ;
        RECT 124.870 108.330 126.110 108.460 ;
        RECT 123.010 108.290 126.110 108.330 ;
        RECT 123.010 108.160 125.040 108.290 ;
      LAYER li1 ;
        RECT 122.660 107.980 122.830 108.110 ;
        RECT 122.660 107.810 124.550 107.980 ;
      LAYER li1 ;
        RECT 117.850 106.210 117.860 106.380 ;
        RECT 118.030 106.210 118.220 106.380 ;
        RECT 118.390 106.210 118.410 106.380 ;
        RECT 117.850 106.130 118.410 106.210 ;
        RECT 119.770 106.330 121.220 107.200 ;
        RECT 119.770 106.160 120.020 106.330 ;
        RECT 120.190 106.160 120.380 106.330 ;
        RECT 120.550 106.160 120.820 106.330 ;
        RECT 120.990 106.160 121.220 106.330 ;
        RECT 119.770 106.130 121.220 106.160 ;
        RECT 121.530 106.380 122.480 107.710 ;
        RECT 121.530 106.210 121.560 106.380 ;
        RECT 121.730 106.210 121.920 106.380 ;
        RECT 122.090 106.210 122.280 106.380 ;
        RECT 122.450 106.210 122.480 106.380 ;
        RECT 121.530 106.130 122.480 106.210 ;
      LAYER li1 ;
        RECT 122.660 106.130 122.910 107.810 ;
      LAYER li1 ;
        RECT 123.090 106.380 124.040 107.630 ;
        RECT 123.090 106.210 123.120 106.380 ;
        RECT 123.290 106.210 123.480 106.380 ;
        RECT 123.650 106.210 123.840 106.380 ;
        RECT 124.010 106.210 124.040 106.380 ;
        RECT 123.090 106.130 124.040 106.210 ;
      LAYER li1 ;
        RECT 124.220 106.130 124.550 107.810 ;
        RECT 125.330 107.770 125.660 108.110 ;
      LAYER li1 ;
        RECT 124.730 106.380 125.680 107.590 ;
        RECT 124.730 106.210 124.760 106.380 ;
        RECT 124.930 106.210 125.120 106.380 ;
        RECT 125.290 106.210 125.480 106.380 ;
        RECT 125.650 106.210 125.680 106.380 ;
        RECT 124.730 106.130 125.680 106.210 ;
        RECT 125.860 106.130 126.110 108.290 ;
        RECT 126.980 107.860 127.310 108.530 ;
        RECT 127.710 107.210 128.040 108.190 ;
        RECT 128.260 107.860 128.590 108.530 ;
        RECT 128.990 107.210 129.320 108.190 ;
        RECT 130.820 107.860 131.150 108.530 ;
        RECT 131.550 107.210 131.880 108.190 ;
        RECT 132.100 107.860 132.430 108.530 ;
        RECT 132.830 107.210 133.160 108.190 ;
        RECT 134.660 107.860 134.990 108.530 ;
        RECT 135.390 107.210 135.720 108.190 ;
        RECT 135.940 107.860 136.270 108.530 ;
        RECT 136.670 107.210 137.000 108.190 ;
        RECT 138.500 107.860 138.830 108.530 ;
        RECT 139.230 107.210 139.560 108.190 ;
        RECT 139.780 107.860 140.110 108.530 ;
        RECT 140.510 107.210 140.840 108.190 ;
        RECT 126.740 106.330 129.480 107.210 ;
        RECT 126.740 106.160 126.950 106.330 ;
        RECT 127.120 106.160 127.390 106.330 ;
        RECT 127.560 106.160 127.800 106.330 ;
        RECT 127.970 106.160 128.230 106.330 ;
        RECT 128.400 106.160 128.670 106.330 ;
        RECT 128.840 106.160 129.080 106.330 ;
        RECT 129.250 106.160 129.480 106.330 ;
        RECT 126.740 106.140 129.480 106.160 ;
        RECT 130.580 106.330 133.320 107.210 ;
        RECT 130.580 106.160 130.790 106.330 ;
        RECT 130.960 106.160 131.230 106.330 ;
        RECT 131.400 106.160 131.640 106.330 ;
        RECT 131.810 106.160 132.070 106.330 ;
        RECT 132.240 106.160 132.510 106.330 ;
        RECT 132.680 106.160 132.920 106.330 ;
        RECT 133.090 106.160 133.320 106.330 ;
        RECT 130.580 106.140 133.320 106.160 ;
        RECT 134.420 106.330 137.160 107.210 ;
        RECT 134.420 106.160 134.630 106.330 ;
        RECT 134.800 106.160 135.070 106.330 ;
        RECT 135.240 106.160 135.480 106.330 ;
        RECT 135.650 106.160 135.910 106.330 ;
        RECT 136.080 106.160 136.350 106.330 ;
        RECT 136.520 106.160 136.760 106.330 ;
        RECT 136.930 106.160 137.160 106.330 ;
        RECT 134.420 106.140 137.160 106.160 ;
        RECT 138.260 106.330 141.000 107.210 ;
        RECT 138.260 106.160 138.470 106.330 ;
        RECT 138.640 106.160 138.910 106.330 ;
        RECT 139.080 106.160 139.320 106.330 ;
        RECT 139.490 106.160 139.750 106.330 ;
        RECT 139.920 106.160 140.190 106.330 ;
        RECT 140.360 106.160 140.600 106.330 ;
        RECT 140.770 106.160 141.000 106.330 ;
        RECT 138.260 106.140 141.000 106.160 ;
        RECT 5.760 105.730 5.920 105.910 ;
        RECT 6.090 105.730 6.400 105.910 ;
        RECT 6.570 105.730 6.880 105.910 ;
        RECT 7.050 105.730 7.360 105.910 ;
        RECT 7.530 105.730 7.840 105.910 ;
        RECT 8.010 105.730 8.320 105.910 ;
        RECT 8.490 105.730 8.800 105.910 ;
        RECT 8.970 105.730 9.280 105.910 ;
        RECT 9.450 105.730 9.760 105.910 ;
        RECT 9.930 105.730 10.240 105.910 ;
        RECT 10.410 105.730 10.720 105.910 ;
        RECT 10.890 105.730 11.200 105.910 ;
        RECT 11.370 105.730 11.680 105.910 ;
        RECT 11.850 105.730 12.160 105.910 ;
        RECT 12.330 105.730 12.640 105.910 ;
        RECT 12.810 105.730 13.120 105.910 ;
        RECT 13.290 105.730 13.600 105.910 ;
        RECT 13.770 105.730 14.080 105.910 ;
        RECT 14.250 105.730 14.560 105.910 ;
        RECT 14.730 105.730 15.040 105.910 ;
        RECT 15.210 105.730 15.520 105.910 ;
        RECT 15.690 105.730 16.000 105.910 ;
        RECT 16.170 105.730 16.480 105.910 ;
        RECT 16.650 105.730 16.960 105.910 ;
        RECT 17.130 105.730 17.440 105.910 ;
        RECT 17.610 105.730 17.920 105.910 ;
        RECT 18.090 105.730 18.400 105.910 ;
        RECT 18.570 105.730 18.880 105.910 ;
        RECT 19.050 105.730 19.360 105.910 ;
        RECT 19.530 105.730 19.840 105.910 ;
        RECT 20.010 105.730 20.320 105.910 ;
        RECT 20.490 105.730 20.800 105.910 ;
        RECT 20.970 105.730 21.280 105.910 ;
        RECT 21.450 105.730 21.760 105.910 ;
        RECT 21.930 105.730 22.240 105.910 ;
        RECT 22.410 105.730 22.720 105.910 ;
        RECT 22.890 105.730 23.200 105.910 ;
        RECT 23.370 105.730 23.680 105.910 ;
        RECT 23.850 105.730 24.160 105.910 ;
        RECT 24.330 105.730 24.640 105.910 ;
        RECT 24.810 105.730 25.120 105.910 ;
        RECT 25.290 105.730 25.600 105.910 ;
        RECT 25.770 105.730 26.080 105.910 ;
        RECT 26.250 105.730 26.560 105.910 ;
        RECT 26.730 105.730 27.040 105.910 ;
        RECT 27.210 105.730 27.520 105.910 ;
        RECT 27.690 105.730 28.000 105.910 ;
        RECT 28.170 105.730 28.480 105.910 ;
        RECT 28.650 105.730 28.960 105.910 ;
        RECT 29.130 105.730 29.440 105.910 ;
        RECT 29.610 105.730 29.920 105.910 ;
        RECT 30.090 105.730 30.400 105.910 ;
        RECT 30.570 105.730 30.880 105.910 ;
        RECT 31.050 105.730 31.360 105.910 ;
        RECT 31.530 105.730 31.840 105.910 ;
        RECT 32.010 105.730 32.320 105.910 ;
        RECT 32.490 105.730 32.800 105.910 ;
        RECT 32.970 105.730 33.280 105.910 ;
        RECT 33.450 105.730 33.760 105.910 ;
        RECT 33.930 105.730 34.240 105.910 ;
        RECT 34.410 105.730 34.720 105.910 ;
        RECT 34.890 105.730 35.200 105.910 ;
        RECT 35.370 105.730 35.680 105.910 ;
        RECT 35.850 105.730 36.160 105.910 ;
        RECT 36.330 105.730 36.640 105.910 ;
        RECT 36.810 105.730 37.120 105.910 ;
        RECT 37.290 105.730 37.600 105.910 ;
        RECT 37.770 105.730 38.080 105.910 ;
        RECT 38.250 105.730 38.560 105.910 ;
        RECT 38.730 105.730 39.040 105.910 ;
        RECT 39.210 105.730 39.520 105.910 ;
        RECT 39.690 105.730 40.000 105.910 ;
        RECT 40.170 105.900 40.320 105.910 ;
        RECT 40.800 105.900 40.960 105.910 ;
        RECT 40.170 105.730 40.480 105.900 ;
        RECT 40.650 105.730 40.960 105.900 ;
        RECT 41.130 105.730 41.440 105.910 ;
        RECT 41.610 105.730 41.920 105.910 ;
        RECT 42.090 105.730 42.400 105.910 ;
        RECT 42.570 105.730 42.880 105.910 ;
        RECT 43.050 105.730 43.360 105.910 ;
        RECT 43.530 105.730 43.840 105.910 ;
        RECT 44.010 105.730 44.320 105.910 ;
        RECT 44.490 105.730 44.800 105.910 ;
        RECT 44.970 105.730 45.280 105.910 ;
        RECT 45.450 105.730 45.760 105.910 ;
        RECT 45.930 105.730 46.240 105.910 ;
        RECT 46.410 105.730 46.720 105.910 ;
        RECT 46.890 105.730 47.200 105.910 ;
        RECT 47.370 105.730 47.680 105.910 ;
        RECT 47.850 105.730 48.160 105.910 ;
        RECT 48.330 105.730 48.640 105.910 ;
        RECT 48.810 105.730 49.120 105.910 ;
        RECT 49.290 105.730 49.600 105.910 ;
        RECT 49.770 105.730 50.080 105.910 ;
        RECT 50.250 105.730 50.560 105.910 ;
        RECT 50.730 105.730 51.040 105.910 ;
        RECT 51.210 105.730 51.520 105.910 ;
        RECT 51.690 105.730 52.000 105.910 ;
        RECT 52.170 105.730 52.480 105.910 ;
        RECT 52.650 105.730 52.960 105.910 ;
        RECT 53.130 105.730 53.440 105.910 ;
        RECT 53.610 105.730 53.920 105.910 ;
        RECT 54.090 105.730 54.400 105.910 ;
        RECT 54.570 105.730 54.880 105.910 ;
        RECT 55.050 105.730 55.360 105.910 ;
        RECT 55.530 105.730 55.840 105.910 ;
        RECT 56.010 105.730 56.320 105.910 ;
        RECT 56.490 105.730 56.800 105.910 ;
        RECT 56.970 105.730 57.280 105.910 ;
        RECT 57.450 105.730 57.760 105.910 ;
        RECT 57.930 105.730 58.240 105.910 ;
        RECT 58.410 105.730 58.720 105.910 ;
        RECT 58.890 105.730 59.200 105.910 ;
        RECT 59.370 105.730 59.680 105.910 ;
        RECT 59.850 105.730 60.160 105.910 ;
        RECT 60.330 105.730 60.640 105.910 ;
        RECT 60.810 105.900 60.960 105.910 ;
        RECT 61.440 105.900 61.600 105.910 ;
        RECT 60.810 105.730 61.120 105.900 ;
        RECT 61.290 105.730 61.600 105.900 ;
        RECT 61.770 105.730 62.080 105.910 ;
        RECT 62.250 105.730 62.560 105.910 ;
        RECT 62.730 105.730 63.040 105.910 ;
        RECT 63.210 105.730 63.520 105.910 ;
        RECT 63.690 105.730 64.000 105.910 ;
        RECT 64.170 105.730 64.480 105.910 ;
        RECT 64.650 105.730 64.960 105.910 ;
        RECT 65.130 105.730 65.440 105.910 ;
        RECT 65.610 105.730 65.920 105.910 ;
        RECT 66.090 105.730 66.400 105.910 ;
        RECT 66.570 105.730 66.880 105.910 ;
        RECT 67.050 105.730 67.360 105.910 ;
        RECT 67.530 105.730 67.840 105.910 ;
        RECT 68.010 105.730 68.320 105.910 ;
        RECT 68.490 105.730 68.800 105.910 ;
        RECT 68.970 105.730 69.280 105.910 ;
        RECT 69.450 105.730 69.760 105.910 ;
        RECT 69.930 105.730 70.240 105.910 ;
        RECT 70.410 105.730 70.720 105.910 ;
        RECT 70.890 105.730 71.200 105.910 ;
        RECT 71.370 105.730 71.680 105.910 ;
        RECT 71.850 105.730 72.160 105.910 ;
        RECT 72.330 105.730 72.640 105.910 ;
        RECT 72.810 105.730 73.120 105.910 ;
        RECT 73.290 105.900 73.600 105.910 ;
        RECT 73.770 105.900 74.080 105.910 ;
        RECT 73.290 105.730 73.440 105.900 ;
        RECT 73.920 105.730 74.080 105.900 ;
        RECT 74.250 105.730 74.560 105.910 ;
        RECT 74.730 105.730 75.040 105.910 ;
        RECT 75.210 105.730 75.520 105.910 ;
        RECT 75.690 105.730 76.000 105.910 ;
        RECT 76.170 105.730 76.480 105.910 ;
        RECT 76.650 105.730 76.960 105.910 ;
        RECT 77.130 105.730 77.440 105.910 ;
        RECT 77.610 105.730 77.920 105.910 ;
        RECT 78.090 105.730 78.400 105.910 ;
        RECT 78.570 105.730 78.880 105.910 ;
        RECT 79.050 105.730 79.360 105.910 ;
        RECT 79.530 105.730 79.840 105.910 ;
        RECT 80.010 105.730 80.320 105.910 ;
        RECT 80.490 105.730 80.800 105.910 ;
        RECT 80.970 105.730 81.280 105.910 ;
        RECT 81.450 105.730 81.760 105.910 ;
        RECT 81.930 105.730 82.240 105.910 ;
        RECT 82.410 105.730 82.720 105.910 ;
        RECT 82.890 105.730 83.200 105.910 ;
        RECT 83.370 105.730 83.680 105.910 ;
        RECT 83.850 105.730 84.160 105.910 ;
        RECT 84.330 105.730 84.640 105.910 ;
        RECT 84.810 105.730 85.120 105.910 ;
        RECT 85.290 105.730 85.600 105.910 ;
        RECT 85.770 105.730 86.080 105.910 ;
        RECT 86.250 105.730 86.560 105.910 ;
        RECT 86.730 105.730 87.040 105.910 ;
        RECT 87.210 105.730 87.520 105.910 ;
        RECT 87.690 105.730 88.000 105.910 ;
        RECT 88.170 105.730 88.480 105.910 ;
        RECT 88.650 105.730 88.960 105.910 ;
        RECT 89.130 105.730 89.440 105.910 ;
        RECT 89.610 105.730 89.920 105.910 ;
        RECT 90.090 105.730 90.400 105.910 ;
        RECT 90.570 105.730 90.880 105.910 ;
        RECT 91.050 105.730 91.360 105.910 ;
        RECT 91.530 105.730 91.840 105.910 ;
        RECT 92.010 105.730 92.320 105.910 ;
        RECT 92.490 105.730 92.800 105.910 ;
        RECT 92.970 105.730 93.280 105.910 ;
        RECT 93.450 105.730 93.760 105.910 ;
        RECT 93.930 105.730 94.240 105.910 ;
        RECT 94.410 105.730 94.720 105.910 ;
        RECT 94.890 105.730 95.200 105.910 ;
        RECT 95.370 105.730 95.680 105.910 ;
        RECT 95.850 105.730 96.160 105.910 ;
        RECT 96.330 105.730 96.640 105.910 ;
        RECT 96.810 105.730 97.120 105.910 ;
        RECT 97.290 105.730 97.600 105.910 ;
        RECT 97.770 105.730 98.080 105.910 ;
        RECT 98.250 105.730 98.560 105.910 ;
        RECT 98.730 105.730 99.040 105.910 ;
        RECT 99.210 105.730 99.520 105.910 ;
        RECT 99.690 105.730 100.000 105.910 ;
        RECT 100.170 105.730 100.480 105.910 ;
        RECT 100.650 105.730 100.960 105.910 ;
        RECT 101.130 105.730 101.440 105.910 ;
        RECT 101.610 105.730 101.920 105.910 ;
        RECT 102.090 105.730 102.400 105.910 ;
        RECT 102.570 105.730 102.880 105.910 ;
        RECT 103.050 105.730 103.360 105.910 ;
        RECT 103.530 105.730 103.840 105.910 ;
        RECT 104.010 105.730 104.320 105.910 ;
        RECT 104.490 105.730 104.800 105.910 ;
        RECT 104.970 105.730 105.280 105.910 ;
        RECT 105.450 105.730 105.760 105.910 ;
        RECT 105.930 105.730 106.240 105.910 ;
        RECT 106.410 105.730 106.720 105.910 ;
        RECT 106.890 105.730 107.200 105.910 ;
        RECT 107.370 105.730 107.680 105.910 ;
        RECT 107.850 105.730 108.160 105.910 ;
        RECT 108.330 105.730 108.640 105.910 ;
        RECT 108.810 105.730 109.120 105.910 ;
        RECT 109.290 105.730 109.600 105.910 ;
        RECT 109.770 105.730 110.080 105.910 ;
        RECT 110.250 105.730 110.560 105.910 ;
        RECT 110.730 105.730 111.040 105.910 ;
        RECT 111.210 105.730 111.520 105.910 ;
        RECT 111.690 105.730 112.000 105.910 ;
        RECT 112.170 105.730 112.480 105.910 ;
        RECT 112.650 105.730 112.960 105.910 ;
        RECT 113.130 105.730 113.440 105.910 ;
        RECT 113.610 105.730 113.920 105.910 ;
        RECT 114.090 105.730 114.400 105.910 ;
        RECT 114.570 105.730 114.880 105.910 ;
        RECT 115.050 105.730 115.360 105.910 ;
        RECT 115.530 105.730 115.840 105.910 ;
        RECT 116.010 105.730 116.320 105.910 ;
        RECT 116.490 105.900 116.800 105.910 ;
        RECT 116.970 105.900 117.280 105.910 ;
        RECT 116.490 105.730 116.640 105.900 ;
        RECT 117.120 105.730 117.280 105.900 ;
        RECT 117.450 105.730 117.760 105.910 ;
        RECT 117.930 105.730 118.240 105.910 ;
        RECT 118.410 105.730 118.720 105.910 ;
        RECT 118.890 105.730 119.200 105.910 ;
        RECT 119.370 105.730 119.680 105.910 ;
        RECT 119.850 105.730 120.160 105.910 ;
        RECT 120.330 105.730 120.640 105.910 ;
        RECT 120.810 105.900 120.960 105.910 ;
        RECT 121.440 105.900 121.600 105.910 ;
        RECT 120.810 105.730 121.120 105.900 ;
        RECT 121.290 105.730 121.600 105.900 ;
        RECT 121.770 105.730 122.080 105.910 ;
        RECT 122.250 105.730 122.560 105.910 ;
        RECT 122.730 105.730 123.040 105.910 ;
        RECT 123.210 105.730 123.520 105.910 ;
        RECT 123.690 105.730 124.000 105.910 ;
        RECT 124.170 105.730 124.480 105.910 ;
        RECT 124.650 105.730 124.960 105.910 ;
        RECT 125.130 105.730 125.440 105.910 ;
        RECT 125.610 105.730 125.920 105.910 ;
        RECT 126.090 105.730 126.400 105.910 ;
        RECT 126.570 105.730 126.880 105.910 ;
        RECT 127.050 105.730 127.360 105.910 ;
        RECT 127.530 105.730 127.840 105.910 ;
        RECT 128.010 105.730 128.320 105.910 ;
        RECT 128.490 105.730 128.800 105.910 ;
        RECT 128.970 105.730 129.280 105.910 ;
        RECT 129.450 105.730 129.760 105.910 ;
        RECT 129.930 105.730 130.240 105.910 ;
        RECT 130.410 105.730 130.720 105.910 ;
        RECT 130.890 105.730 131.200 105.910 ;
        RECT 131.370 105.730 131.680 105.910 ;
        RECT 131.850 105.730 132.160 105.910 ;
        RECT 132.330 105.730 132.640 105.910 ;
        RECT 132.810 105.730 133.120 105.910 ;
        RECT 133.290 105.730 133.600 105.910 ;
        RECT 133.770 105.730 134.080 105.910 ;
        RECT 134.250 105.730 134.560 105.910 ;
        RECT 134.730 105.730 135.040 105.910 ;
        RECT 135.210 105.730 135.520 105.910 ;
        RECT 135.690 105.730 136.000 105.910 ;
        RECT 136.170 105.730 136.480 105.910 ;
        RECT 136.650 105.730 136.960 105.910 ;
        RECT 137.130 105.730 137.440 105.910 ;
        RECT 137.610 105.730 137.920 105.910 ;
        RECT 138.090 105.730 138.400 105.910 ;
        RECT 138.570 105.730 138.880 105.910 ;
        RECT 139.050 105.730 139.360 105.910 ;
        RECT 139.530 105.730 139.840 105.910 ;
        RECT 140.010 105.730 140.320 105.910 ;
        RECT 140.490 105.730 140.800 105.910 ;
        RECT 140.970 105.730 141.280 105.910 ;
        RECT 141.450 105.900 141.760 105.910 ;
        RECT 141.930 105.900 142.080 105.910 ;
        RECT 141.450 105.730 141.600 105.900 ;
        RECT 6.260 105.480 9.000 105.500 ;
        RECT 6.260 105.310 6.470 105.480 ;
        RECT 6.640 105.310 6.910 105.480 ;
        RECT 7.080 105.310 7.320 105.480 ;
        RECT 7.490 105.310 7.750 105.480 ;
        RECT 7.920 105.310 8.190 105.480 ;
        RECT 8.360 105.310 8.600 105.480 ;
        RECT 8.770 105.310 9.000 105.480 ;
        RECT 6.260 104.430 9.000 105.310 ;
        RECT 10.230 105.430 10.820 105.460 ;
        RECT 10.230 105.260 10.260 105.430 ;
        RECT 10.430 105.260 10.620 105.430 ;
        RECT 10.790 105.260 10.820 105.430 ;
        RECT 6.500 103.110 6.830 103.780 ;
        RECT 7.230 103.450 7.560 104.430 ;
        RECT 7.780 103.110 8.110 103.780 ;
        RECT 8.510 103.450 8.840 104.430 ;
        RECT 9.710 104.280 10.040 105.210 ;
        RECT 10.230 104.480 10.820 105.260 ;
        RECT 11.000 105.390 12.440 105.560 ;
        RECT 11.000 104.280 11.170 105.390 ;
        RECT 9.710 104.110 11.170 104.280 ;
        RECT 6.340 102.110 9.070 103.110 ;
        RECT 9.710 102.250 9.980 104.110 ;
        RECT 10.840 103.610 11.170 104.110 ;
        RECT 11.350 103.900 11.600 105.210 ;
        RECT 11.840 104.590 12.090 105.210 ;
        RECT 12.270 104.940 12.440 105.390 ;
        RECT 12.620 105.430 12.950 105.460 ;
        RECT 12.620 105.260 12.650 105.430 ;
        RECT 12.820 105.260 12.950 105.430 ;
        RECT 12.620 105.120 12.950 105.260 ;
        RECT 13.130 105.390 14.870 105.560 ;
        RECT 13.130 104.940 13.300 105.390 ;
        RECT 12.270 104.770 13.300 104.940 ;
        RECT 13.480 104.590 13.650 105.210 ;
        RECT 14.180 104.950 14.510 105.210 ;
        RECT 11.840 104.420 13.650 104.590 ;
        RECT 13.830 104.420 14.050 104.750 ;
        RECT 13.480 104.240 13.650 104.420 ;
        RECT 11.350 103.670 11.880 103.900 ;
        RECT 11.350 102.750 11.620 103.670 ;
      LAYER li1 ;
        RECT 12.300 103.370 12.840 104.240 ;
      LAYER li1 ;
        RECT 13.480 104.070 13.700 104.240 ;
        RECT 10.160 102.120 11.110 102.750 ;
        RECT 11.290 102.250 11.620 102.750 ;
        RECT 11.800 102.120 12.390 103.000 ;
      LAYER li1 ;
        RECT 12.670 102.380 12.840 103.370 ;
        RECT 13.020 102.560 13.350 103.860 ;
      LAYER li1 ;
        RECT 13.530 103.080 13.700 104.070 ;
        RECT 13.880 103.900 14.050 104.420 ;
        RECT 14.230 104.250 14.400 104.950 ;
        RECT 14.700 104.800 14.870 105.390 ;
        RECT 15.050 105.430 16.000 105.460 ;
        RECT 15.050 105.260 15.080 105.430 ;
        RECT 15.250 105.260 15.440 105.430 ;
        RECT 15.610 105.260 15.800 105.430 ;
        RECT 15.970 105.260 16.000 105.430 ;
        RECT 15.050 104.980 16.000 105.260 ;
        RECT 16.180 105.390 17.210 105.560 ;
        RECT 16.180 104.800 16.350 105.390 ;
        RECT 14.700 104.750 16.350 104.800 ;
        RECT 14.580 104.630 16.350 104.750 ;
        RECT 14.580 104.430 14.910 104.630 ;
        RECT 16.530 104.450 16.860 105.210 ;
        RECT 17.040 105.030 17.210 105.390 ;
        RECT 17.390 105.430 18.340 105.510 ;
        RECT 17.390 105.260 17.420 105.430 ;
        RECT 17.590 105.260 17.780 105.430 ;
        RECT 17.950 105.260 18.140 105.430 ;
        RECT 18.310 105.260 18.340 105.430 ;
        RECT 17.390 105.210 18.340 105.260 ;
        RECT 17.040 104.860 18.850 105.030 ;
        RECT 15.090 104.280 16.860 104.450 ;
        RECT 15.090 104.250 15.260 104.280 ;
        RECT 14.230 104.080 15.260 104.250 ;
        RECT 18.170 104.100 18.500 104.680 ;
        RECT 13.880 103.670 14.910 103.900 ;
        RECT 14.580 103.180 14.910 103.670 ;
        RECT 15.090 103.400 15.260 104.080 ;
        RECT 15.440 103.930 18.500 104.100 ;
        RECT 15.440 103.580 15.770 103.930 ;
      LAYER li1 ;
        RECT 16.210 103.580 18.060 103.750 ;
      LAYER li1 ;
        RECT 15.090 103.230 17.710 103.400 ;
        RECT 13.530 102.580 13.800 103.080 ;
        RECT 15.090 103.000 15.260 103.230 ;
      LAYER li1 ;
        RECT 17.890 103.050 18.060 103.580 ;
      LAYER li1 ;
        RECT 14.250 102.830 15.260 103.000 ;
      LAYER li1 ;
        RECT 15.440 102.880 18.060 103.050 ;
      LAYER li1 ;
        RECT 14.250 102.580 14.580 102.830 ;
      LAYER li1 ;
        RECT 15.440 102.380 15.610 102.880 ;
        RECT 12.670 102.210 15.610 102.380 ;
      LAYER li1 ;
        RECT 16.760 102.120 17.710 102.700 ;
      LAYER li1 ;
        RECT 17.890 102.190 18.060 102.880 ;
      LAYER li1 ;
        RECT 18.240 103.080 18.500 103.930 ;
        RECT 18.680 103.510 18.850 104.860 ;
        RECT 19.030 104.600 19.280 105.510 ;
        RECT 20.090 105.430 21.040 105.460 ;
        RECT 21.870 105.430 22.770 105.460 ;
        RECT 20.090 105.260 20.120 105.430 ;
        RECT 20.290 105.260 20.480 105.430 ;
        RECT 20.650 105.260 20.840 105.430 ;
        RECT 21.010 105.260 21.040 105.430 ;
        RECT 22.040 105.260 22.230 105.430 ;
        RECT 22.400 105.260 22.590 105.430 ;
        RECT 22.760 105.260 22.770 105.430 ;
        RECT 19.030 104.430 19.910 104.600 ;
        RECT 20.090 104.430 21.040 105.260 ;
        RECT 21.440 104.460 21.690 104.930 ;
        RECT 21.870 104.640 22.770 105.260 ;
        RECT 23.380 105.430 24.320 105.490 ;
        RECT 23.380 105.260 23.400 105.430 ;
        RECT 23.570 105.260 23.760 105.430 ;
        RECT 23.930 105.260 24.120 105.430 ;
        RECT 24.290 105.260 24.320 105.430 ;
        RECT 19.230 103.690 19.560 104.190 ;
        RECT 19.740 104.110 19.910 104.430 ;
        RECT 21.440 104.290 22.450 104.460 ;
        RECT 19.740 103.940 22.100 104.110 ;
        RECT 18.680 103.340 19.850 103.510 ;
        RECT 18.240 102.370 18.570 103.080 ;
        RECT 19.030 102.540 19.360 103.080 ;
        RECT 19.570 102.840 19.850 103.340 ;
        RECT 20.030 102.540 20.200 103.940 ;
        RECT 22.280 103.760 22.450 104.290 ;
        RECT 20.410 103.590 22.450 103.760 ;
        RECT 20.410 103.200 20.740 103.590 ;
      LAYER li1 ;
        RECT 21.060 103.130 21.390 103.410 ;
        RECT 21.060 103.020 21.440 103.130 ;
      LAYER li1 ;
        RECT 19.030 102.370 20.200 102.540 ;
      LAYER li1 ;
        RECT 20.380 102.960 21.440 103.020 ;
        RECT 20.380 102.850 21.390 102.960 ;
        RECT 20.380 102.190 20.550 102.850 ;
      LAYER li1 ;
        RECT 22.220 102.750 22.450 103.590 ;
        RECT 22.950 103.760 23.200 104.760 ;
        RECT 23.380 103.950 24.320 105.260 ;
        RECT 22.950 103.430 24.320 103.760 ;
        RECT 22.950 103.250 23.160 103.430 ;
        RECT 22.830 102.750 23.160 103.250 ;
      LAYER li1 ;
        RECT 17.890 102.020 20.550 102.190 ;
      LAYER li1 ;
        RECT 20.730 102.120 21.680 102.670 ;
        RECT 22.220 102.250 22.550 102.750 ;
        RECT 23.340 102.120 24.290 103.250 ;
      LAYER li1 ;
        RECT 24.500 102.420 24.840 105.490 ;
      LAYER li1 ;
        RECT 25.210 105.480 26.660 105.510 ;
        RECT 25.210 105.310 25.460 105.480 ;
        RECT 25.630 105.310 25.820 105.480 ;
        RECT 25.990 105.310 26.260 105.480 ;
        RECT 26.430 105.310 26.660 105.480 ;
        RECT 25.210 104.440 26.660 105.310 ;
        RECT 26.970 105.430 27.560 105.510 ;
        RECT 26.970 105.260 27.000 105.430 ;
        RECT 27.170 105.260 27.360 105.430 ;
        RECT 27.530 105.260 27.560 105.430 ;
        RECT 25.440 103.000 25.770 103.780 ;
        RECT 25.980 103.450 26.310 104.440 ;
        RECT 26.970 103.930 27.560 105.260 ;
      LAYER li1 ;
        RECT 27.840 103.930 28.230 105.510 ;
      LAYER li1 ;
        RECT 28.570 105.480 30.020 105.510 ;
        RECT 28.570 105.310 28.820 105.480 ;
        RECT 28.990 105.310 29.180 105.480 ;
        RECT 29.350 105.310 29.620 105.480 ;
        RECT 29.790 105.310 30.020 105.480 ;
        RECT 28.570 104.440 30.020 105.310 ;
      LAYER li1 ;
        RECT 27.010 103.300 27.720 103.690 ;
      LAYER li1 ;
        RECT 25.440 102.600 26.740 103.000 ;
        RECT 25.130 102.120 26.740 102.600 ;
        RECT 26.970 102.120 27.560 103.080 ;
      LAYER li1 ;
        RECT 27.900 102.250 28.230 103.930 ;
      LAYER li1 ;
        RECT 28.800 103.000 29.130 103.780 ;
        RECT 29.340 103.450 29.670 104.440 ;
        RECT 28.800 102.600 30.100 103.000 ;
        RECT 28.490 102.120 30.100 102.600 ;
      LAYER li1 ;
        RECT 31.310 102.250 31.580 105.510 ;
      LAYER li1 ;
        RECT 31.760 105.430 32.660 105.510 ;
        RECT 31.760 105.260 31.770 105.430 ;
        RECT 31.940 105.260 32.130 105.430 ;
        RECT 32.300 105.260 32.490 105.430 ;
        RECT 32.840 105.390 34.730 105.560 ;
        RECT 31.760 103.930 32.660 105.260 ;
        RECT 32.840 103.930 33.010 105.390 ;
      LAYER li1 ;
        RECT 33.190 103.530 33.520 105.010 ;
      LAYER li1 ;
        RECT 31.790 103.350 32.120 103.510 ;
        RECT 33.700 103.350 34.030 105.210 ;
        RECT 34.480 103.850 34.730 105.390 ;
        RECT 34.910 105.430 35.860 105.510 ;
        RECT 34.910 105.260 34.940 105.430 ;
        RECT 35.110 105.260 35.300 105.430 ;
        RECT 35.470 105.260 35.660 105.430 ;
        RECT 35.830 105.260 35.860 105.430 ;
        RECT 34.910 104.030 35.860 105.260 ;
        RECT 36.040 103.850 36.370 105.490 ;
        RECT 36.980 105.480 39.720 105.500 ;
        RECT 36.980 105.310 37.190 105.480 ;
        RECT 37.360 105.310 37.630 105.480 ;
        RECT 37.800 105.310 38.040 105.480 ;
        RECT 38.210 105.310 38.470 105.480 ;
        RECT 38.640 105.310 38.910 105.480 ;
        RECT 39.080 105.310 39.320 105.480 ;
        RECT 39.490 105.310 39.720 105.480 ;
        RECT 36.980 104.430 39.720 105.310 ;
        RECT 40.890 105.430 41.840 105.510 ;
        RECT 40.890 105.260 40.920 105.430 ;
        RECT 41.090 105.260 41.280 105.430 ;
        RECT 41.450 105.260 41.640 105.430 ;
        RECT 41.810 105.260 41.840 105.430 ;
        RECT 34.480 103.680 36.370 103.850 ;
        RECT 31.790 103.180 34.060 103.350 ;
      LAYER li1 ;
        RECT 34.230 103.330 34.410 103.500 ;
      LAYER li1 ;
        RECT 31.750 102.120 33.460 103.000 ;
        RECT 33.890 102.380 34.060 103.180 ;
      LAYER li1 ;
        RECT 34.240 102.560 34.410 103.330 ;
        RECT 36.030 103.260 36.360 103.500 ;
      LAYER li1 ;
        RECT 37.220 103.110 37.550 103.780 ;
        RECT 37.950 103.450 38.280 104.430 ;
        RECT 38.500 103.110 38.830 103.780 ;
        RECT 39.230 103.450 39.560 104.430 ;
        RECT 40.890 103.930 41.840 105.260 ;
      LAYER li1 ;
        RECT 42.020 103.830 42.270 105.510 ;
      LAYER li1 ;
        RECT 42.450 105.430 43.400 105.510 ;
        RECT 42.450 105.260 42.480 105.430 ;
        RECT 42.650 105.260 42.840 105.430 ;
        RECT 43.010 105.260 43.200 105.430 ;
        RECT 43.370 105.260 43.400 105.430 ;
        RECT 42.450 104.010 43.400 105.260 ;
      LAYER li1 ;
        RECT 43.580 103.830 43.910 105.510 ;
      LAYER li1 ;
        RECT 44.090 105.430 45.040 105.510 ;
        RECT 44.090 105.260 44.120 105.430 ;
        RECT 44.290 105.260 44.480 105.430 ;
        RECT 44.650 105.260 44.840 105.430 ;
        RECT 45.010 105.260 45.040 105.430 ;
        RECT 44.090 104.050 45.040 105.260 ;
      LAYER li1 ;
        RECT 42.020 103.660 43.910 103.830 ;
        RECT 42.020 103.530 42.190 103.660 ;
        RECT 44.690 103.530 45.020 103.870 ;
        RECT 40.930 103.300 42.190 103.530 ;
      LAYER li1 ;
        RECT 42.370 103.350 44.400 103.480 ;
        RECT 45.220 103.350 45.470 105.510 ;
        RECT 45.850 105.480 47.300 105.510 ;
        RECT 45.850 105.310 46.100 105.480 ;
        RECT 46.270 105.310 46.460 105.480 ;
        RECT 46.630 105.310 46.900 105.480 ;
        RECT 47.070 105.310 47.300 105.480 ;
        RECT 45.850 104.440 47.300 105.310 ;
        RECT 47.610 105.430 48.560 105.510 ;
        RECT 47.610 105.260 47.640 105.430 ;
        RECT 47.810 105.260 48.000 105.430 ;
        RECT 48.170 105.260 48.360 105.430 ;
        RECT 48.530 105.260 48.560 105.430 ;
        RECT 42.370 103.310 45.470 103.350 ;
      LAYER li1 ;
        RECT 42.020 103.130 42.190 103.300 ;
      LAYER li1 ;
        RECT 44.230 103.180 45.470 103.310 ;
        RECT 34.590 102.380 34.840 103.080 ;
        RECT 33.890 102.210 34.840 102.380 ;
        RECT 35.020 102.120 36.330 103.080 ;
        RECT 37.060 102.110 39.790 103.110 ;
        RECT 40.890 102.120 41.840 103.080 ;
      LAYER li1 ;
        RECT 42.020 102.960 43.830 103.130 ;
        RECT 42.020 102.250 42.270 102.960 ;
      LAYER li1 ;
        RECT 42.450 102.120 43.400 102.780 ;
      LAYER li1 ;
        RECT 43.580 102.250 43.830 102.960 ;
      LAYER li1 ;
        RECT 44.010 102.120 44.960 103.000 ;
        RECT 45.140 102.250 45.470 103.180 ;
        RECT 46.080 103.000 46.410 103.780 ;
        RECT 46.620 103.450 46.950 104.440 ;
        RECT 47.610 103.930 48.560 105.260 ;
      LAYER li1 ;
        RECT 48.740 103.830 48.990 105.510 ;
      LAYER li1 ;
        RECT 49.170 105.430 50.120 105.510 ;
        RECT 49.170 105.260 49.200 105.430 ;
        RECT 49.370 105.260 49.560 105.430 ;
        RECT 49.730 105.260 49.920 105.430 ;
        RECT 50.090 105.260 50.120 105.430 ;
        RECT 49.170 104.010 50.120 105.260 ;
      LAYER li1 ;
        RECT 50.300 103.830 50.630 105.510 ;
      LAYER li1 ;
        RECT 50.810 105.430 51.760 105.510 ;
        RECT 50.810 105.260 50.840 105.430 ;
        RECT 51.010 105.260 51.200 105.430 ;
        RECT 51.370 105.260 51.560 105.430 ;
        RECT 51.730 105.260 51.760 105.430 ;
        RECT 50.810 104.050 51.760 105.260 ;
      LAYER li1 ;
        RECT 48.740 103.660 50.630 103.830 ;
        RECT 48.740 103.530 48.910 103.660 ;
        RECT 51.410 103.530 51.740 103.870 ;
        RECT 47.650 103.300 48.910 103.530 ;
      LAYER li1 ;
        RECT 49.090 103.350 51.120 103.480 ;
        RECT 51.940 103.350 52.190 105.510 ;
        RECT 52.570 105.480 54.020 105.510 ;
        RECT 52.570 105.310 52.820 105.480 ;
        RECT 52.990 105.310 53.180 105.480 ;
        RECT 53.350 105.310 53.620 105.480 ;
        RECT 53.790 105.310 54.020 105.480 ;
        RECT 52.570 104.440 54.020 105.310 ;
        RECT 54.330 105.430 55.280 105.510 ;
        RECT 54.330 105.260 54.360 105.430 ;
        RECT 54.530 105.260 54.720 105.430 ;
        RECT 54.890 105.260 55.080 105.430 ;
        RECT 55.250 105.260 55.280 105.430 ;
        RECT 49.090 103.310 52.190 103.350 ;
      LAYER li1 ;
        RECT 48.740 103.130 48.910 103.300 ;
      LAYER li1 ;
        RECT 50.950 103.180 52.190 103.310 ;
        RECT 46.080 102.600 47.380 103.000 ;
        RECT 45.770 102.120 47.380 102.600 ;
        RECT 47.610 102.120 48.560 103.080 ;
      LAYER li1 ;
        RECT 48.740 102.960 50.550 103.130 ;
        RECT 48.740 102.250 48.990 102.960 ;
      LAYER li1 ;
        RECT 49.170 102.120 50.120 102.780 ;
      LAYER li1 ;
        RECT 50.300 102.250 50.550 102.960 ;
      LAYER li1 ;
        RECT 50.730 102.120 51.680 103.000 ;
        RECT 51.860 102.250 52.190 103.180 ;
        RECT 52.800 103.000 53.130 103.780 ;
        RECT 53.340 103.450 53.670 104.440 ;
        RECT 54.330 103.930 55.280 105.260 ;
      LAYER li1 ;
        RECT 55.460 103.830 55.710 105.510 ;
      LAYER li1 ;
        RECT 55.890 105.430 56.840 105.510 ;
        RECT 55.890 105.260 55.920 105.430 ;
        RECT 56.090 105.260 56.280 105.430 ;
        RECT 56.450 105.260 56.640 105.430 ;
        RECT 56.810 105.260 56.840 105.430 ;
        RECT 55.890 104.010 56.840 105.260 ;
      LAYER li1 ;
        RECT 57.020 103.830 57.350 105.510 ;
      LAYER li1 ;
        RECT 57.530 105.430 58.480 105.510 ;
        RECT 57.530 105.260 57.560 105.430 ;
        RECT 57.730 105.260 57.920 105.430 ;
        RECT 58.090 105.260 58.280 105.430 ;
        RECT 58.450 105.260 58.480 105.430 ;
        RECT 57.530 104.050 58.480 105.260 ;
      LAYER li1 ;
        RECT 55.460 103.660 57.350 103.830 ;
        RECT 55.460 103.530 55.630 103.660 ;
        RECT 58.130 103.530 58.460 103.870 ;
        RECT 54.370 103.300 55.630 103.530 ;
      LAYER li1 ;
        RECT 55.810 103.350 57.840 103.480 ;
        RECT 58.660 103.350 58.910 105.510 ;
        RECT 59.290 105.480 60.740 105.510 ;
        RECT 59.290 105.310 59.540 105.480 ;
        RECT 59.710 105.310 59.900 105.480 ;
        RECT 60.070 105.310 60.340 105.480 ;
        RECT 60.510 105.310 60.740 105.480 ;
        RECT 59.290 104.440 60.740 105.310 ;
        RECT 61.530 105.430 62.120 105.510 ;
        RECT 61.530 105.260 61.560 105.430 ;
        RECT 61.730 105.260 61.920 105.430 ;
        RECT 62.090 105.260 62.120 105.430 ;
        RECT 55.810 103.310 58.910 103.350 ;
      LAYER li1 ;
        RECT 55.460 103.130 55.630 103.300 ;
      LAYER li1 ;
        RECT 57.670 103.180 58.910 103.310 ;
        RECT 52.800 102.600 54.100 103.000 ;
        RECT 52.490 102.120 54.100 102.600 ;
        RECT 54.330 102.120 55.280 103.080 ;
      LAYER li1 ;
        RECT 55.460 102.960 57.270 103.130 ;
        RECT 55.460 102.250 55.710 102.960 ;
      LAYER li1 ;
        RECT 55.890 102.120 56.840 102.780 ;
      LAYER li1 ;
        RECT 57.020 102.250 57.270 102.960 ;
      LAYER li1 ;
        RECT 57.450 102.120 58.400 103.000 ;
        RECT 58.580 102.250 58.910 103.180 ;
        RECT 59.520 103.000 59.850 103.780 ;
        RECT 60.060 103.450 60.390 104.440 ;
        RECT 61.530 103.930 62.120 105.260 ;
      LAYER li1 ;
        RECT 62.400 103.930 62.790 105.510 ;
      LAYER li1 ;
        RECT 63.130 105.480 64.580 105.510 ;
        RECT 63.130 105.310 63.380 105.480 ;
        RECT 63.550 105.310 63.740 105.480 ;
        RECT 63.910 105.310 64.180 105.480 ;
        RECT 64.350 105.310 64.580 105.480 ;
        RECT 63.130 104.440 64.580 105.310 ;
        RECT 65.430 105.430 66.020 105.460 ;
        RECT 65.430 105.260 65.460 105.430 ;
        RECT 65.630 105.260 65.820 105.430 ;
        RECT 65.990 105.260 66.020 105.430 ;
        RECT 59.520 102.600 60.820 103.000 ;
        RECT 59.210 102.120 60.820 102.600 ;
        RECT 61.530 102.120 62.120 103.080 ;
      LAYER li1 ;
        RECT 62.460 102.250 62.790 103.930 ;
      LAYER li1 ;
        RECT 63.360 103.000 63.690 103.780 ;
        RECT 63.900 103.450 64.230 104.440 ;
        RECT 64.910 104.280 65.240 105.210 ;
        RECT 65.430 104.480 66.020 105.260 ;
        RECT 66.200 105.390 67.640 105.560 ;
        RECT 66.200 104.280 66.370 105.390 ;
        RECT 64.910 104.110 66.370 104.280 ;
        RECT 63.360 102.600 64.660 103.000 ;
        RECT 63.050 102.120 64.660 102.600 ;
        RECT 64.910 102.250 65.180 104.110 ;
      LAYER li1 ;
        RECT 65.360 102.930 65.690 103.900 ;
      LAYER li1 ;
        RECT 66.040 103.610 66.370 104.110 ;
        RECT 66.550 103.900 66.800 105.210 ;
        RECT 67.040 104.590 67.290 105.210 ;
        RECT 67.470 104.940 67.640 105.390 ;
        RECT 67.820 105.430 68.150 105.460 ;
        RECT 67.820 105.260 67.850 105.430 ;
        RECT 68.020 105.260 68.150 105.430 ;
        RECT 67.820 105.120 68.150 105.260 ;
        RECT 68.330 105.390 70.070 105.560 ;
        RECT 68.330 104.940 68.500 105.390 ;
        RECT 67.470 104.770 68.500 104.940 ;
        RECT 68.680 104.590 68.850 105.210 ;
        RECT 69.380 104.950 69.710 105.210 ;
        RECT 67.040 104.420 68.850 104.590 ;
        RECT 69.030 104.420 69.250 104.750 ;
        RECT 68.680 104.240 68.850 104.420 ;
        RECT 66.550 103.670 67.080 103.900 ;
        RECT 66.550 102.750 66.820 103.670 ;
      LAYER li1 ;
        RECT 67.500 103.370 68.040 104.240 ;
      LAYER li1 ;
        RECT 68.680 104.070 68.900 104.240 ;
        RECT 65.360 102.120 66.310 102.750 ;
        RECT 66.490 102.250 66.820 102.750 ;
        RECT 67.000 102.120 67.590 103.000 ;
      LAYER li1 ;
        RECT 67.870 102.380 68.040 103.370 ;
        RECT 68.220 102.560 68.550 103.860 ;
      LAYER li1 ;
        RECT 68.730 103.080 68.900 104.070 ;
        RECT 69.080 103.900 69.250 104.420 ;
        RECT 69.430 104.250 69.600 104.950 ;
        RECT 69.900 104.800 70.070 105.390 ;
        RECT 70.250 105.430 71.200 105.460 ;
        RECT 70.250 105.260 70.280 105.430 ;
        RECT 70.450 105.260 70.640 105.430 ;
        RECT 70.810 105.260 71.000 105.430 ;
        RECT 71.170 105.260 71.200 105.430 ;
        RECT 70.250 104.980 71.200 105.260 ;
        RECT 71.380 105.390 72.410 105.560 ;
        RECT 71.380 104.800 71.550 105.390 ;
        RECT 69.900 104.750 71.550 104.800 ;
        RECT 69.780 104.630 71.550 104.750 ;
        RECT 69.780 104.430 70.110 104.630 ;
        RECT 71.730 104.450 72.060 105.210 ;
        RECT 72.240 105.030 72.410 105.390 ;
        RECT 72.590 105.430 73.540 105.510 ;
        RECT 72.590 105.260 72.620 105.430 ;
        RECT 72.790 105.260 72.980 105.430 ;
        RECT 73.150 105.260 73.340 105.430 ;
        RECT 73.510 105.260 73.540 105.430 ;
        RECT 72.590 105.210 73.540 105.260 ;
        RECT 72.240 104.860 74.050 105.030 ;
        RECT 70.290 104.280 72.060 104.450 ;
        RECT 70.290 104.250 70.460 104.280 ;
        RECT 69.430 104.080 70.460 104.250 ;
        RECT 73.370 104.100 73.700 104.680 ;
        RECT 69.080 103.670 70.110 103.900 ;
        RECT 69.780 103.180 70.110 103.670 ;
        RECT 70.290 103.400 70.460 104.080 ;
        RECT 70.640 103.930 73.700 104.100 ;
        RECT 70.640 103.580 70.970 103.930 ;
      LAYER li1 ;
        RECT 71.410 103.580 73.260 103.750 ;
      LAYER li1 ;
        RECT 70.290 103.230 72.910 103.400 ;
        RECT 68.730 102.580 69.000 103.080 ;
        RECT 70.290 103.000 70.460 103.230 ;
      LAYER li1 ;
        RECT 73.090 103.050 73.260 103.580 ;
      LAYER li1 ;
        RECT 69.450 102.830 70.460 103.000 ;
      LAYER li1 ;
        RECT 70.640 102.880 73.260 103.050 ;
      LAYER li1 ;
        RECT 69.450 102.580 69.780 102.830 ;
      LAYER li1 ;
        RECT 70.640 102.380 70.810 102.880 ;
        RECT 67.870 102.210 70.810 102.380 ;
      LAYER li1 ;
        RECT 71.960 102.120 72.910 102.700 ;
      LAYER li1 ;
        RECT 73.090 102.190 73.260 102.880 ;
      LAYER li1 ;
        RECT 73.440 103.080 73.700 103.930 ;
        RECT 73.880 103.510 74.050 104.860 ;
        RECT 74.230 104.600 74.480 105.510 ;
        RECT 75.290 105.430 76.240 105.460 ;
        RECT 77.070 105.430 77.970 105.460 ;
        RECT 75.290 105.260 75.320 105.430 ;
        RECT 75.490 105.260 75.680 105.430 ;
        RECT 75.850 105.260 76.040 105.430 ;
        RECT 76.210 105.260 76.240 105.430 ;
        RECT 77.240 105.260 77.430 105.430 ;
        RECT 77.600 105.260 77.790 105.430 ;
        RECT 77.960 105.260 77.970 105.430 ;
        RECT 74.230 104.430 75.110 104.600 ;
        RECT 75.290 104.430 76.240 105.260 ;
        RECT 76.640 104.460 76.890 104.930 ;
        RECT 77.070 104.640 77.970 105.260 ;
        RECT 78.580 105.430 79.520 105.490 ;
        RECT 78.580 105.260 78.600 105.430 ;
        RECT 78.770 105.260 78.960 105.430 ;
        RECT 79.130 105.260 79.320 105.430 ;
        RECT 79.490 105.260 79.520 105.430 ;
        RECT 74.430 103.690 74.760 104.190 ;
        RECT 74.940 104.110 75.110 104.430 ;
        RECT 76.640 104.290 77.650 104.460 ;
        RECT 74.940 103.940 77.300 104.110 ;
        RECT 73.880 103.340 75.050 103.510 ;
        RECT 73.440 102.370 73.770 103.080 ;
        RECT 74.230 102.540 74.560 103.080 ;
        RECT 74.770 102.840 75.050 103.340 ;
        RECT 75.230 102.540 75.400 103.940 ;
        RECT 77.480 103.760 77.650 104.290 ;
        RECT 75.610 103.590 77.650 103.760 ;
        RECT 75.610 103.200 75.940 103.590 ;
      LAYER li1 ;
        RECT 76.260 103.130 76.590 103.410 ;
        RECT 76.260 103.020 76.640 103.130 ;
      LAYER li1 ;
        RECT 74.230 102.370 75.400 102.540 ;
      LAYER li1 ;
        RECT 75.580 102.960 76.640 103.020 ;
        RECT 75.580 102.850 76.590 102.960 ;
        RECT 75.580 102.190 75.750 102.850 ;
      LAYER li1 ;
        RECT 77.420 102.750 77.650 103.590 ;
        RECT 78.150 103.760 78.400 104.760 ;
        RECT 78.580 103.950 79.520 105.260 ;
        RECT 78.150 103.430 79.520 103.760 ;
        RECT 78.150 103.250 78.360 103.430 ;
        RECT 78.030 102.750 78.360 103.250 ;
      LAYER li1 ;
        RECT 73.090 102.020 75.750 102.190 ;
      LAYER li1 ;
        RECT 75.930 102.120 76.880 102.670 ;
        RECT 77.420 102.250 77.750 102.750 ;
        RECT 78.540 102.120 79.490 103.250 ;
      LAYER li1 ;
        RECT 79.700 102.420 80.040 105.490 ;
      LAYER li1 ;
        RECT 80.410 105.480 81.860 105.510 ;
        RECT 80.410 105.310 80.660 105.480 ;
        RECT 80.830 105.310 81.020 105.480 ;
        RECT 81.190 105.310 81.460 105.480 ;
        RECT 81.630 105.310 81.860 105.480 ;
        RECT 80.410 104.440 81.860 105.310 ;
        RECT 82.170 105.430 83.120 105.510 ;
        RECT 82.170 105.260 82.200 105.430 ;
        RECT 82.370 105.260 82.560 105.430 ;
        RECT 82.730 105.260 82.920 105.430 ;
        RECT 83.090 105.260 83.120 105.430 ;
        RECT 80.640 103.000 80.970 103.780 ;
        RECT 81.180 103.450 81.510 104.440 ;
        RECT 82.170 103.930 83.120 105.260 ;
      LAYER li1 ;
        RECT 83.300 103.830 83.550 105.510 ;
      LAYER li1 ;
        RECT 83.730 105.430 84.680 105.510 ;
        RECT 83.730 105.260 83.760 105.430 ;
        RECT 83.930 105.260 84.120 105.430 ;
        RECT 84.290 105.260 84.480 105.430 ;
        RECT 84.650 105.260 84.680 105.430 ;
        RECT 83.730 104.010 84.680 105.260 ;
      LAYER li1 ;
        RECT 84.860 103.830 85.190 105.510 ;
      LAYER li1 ;
        RECT 85.370 105.430 86.320 105.510 ;
        RECT 85.370 105.260 85.400 105.430 ;
        RECT 85.570 105.260 85.760 105.430 ;
        RECT 85.930 105.260 86.120 105.430 ;
        RECT 86.290 105.260 86.320 105.430 ;
        RECT 85.370 104.050 86.320 105.260 ;
      LAYER li1 ;
        RECT 83.300 103.660 85.190 103.830 ;
        RECT 83.300 103.530 83.470 103.660 ;
        RECT 85.970 103.530 86.300 103.870 ;
        RECT 82.210 103.300 83.470 103.530 ;
      LAYER li1 ;
        RECT 83.650 103.350 85.680 103.480 ;
        RECT 86.500 103.350 86.750 105.510 ;
        RECT 87.130 105.480 88.580 105.510 ;
        RECT 87.130 105.310 87.380 105.480 ;
        RECT 87.550 105.310 87.740 105.480 ;
        RECT 87.910 105.310 88.180 105.480 ;
        RECT 88.350 105.310 88.580 105.480 ;
        RECT 87.130 104.440 88.580 105.310 ;
        RECT 88.890 105.430 89.840 105.510 ;
        RECT 88.890 105.260 88.920 105.430 ;
        RECT 89.090 105.260 89.280 105.430 ;
        RECT 89.450 105.260 89.640 105.430 ;
        RECT 89.810 105.260 89.840 105.430 ;
        RECT 83.650 103.310 86.750 103.350 ;
      LAYER li1 ;
        RECT 83.300 103.130 83.470 103.300 ;
      LAYER li1 ;
        RECT 85.510 103.180 86.750 103.310 ;
        RECT 80.640 102.600 81.940 103.000 ;
        RECT 80.330 102.120 81.940 102.600 ;
        RECT 82.170 102.120 83.120 103.080 ;
      LAYER li1 ;
        RECT 83.300 102.960 85.110 103.130 ;
        RECT 83.300 102.250 83.550 102.960 ;
      LAYER li1 ;
        RECT 83.730 102.120 84.680 102.780 ;
      LAYER li1 ;
        RECT 84.860 102.250 85.110 102.960 ;
      LAYER li1 ;
        RECT 85.290 102.120 86.240 103.000 ;
        RECT 86.420 102.250 86.750 103.180 ;
        RECT 87.360 103.000 87.690 103.780 ;
        RECT 87.900 103.450 88.230 104.440 ;
        RECT 88.890 103.930 89.840 105.260 ;
      LAYER li1 ;
        RECT 90.020 103.830 90.270 105.510 ;
      LAYER li1 ;
        RECT 90.450 105.430 91.400 105.510 ;
        RECT 90.450 105.260 90.480 105.430 ;
        RECT 90.650 105.260 90.840 105.430 ;
        RECT 91.010 105.260 91.200 105.430 ;
        RECT 91.370 105.260 91.400 105.430 ;
        RECT 90.450 104.010 91.400 105.260 ;
      LAYER li1 ;
        RECT 91.580 103.830 91.910 105.510 ;
      LAYER li1 ;
        RECT 92.090 105.430 93.040 105.510 ;
        RECT 92.090 105.260 92.120 105.430 ;
        RECT 92.290 105.260 92.480 105.430 ;
        RECT 92.650 105.260 92.840 105.430 ;
        RECT 93.010 105.260 93.040 105.430 ;
        RECT 92.090 104.050 93.040 105.260 ;
      LAYER li1 ;
        RECT 90.020 103.660 91.910 103.830 ;
        RECT 90.020 103.530 90.190 103.660 ;
        RECT 92.690 103.530 93.020 103.870 ;
        RECT 88.930 103.300 90.190 103.530 ;
      LAYER li1 ;
        RECT 90.370 103.350 92.400 103.480 ;
        RECT 93.220 103.350 93.470 105.510 ;
        RECT 94.100 105.480 96.840 105.500 ;
        RECT 94.100 105.310 94.310 105.480 ;
        RECT 94.480 105.310 94.750 105.480 ;
        RECT 94.920 105.310 95.160 105.480 ;
        RECT 95.330 105.310 95.590 105.480 ;
        RECT 95.760 105.310 96.030 105.480 ;
        RECT 96.200 105.310 96.440 105.480 ;
        RECT 96.610 105.310 96.840 105.480 ;
        RECT 94.100 104.430 96.840 105.310 ;
        RECT 90.370 103.310 93.470 103.350 ;
      LAYER li1 ;
        RECT 90.020 103.130 90.190 103.300 ;
      LAYER li1 ;
        RECT 92.230 103.180 93.470 103.310 ;
        RECT 87.360 102.600 88.660 103.000 ;
        RECT 87.050 102.120 88.660 102.600 ;
        RECT 88.890 102.120 89.840 103.080 ;
      LAYER li1 ;
        RECT 90.020 102.960 91.830 103.130 ;
        RECT 90.020 102.250 90.270 102.960 ;
      LAYER li1 ;
        RECT 90.450 102.120 91.400 102.780 ;
      LAYER li1 ;
        RECT 91.580 102.250 91.830 102.960 ;
      LAYER li1 ;
        RECT 92.010 102.120 92.960 103.000 ;
        RECT 93.140 102.250 93.470 103.180 ;
        RECT 94.340 103.110 94.670 103.780 ;
        RECT 95.070 103.450 95.400 104.430 ;
        RECT 95.620 103.110 95.950 103.780 ;
        RECT 96.350 103.450 96.680 104.430 ;
        RECT 94.180 102.110 96.910 103.110 ;
      LAYER li1 ;
        RECT 98.530 102.250 98.780 105.510 ;
      LAYER li1 ;
        RECT 98.960 105.430 101.650 105.510 ;
        RECT 99.130 105.260 99.320 105.430 ;
        RECT 99.490 105.260 99.680 105.430 ;
        RECT 99.850 105.260 100.040 105.430 ;
        RECT 100.210 105.260 100.400 105.430 ;
        RECT 100.570 105.260 100.760 105.430 ;
        RECT 100.930 105.260 101.120 105.430 ;
        RECT 101.290 105.260 101.480 105.430 ;
        RECT 98.960 104.400 101.650 105.260 ;
        RECT 101.830 104.220 102.080 105.510 ;
        RECT 98.990 104.050 102.080 104.220 ;
        RECT 98.990 103.350 99.320 104.050 ;
        RECT 101.830 103.930 102.080 104.050 ;
        RECT 102.260 105.430 103.570 105.490 ;
        RECT 102.260 105.260 102.290 105.430 ;
        RECT 102.460 105.260 102.650 105.430 ;
        RECT 102.820 105.260 103.010 105.430 ;
        RECT 103.180 105.260 103.370 105.430 ;
        RECT 103.540 105.260 103.570 105.430 ;
        RECT 102.260 103.950 103.570 105.260 ;
        RECT 103.930 105.480 105.380 105.510 ;
        RECT 103.930 105.310 104.180 105.480 ;
        RECT 104.350 105.310 104.540 105.480 ;
        RECT 104.710 105.310 104.980 105.480 ;
        RECT 105.150 105.310 105.380 105.480 ;
        RECT 103.930 104.440 105.380 105.310 ;
        RECT 105.690 105.430 106.640 105.510 ;
        RECT 105.690 105.260 105.720 105.430 ;
        RECT 105.890 105.260 106.080 105.430 ;
        RECT 106.250 105.260 106.440 105.430 ;
        RECT 106.610 105.260 106.640 105.430 ;
      LAYER li1 ;
        RECT 99.990 103.810 100.160 103.870 ;
        RECT 99.820 103.530 100.550 103.810 ;
      LAYER li1 ;
        RECT 98.990 103.180 100.200 103.350 ;
        RECT 98.960 102.120 99.850 103.000 ;
        RECT 100.030 102.970 100.200 103.180 ;
      LAYER li1 ;
        RECT 100.380 103.320 100.550 103.530 ;
        RECT 101.360 103.330 101.650 103.870 ;
        RECT 101.890 103.330 102.600 103.660 ;
        RECT 100.380 103.150 101.180 103.320 ;
        RECT 102.950 103.150 103.280 103.770 ;
        RECT 101.010 102.980 103.280 103.150 ;
      LAYER li1 ;
        RECT 104.160 103.000 104.490 103.780 ;
        RECT 104.700 103.450 105.030 104.440 ;
        RECT 105.690 103.930 106.640 105.260 ;
      LAYER li1 ;
        RECT 106.820 103.830 107.070 105.510 ;
      LAYER li1 ;
        RECT 107.250 105.430 108.200 105.510 ;
        RECT 107.250 105.260 107.280 105.430 ;
        RECT 107.450 105.260 107.640 105.430 ;
        RECT 107.810 105.260 108.000 105.430 ;
        RECT 108.170 105.260 108.200 105.430 ;
        RECT 107.250 104.010 108.200 105.260 ;
      LAYER li1 ;
        RECT 108.380 103.830 108.710 105.510 ;
      LAYER li1 ;
        RECT 108.890 105.430 109.840 105.510 ;
        RECT 108.890 105.260 108.920 105.430 ;
        RECT 109.090 105.260 109.280 105.430 ;
        RECT 109.450 105.260 109.640 105.430 ;
        RECT 109.810 105.260 109.840 105.430 ;
        RECT 108.890 104.050 109.840 105.260 ;
      LAYER li1 ;
        RECT 106.820 103.660 108.710 103.830 ;
        RECT 106.820 103.530 106.990 103.660 ;
        RECT 109.490 103.530 109.820 103.870 ;
        RECT 105.730 103.300 106.990 103.530 ;
      LAYER li1 ;
        RECT 107.170 103.350 109.200 103.480 ;
        RECT 110.020 103.350 110.270 105.510 ;
        RECT 110.650 105.480 112.100 105.510 ;
        RECT 110.650 105.310 110.900 105.480 ;
        RECT 111.070 105.310 111.260 105.480 ;
        RECT 111.430 105.310 111.700 105.480 ;
        RECT 111.870 105.310 112.100 105.480 ;
        RECT 110.650 104.440 112.100 105.310 ;
        RECT 112.410 105.430 113.360 105.510 ;
        RECT 112.410 105.260 112.440 105.430 ;
        RECT 112.610 105.260 112.800 105.430 ;
        RECT 112.970 105.260 113.160 105.430 ;
        RECT 113.330 105.260 113.360 105.430 ;
        RECT 107.170 103.310 110.270 103.350 ;
      LAYER li1 ;
        RECT 106.820 103.130 106.990 103.300 ;
      LAYER li1 ;
        RECT 109.030 103.180 110.270 103.310 ;
        RECT 100.030 102.800 100.830 102.970 ;
      LAYER li1 ;
        RECT 101.440 102.960 102.110 102.980 ;
      LAYER li1 ;
        RECT 100.660 102.630 101.260 102.800 ;
        RECT 100.150 102.190 100.480 102.620 ;
        RECT 100.930 102.370 101.260 102.630 ;
        RECT 101.750 102.190 102.080 102.780 ;
        RECT 100.150 102.020 102.080 102.190 ;
        RECT 102.290 102.120 103.590 102.800 ;
        RECT 104.160 102.600 105.460 103.000 ;
        RECT 103.850 102.120 105.460 102.600 ;
        RECT 105.690 102.120 106.640 103.080 ;
      LAYER li1 ;
        RECT 106.820 102.960 108.630 103.130 ;
        RECT 106.820 102.250 107.070 102.960 ;
      LAYER li1 ;
        RECT 107.250 102.120 108.200 102.780 ;
      LAYER li1 ;
        RECT 108.380 102.250 108.630 102.960 ;
      LAYER li1 ;
        RECT 108.810 102.120 109.760 103.000 ;
        RECT 109.940 102.250 110.270 103.180 ;
        RECT 110.880 103.000 111.210 103.780 ;
        RECT 111.420 103.450 111.750 104.440 ;
        RECT 112.410 103.930 113.360 105.260 ;
      LAYER li1 ;
        RECT 113.540 103.830 113.790 105.510 ;
      LAYER li1 ;
        RECT 113.970 105.430 114.920 105.510 ;
        RECT 113.970 105.260 114.000 105.430 ;
        RECT 114.170 105.260 114.360 105.430 ;
        RECT 114.530 105.260 114.720 105.430 ;
        RECT 114.890 105.260 114.920 105.430 ;
        RECT 113.970 104.010 114.920 105.260 ;
      LAYER li1 ;
        RECT 115.100 103.830 115.430 105.510 ;
      LAYER li1 ;
        RECT 115.610 105.430 116.560 105.510 ;
        RECT 115.610 105.260 115.640 105.430 ;
        RECT 115.810 105.260 116.000 105.430 ;
        RECT 116.170 105.260 116.360 105.430 ;
        RECT 116.530 105.260 116.560 105.430 ;
        RECT 115.610 104.050 116.560 105.260 ;
      LAYER li1 ;
        RECT 113.540 103.660 115.430 103.830 ;
        RECT 113.540 103.530 113.710 103.660 ;
        RECT 116.210 103.530 116.540 103.870 ;
        RECT 112.450 103.300 113.710 103.530 ;
      LAYER li1 ;
        RECT 113.890 103.350 115.920 103.480 ;
        RECT 116.740 103.350 116.990 105.510 ;
        RECT 117.620 105.480 120.360 105.500 ;
        RECT 117.620 105.310 117.830 105.480 ;
        RECT 118.000 105.310 118.270 105.480 ;
        RECT 118.440 105.310 118.680 105.480 ;
        RECT 118.850 105.310 119.110 105.480 ;
        RECT 119.280 105.310 119.550 105.480 ;
        RECT 119.720 105.310 119.960 105.480 ;
        RECT 120.130 105.310 120.360 105.480 ;
        RECT 117.620 104.430 120.360 105.310 ;
        RECT 121.530 105.430 122.480 105.510 ;
        RECT 121.530 105.260 121.560 105.430 ;
        RECT 121.730 105.260 121.920 105.430 ;
        RECT 122.090 105.260 122.280 105.430 ;
        RECT 122.450 105.260 122.480 105.430 ;
        RECT 113.890 103.310 116.990 103.350 ;
      LAYER li1 ;
        RECT 113.540 103.130 113.710 103.300 ;
      LAYER li1 ;
        RECT 115.750 103.180 116.990 103.310 ;
        RECT 110.880 102.600 112.180 103.000 ;
        RECT 110.570 102.120 112.180 102.600 ;
        RECT 112.410 102.120 113.360 103.080 ;
      LAYER li1 ;
        RECT 113.540 102.960 115.350 103.130 ;
        RECT 113.540 102.250 113.790 102.960 ;
      LAYER li1 ;
        RECT 113.970 102.120 114.920 102.780 ;
      LAYER li1 ;
        RECT 115.100 102.250 115.350 102.960 ;
      LAYER li1 ;
        RECT 115.530 102.120 116.480 103.000 ;
        RECT 116.660 102.250 116.990 103.180 ;
        RECT 117.860 103.110 118.190 103.780 ;
        RECT 118.590 103.450 118.920 104.430 ;
        RECT 119.140 103.110 119.470 103.780 ;
        RECT 119.870 103.450 120.200 104.430 ;
        RECT 121.530 103.930 122.480 105.260 ;
      LAYER li1 ;
        RECT 122.660 103.830 122.910 105.510 ;
      LAYER li1 ;
        RECT 123.090 105.430 124.040 105.510 ;
        RECT 123.090 105.260 123.120 105.430 ;
        RECT 123.290 105.260 123.480 105.430 ;
        RECT 123.650 105.260 123.840 105.430 ;
        RECT 124.010 105.260 124.040 105.430 ;
        RECT 123.090 104.010 124.040 105.260 ;
      LAYER li1 ;
        RECT 124.220 103.830 124.550 105.510 ;
      LAYER li1 ;
        RECT 124.730 105.430 125.680 105.510 ;
        RECT 124.730 105.260 124.760 105.430 ;
        RECT 124.930 105.260 125.120 105.430 ;
        RECT 125.290 105.260 125.480 105.430 ;
        RECT 125.650 105.260 125.680 105.430 ;
        RECT 124.730 104.050 125.680 105.260 ;
      LAYER li1 ;
        RECT 122.660 103.660 124.550 103.830 ;
        RECT 122.660 103.530 122.830 103.660 ;
        RECT 125.330 103.530 125.660 103.870 ;
        RECT 121.570 103.300 122.830 103.530 ;
      LAYER li1 ;
        RECT 123.010 103.350 125.040 103.480 ;
        RECT 125.860 103.350 126.110 105.510 ;
        RECT 126.740 105.480 129.480 105.500 ;
        RECT 126.740 105.310 126.950 105.480 ;
        RECT 127.120 105.310 127.390 105.480 ;
        RECT 127.560 105.310 127.800 105.480 ;
        RECT 127.970 105.310 128.230 105.480 ;
        RECT 128.400 105.310 128.670 105.480 ;
        RECT 128.840 105.310 129.080 105.480 ;
        RECT 129.250 105.310 129.480 105.480 ;
        RECT 126.740 104.430 129.480 105.310 ;
        RECT 130.580 105.480 133.320 105.500 ;
        RECT 130.580 105.310 130.790 105.480 ;
        RECT 130.960 105.310 131.230 105.480 ;
        RECT 131.400 105.310 131.640 105.480 ;
        RECT 131.810 105.310 132.070 105.480 ;
        RECT 132.240 105.310 132.510 105.480 ;
        RECT 132.680 105.310 132.920 105.480 ;
        RECT 133.090 105.310 133.320 105.480 ;
        RECT 130.580 104.430 133.320 105.310 ;
        RECT 134.970 105.430 135.560 105.510 ;
        RECT 134.970 105.260 135.000 105.430 ;
        RECT 135.170 105.260 135.360 105.430 ;
        RECT 135.530 105.260 135.560 105.430 ;
        RECT 123.010 103.310 126.110 103.350 ;
      LAYER li1 ;
        RECT 122.660 103.130 122.830 103.300 ;
      LAYER li1 ;
        RECT 124.870 103.180 126.110 103.310 ;
        RECT 117.700 102.110 120.430 103.110 ;
        RECT 121.530 102.120 122.480 103.080 ;
      LAYER li1 ;
        RECT 122.660 102.960 124.470 103.130 ;
        RECT 122.660 102.250 122.910 102.960 ;
      LAYER li1 ;
        RECT 123.090 102.120 124.040 102.780 ;
      LAYER li1 ;
        RECT 124.220 102.250 124.470 102.960 ;
      LAYER li1 ;
        RECT 124.650 102.120 125.600 103.000 ;
        RECT 125.780 102.250 126.110 103.180 ;
        RECT 126.980 103.110 127.310 103.780 ;
        RECT 127.710 103.450 128.040 104.430 ;
        RECT 128.260 103.110 128.590 103.780 ;
        RECT 128.990 103.450 129.320 104.430 ;
        RECT 130.820 103.110 131.150 103.780 ;
        RECT 131.550 103.450 131.880 104.430 ;
        RECT 132.100 103.110 132.430 103.780 ;
        RECT 132.830 103.450 133.160 104.430 ;
        RECT 134.970 103.930 135.560 105.260 ;
      LAYER li1 ;
        RECT 135.840 103.930 136.230 105.510 ;
      LAYER li1 ;
        RECT 136.820 105.480 139.560 105.500 ;
        RECT 136.820 105.310 137.030 105.480 ;
        RECT 137.200 105.310 137.470 105.480 ;
        RECT 137.640 105.310 137.880 105.480 ;
        RECT 138.050 105.310 138.310 105.480 ;
        RECT 138.480 105.310 138.750 105.480 ;
        RECT 138.920 105.310 139.160 105.480 ;
        RECT 139.330 105.310 139.560 105.480 ;
        RECT 136.820 104.430 139.560 105.310 ;
        RECT 140.410 105.480 141.860 105.510 ;
        RECT 140.410 105.310 140.660 105.480 ;
        RECT 140.830 105.310 141.020 105.480 ;
        RECT 141.190 105.310 141.460 105.480 ;
        RECT 141.630 105.310 141.860 105.480 ;
        RECT 140.410 104.440 141.860 105.310 ;
        RECT 126.820 102.110 129.550 103.110 ;
        RECT 130.660 102.110 133.390 103.110 ;
        RECT 134.970 102.120 135.560 103.080 ;
      LAYER li1 ;
        RECT 135.900 102.250 136.230 103.930 ;
      LAYER li1 ;
        RECT 137.060 103.110 137.390 103.780 ;
        RECT 137.790 103.450 138.120 104.430 ;
        RECT 138.340 103.110 138.670 103.780 ;
        RECT 139.070 103.450 139.400 104.430 ;
        RECT 136.900 102.110 139.630 103.110 ;
        RECT 140.640 103.000 140.970 103.780 ;
        RECT 141.180 103.450 141.510 104.440 ;
        RECT 140.640 102.600 141.940 103.000 ;
        RECT 140.330 102.120 141.940 102.600 ;
        RECT 5.760 101.660 5.920 101.840 ;
        RECT 6.090 101.660 6.400 101.840 ;
        RECT 6.570 101.660 6.880 101.840 ;
        RECT 7.050 101.660 7.360 101.840 ;
        RECT 7.530 101.660 7.840 101.840 ;
        RECT 8.010 101.660 8.320 101.840 ;
        RECT 8.490 101.660 8.800 101.840 ;
        RECT 8.970 101.660 9.280 101.840 ;
        RECT 9.450 101.660 9.760 101.840 ;
        RECT 9.930 101.660 10.240 101.840 ;
        RECT 10.410 101.660 10.720 101.840 ;
        RECT 10.890 101.660 11.200 101.840 ;
        RECT 11.370 101.660 11.680 101.840 ;
        RECT 11.850 101.660 12.160 101.840 ;
        RECT 12.330 101.660 12.640 101.840 ;
        RECT 12.810 101.660 13.120 101.840 ;
        RECT 13.290 101.660 13.600 101.840 ;
        RECT 13.770 101.660 14.080 101.840 ;
        RECT 14.250 101.660 14.560 101.840 ;
        RECT 14.730 101.660 15.040 101.840 ;
        RECT 15.210 101.660 15.520 101.840 ;
        RECT 15.690 101.660 16.000 101.840 ;
        RECT 16.170 101.660 16.480 101.840 ;
        RECT 16.650 101.660 16.960 101.840 ;
        RECT 17.130 101.660 17.440 101.840 ;
        RECT 17.610 101.660 17.920 101.840 ;
        RECT 18.090 101.660 18.400 101.840 ;
        RECT 18.570 101.660 18.880 101.840 ;
        RECT 19.050 101.660 19.360 101.840 ;
        RECT 19.530 101.660 19.840 101.840 ;
        RECT 20.010 101.660 20.320 101.840 ;
        RECT 20.490 101.660 20.800 101.840 ;
        RECT 20.970 101.660 21.280 101.840 ;
        RECT 21.450 101.660 21.760 101.840 ;
        RECT 21.930 101.660 22.240 101.840 ;
        RECT 22.410 101.660 22.720 101.840 ;
        RECT 22.890 101.660 23.200 101.840 ;
        RECT 23.370 101.660 23.680 101.840 ;
        RECT 23.850 101.660 24.160 101.840 ;
        RECT 24.330 101.660 24.640 101.840 ;
        RECT 24.810 101.660 25.120 101.840 ;
        RECT 25.290 101.660 25.600 101.840 ;
        RECT 25.770 101.660 26.080 101.840 ;
        RECT 26.250 101.660 26.560 101.840 ;
        RECT 26.730 101.660 27.040 101.840 ;
        RECT 27.210 101.660 27.520 101.840 ;
        RECT 27.690 101.660 28.000 101.840 ;
        RECT 28.170 101.660 28.480 101.840 ;
        RECT 28.650 101.660 28.960 101.840 ;
        RECT 29.130 101.660 29.440 101.840 ;
        RECT 29.610 101.660 29.920 101.840 ;
        RECT 30.090 101.660 30.400 101.840 ;
        RECT 30.570 101.660 30.880 101.840 ;
        RECT 31.050 101.660 31.360 101.840 ;
        RECT 31.530 101.660 31.840 101.840 ;
        RECT 32.010 101.660 32.320 101.840 ;
        RECT 32.490 101.660 32.800 101.840 ;
        RECT 32.970 101.660 33.280 101.840 ;
        RECT 33.450 101.660 33.760 101.840 ;
        RECT 33.930 101.660 34.240 101.840 ;
        RECT 34.410 101.660 34.720 101.840 ;
        RECT 34.890 101.660 35.200 101.840 ;
        RECT 35.370 101.660 35.680 101.840 ;
        RECT 35.850 101.660 36.160 101.840 ;
        RECT 36.330 101.660 36.640 101.840 ;
        RECT 36.810 101.660 37.120 101.840 ;
        RECT 37.290 101.660 37.600 101.840 ;
        RECT 37.770 101.660 38.080 101.840 ;
        RECT 38.250 101.660 38.560 101.840 ;
        RECT 38.730 101.660 39.040 101.840 ;
        RECT 39.210 101.660 39.520 101.840 ;
        RECT 39.690 101.660 40.000 101.840 ;
        RECT 40.170 101.660 40.320 101.840 ;
        RECT 40.800 101.660 40.960 101.840 ;
        RECT 41.130 101.660 41.440 101.840 ;
        RECT 41.610 101.660 41.920 101.840 ;
        RECT 42.090 101.660 42.400 101.840 ;
        RECT 42.570 101.660 42.880 101.840 ;
        RECT 43.050 101.660 43.360 101.840 ;
        RECT 43.530 101.660 43.840 101.840 ;
        RECT 44.010 101.660 44.320 101.840 ;
        RECT 44.490 101.660 44.800 101.840 ;
        RECT 44.970 101.660 45.280 101.840 ;
        RECT 45.450 101.660 45.760 101.840 ;
        RECT 45.930 101.660 46.240 101.840 ;
        RECT 46.410 101.660 46.720 101.840 ;
        RECT 46.890 101.660 47.200 101.840 ;
        RECT 47.370 101.660 47.680 101.840 ;
        RECT 47.850 101.660 48.160 101.840 ;
        RECT 48.330 101.660 48.640 101.840 ;
        RECT 48.810 101.660 49.120 101.840 ;
        RECT 49.290 101.660 49.600 101.840 ;
        RECT 49.770 101.660 50.080 101.840 ;
        RECT 50.250 101.660 50.560 101.840 ;
        RECT 50.730 101.660 51.040 101.840 ;
        RECT 51.210 101.660 51.520 101.840 ;
        RECT 51.690 101.660 52.000 101.840 ;
        RECT 52.170 101.660 52.480 101.840 ;
        RECT 52.650 101.660 52.960 101.840 ;
        RECT 53.130 101.660 53.440 101.840 ;
        RECT 53.610 101.660 53.920 101.840 ;
        RECT 54.090 101.660 54.400 101.840 ;
        RECT 54.570 101.660 54.880 101.840 ;
        RECT 55.050 101.660 55.360 101.840 ;
        RECT 55.530 101.660 55.840 101.840 ;
        RECT 56.010 101.660 56.320 101.840 ;
        RECT 56.490 101.660 56.800 101.840 ;
        RECT 56.970 101.660 57.280 101.840 ;
        RECT 57.450 101.660 57.760 101.840 ;
        RECT 57.930 101.660 58.240 101.840 ;
        RECT 58.410 101.660 58.720 101.840 ;
        RECT 58.890 101.660 59.200 101.840 ;
        RECT 59.370 101.660 59.680 101.840 ;
        RECT 59.850 101.660 60.160 101.840 ;
        RECT 60.330 101.660 60.640 101.840 ;
        RECT 60.810 101.660 60.960 101.840 ;
        RECT 61.440 101.660 61.600 101.840 ;
        RECT 61.770 101.660 62.080 101.840 ;
        RECT 62.250 101.660 62.560 101.840 ;
        RECT 62.730 101.660 63.040 101.840 ;
        RECT 63.210 101.660 63.520 101.840 ;
        RECT 63.690 101.660 64.000 101.840 ;
        RECT 64.170 101.660 64.480 101.840 ;
        RECT 64.650 101.660 64.960 101.840 ;
        RECT 65.130 101.660 65.440 101.840 ;
        RECT 65.610 101.660 65.920 101.840 ;
        RECT 66.090 101.660 66.400 101.840 ;
        RECT 66.570 101.660 66.880 101.840 ;
        RECT 67.050 101.660 67.360 101.840 ;
        RECT 67.530 101.660 67.840 101.840 ;
        RECT 68.010 101.660 68.320 101.840 ;
        RECT 68.490 101.660 68.800 101.840 ;
        RECT 68.970 101.660 69.280 101.840 ;
        RECT 69.450 101.660 69.760 101.840 ;
        RECT 69.930 101.660 70.240 101.840 ;
        RECT 70.410 101.660 70.720 101.840 ;
        RECT 70.890 101.660 71.200 101.840 ;
        RECT 71.370 101.660 71.680 101.840 ;
        RECT 71.850 101.660 72.160 101.840 ;
        RECT 72.330 101.660 72.640 101.840 ;
        RECT 72.810 101.660 73.120 101.840 ;
        RECT 73.290 101.660 73.600 101.840 ;
        RECT 73.770 101.660 74.080 101.840 ;
        RECT 74.250 101.660 74.560 101.840 ;
        RECT 74.730 101.660 75.040 101.840 ;
        RECT 75.210 101.660 75.520 101.840 ;
        RECT 75.690 101.660 76.000 101.840 ;
        RECT 76.170 101.660 76.480 101.840 ;
        RECT 76.650 101.660 76.960 101.840 ;
        RECT 77.130 101.660 77.440 101.840 ;
        RECT 77.610 101.660 77.920 101.840 ;
        RECT 78.090 101.660 78.400 101.840 ;
        RECT 78.570 101.660 78.880 101.840 ;
        RECT 79.050 101.660 79.360 101.840 ;
        RECT 79.530 101.660 79.840 101.840 ;
        RECT 80.010 101.660 80.320 101.840 ;
        RECT 80.490 101.660 80.800 101.840 ;
        RECT 80.970 101.660 81.280 101.840 ;
        RECT 81.450 101.660 81.760 101.840 ;
        RECT 81.930 101.660 82.240 101.840 ;
        RECT 82.410 101.660 82.720 101.840 ;
        RECT 82.890 101.660 83.200 101.840 ;
        RECT 83.370 101.660 83.680 101.840 ;
        RECT 83.850 101.660 84.160 101.840 ;
        RECT 84.330 101.660 84.640 101.840 ;
        RECT 84.810 101.660 85.120 101.840 ;
        RECT 85.290 101.660 85.600 101.840 ;
        RECT 85.770 101.660 86.080 101.840 ;
        RECT 86.250 101.660 86.560 101.840 ;
        RECT 86.730 101.660 87.040 101.840 ;
        RECT 87.210 101.660 87.520 101.840 ;
        RECT 87.690 101.660 88.000 101.840 ;
        RECT 88.170 101.660 88.480 101.840 ;
        RECT 88.650 101.660 88.960 101.840 ;
        RECT 89.130 101.660 89.440 101.840 ;
        RECT 89.610 101.660 89.920 101.840 ;
        RECT 90.090 101.660 90.400 101.840 ;
        RECT 90.570 101.660 90.880 101.840 ;
        RECT 91.050 101.660 91.360 101.840 ;
        RECT 91.530 101.660 91.840 101.840 ;
        RECT 92.010 101.660 92.320 101.840 ;
        RECT 92.490 101.660 92.800 101.840 ;
        RECT 92.970 101.660 93.280 101.840 ;
        RECT 93.450 101.660 93.760 101.840 ;
        RECT 93.930 101.660 94.240 101.840 ;
        RECT 94.410 101.660 94.720 101.840 ;
        RECT 94.890 101.660 95.200 101.840 ;
        RECT 95.370 101.660 95.680 101.840 ;
        RECT 95.850 101.660 96.160 101.840 ;
        RECT 96.330 101.660 96.640 101.840 ;
        RECT 96.810 101.660 97.120 101.840 ;
        RECT 97.290 101.660 97.600 101.840 ;
        RECT 97.770 101.660 98.080 101.840 ;
        RECT 98.250 101.660 98.560 101.840 ;
        RECT 98.730 101.660 99.040 101.840 ;
        RECT 99.210 101.660 99.520 101.840 ;
        RECT 99.690 101.660 100.000 101.840 ;
        RECT 100.170 101.660 100.480 101.840 ;
        RECT 100.650 101.660 100.960 101.840 ;
        RECT 101.130 101.660 101.440 101.840 ;
        RECT 101.610 101.660 101.920 101.840 ;
        RECT 102.090 101.660 102.400 101.840 ;
        RECT 102.570 101.660 102.880 101.840 ;
        RECT 103.050 101.660 103.360 101.840 ;
        RECT 103.530 101.660 103.840 101.840 ;
        RECT 104.010 101.660 104.320 101.840 ;
        RECT 104.490 101.660 104.800 101.840 ;
        RECT 104.970 101.660 105.280 101.840 ;
        RECT 105.450 101.660 105.760 101.840 ;
        RECT 105.930 101.660 106.240 101.840 ;
        RECT 106.410 101.660 106.720 101.840 ;
        RECT 106.890 101.660 107.200 101.840 ;
        RECT 107.370 101.660 107.680 101.840 ;
        RECT 107.850 101.660 108.160 101.840 ;
        RECT 108.330 101.660 108.640 101.840 ;
        RECT 108.810 101.660 109.120 101.840 ;
        RECT 109.290 101.660 109.600 101.840 ;
        RECT 109.770 101.660 110.080 101.840 ;
        RECT 110.250 101.660 110.560 101.840 ;
        RECT 110.730 101.660 111.040 101.840 ;
        RECT 111.210 101.660 111.520 101.840 ;
        RECT 111.690 101.660 112.000 101.840 ;
        RECT 112.170 101.660 112.480 101.840 ;
        RECT 112.650 101.660 112.960 101.840 ;
        RECT 113.130 101.660 113.440 101.840 ;
        RECT 113.610 101.660 113.920 101.840 ;
        RECT 114.090 101.660 114.400 101.840 ;
        RECT 114.570 101.660 114.880 101.840 ;
        RECT 115.050 101.660 115.360 101.840 ;
        RECT 115.530 101.660 115.840 101.840 ;
        RECT 116.010 101.660 116.320 101.840 ;
        RECT 116.490 101.660 116.800 101.840 ;
        RECT 116.970 101.660 117.280 101.840 ;
        RECT 117.450 101.660 117.760 101.840 ;
        RECT 117.930 101.660 118.240 101.840 ;
        RECT 118.410 101.660 118.720 101.840 ;
        RECT 118.890 101.660 119.200 101.840 ;
        RECT 119.370 101.660 119.680 101.840 ;
        RECT 119.850 101.660 120.160 101.840 ;
        RECT 120.330 101.660 120.640 101.840 ;
        RECT 120.810 101.660 120.960 101.840 ;
        RECT 121.440 101.660 121.600 101.840 ;
        RECT 121.770 101.660 122.080 101.840 ;
        RECT 122.250 101.660 122.560 101.840 ;
        RECT 122.730 101.660 123.040 101.840 ;
        RECT 123.210 101.660 123.520 101.840 ;
        RECT 123.690 101.660 124.000 101.840 ;
        RECT 124.170 101.660 124.480 101.840 ;
        RECT 124.650 101.660 124.960 101.840 ;
        RECT 125.130 101.660 125.440 101.840 ;
        RECT 125.610 101.660 125.920 101.840 ;
        RECT 126.090 101.660 126.400 101.840 ;
        RECT 126.570 101.660 126.880 101.840 ;
        RECT 127.050 101.660 127.360 101.840 ;
        RECT 127.530 101.660 127.840 101.840 ;
        RECT 128.010 101.660 128.320 101.840 ;
        RECT 128.490 101.660 128.800 101.840 ;
        RECT 128.970 101.660 129.280 101.840 ;
        RECT 129.450 101.660 129.760 101.840 ;
        RECT 129.930 101.660 130.240 101.840 ;
        RECT 130.410 101.660 130.720 101.840 ;
        RECT 130.890 101.660 131.200 101.840 ;
        RECT 131.370 101.660 131.680 101.840 ;
        RECT 131.850 101.660 132.160 101.840 ;
        RECT 132.330 101.660 132.640 101.840 ;
        RECT 132.810 101.660 133.120 101.840 ;
        RECT 133.290 101.660 133.600 101.840 ;
        RECT 133.770 101.660 134.080 101.840 ;
        RECT 134.250 101.660 134.560 101.840 ;
        RECT 134.730 101.660 135.040 101.840 ;
        RECT 135.210 101.660 135.520 101.840 ;
        RECT 135.690 101.660 136.000 101.840 ;
        RECT 136.170 101.660 136.480 101.840 ;
        RECT 136.650 101.660 136.960 101.840 ;
        RECT 137.130 101.660 137.440 101.840 ;
        RECT 137.610 101.660 137.920 101.840 ;
        RECT 138.090 101.660 138.400 101.840 ;
        RECT 138.570 101.660 138.880 101.840 ;
        RECT 139.050 101.660 139.360 101.840 ;
        RECT 139.530 101.660 139.840 101.840 ;
        RECT 140.010 101.660 140.320 101.840 ;
        RECT 140.490 101.660 140.800 101.840 ;
        RECT 140.970 101.660 141.280 101.840 ;
        RECT 141.450 101.660 141.760 101.840 ;
        RECT 141.930 101.660 142.080 101.840 ;
        RECT 6.340 101.360 9.070 101.390 ;
        RECT 6.340 101.190 6.510 101.360 ;
        RECT 6.680 101.190 6.950 101.360 ;
        RECT 7.120 101.190 7.360 101.360 ;
        RECT 7.530 101.190 7.790 101.360 ;
        RECT 7.960 101.190 8.230 101.360 ;
        RECT 8.400 101.190 8.640 101.360 ;
        RECT 8.810 101.190 9.070 101.360 ;
        RECT 6.340 100.390 9.070 101.190 ;
        RECT 10.180 101.360 12.910 101.390 ;
        RECT 10.180 101.190 10.350 101.360 ;
        RECT 10.520 101.190 10.790 101.360 ;
        RECT 10.960 101.190 11.200 101.360 ;
        RECT 11.370 101.190 11.630 101.360 ;
        RECT 11.800 101.190 12.070 101.360 ;
        RECT 12.240 101.190 12.480 101.360 ;
        RECT 12.650 101.190 12.910 101.360 ;
        RECT 10.180 100.390 12.910 101.190 ;
        RECT 13.610 101.350 15.220 101.380 ;
        RECT 16.870 101.350 18.120 101.380 ;
        RECT 18.890 101.350 20.500 101.380 ;
        RECT 13.610 101.180 13.660 101.350 ;
        RECT 13.830 101.180 14.100 101.350 ;
        RECT 14.270 101.180 14.540 101.350 ;
        RECT 14.710 101.180 14.950 101.350 ;
        RECT 15.120 101.180 15.220 101.350 ;
        RECT 13.610 100.900 15.220 101.180 ;
        RECT 13.920 100.500 15.220 100.900 ;
        RECT 6.500 99.720 6.830 100.390 ;
        RECT 7.230 99.070 7.560 100.050 ;
        RECT 7.780 99.720 8.110 100.390 ;
        RECT 8.510 99.070 8.840 100.050 ;
        RECT 10.340 99.720 10.670 100.390 ;
        RECT 11.070 99.070 11.400 100.050 ;
        RECT 11.620 99.720 11.950 100.390 ;
        RECT 12.350 99.070 12.680 100.050 ;
        RECT 13.920 99.720 14.250 100.500 ;
        RECT 6.260 98.190 9.000 99.070 ;
        RECT 6.260 98.020 6.470 98.190 ;
        RECT 6.640 98.020 6.910 98.190 ;
        RECT 7.080 98.020 7.320 98.190 ;
        RECT 7.490 98.020 7.750 98.190 ;
        RECT 7.920 98.020 8.190 98.190 ;
        RECT 8.360 98.020 8.600 98.190 ;
        RECT 8.770 98.020 9.000 98.190 ;
        RECT 6.260 98.000 9.000 98.020 ;
        RECT 10.100 98.190 12.840 99.070 ;
        RECT 14.460 99.060 14.790 100.050 ;
      LAYER li1 ;
        RECT 16.440 99.570 16.690 101.250 ;
      LAYER li1 ;
        RECT 17.040 101.180 17.230 101.350 ;
        RECT 17.400 101.180 17.590 101.350 ;
        RECT 17.760 101.180 17.950 101.350 ;
        RECT 16.870 100.810 18.120 101.180 ;
        RECT 18.300 100.630 18.550 101.250 ;
        RECT 18.890 101.180 18.940 101.350 ;
        RECT 19.110 101.180 19.380 101.350 ;
        RECT 19.550 101.180 19.820 101.350 ;
        RECT 19.990 101.180 20.230 101.350 ;
        RECT 20.400 101.180 20.500 101.350 ;
        RECT 18.890 100.900 20.500 101.180 ;
        RECT 17.000 100.460 18.550 100.630 ;
        RECT 17.000 100.000 17.330 100.460 ;
        RECT 10.100 98.020 10.310 98.190 ;
        RECT 10.480 98.020 10.750 98.190 ;
        RECT 10.920 98.020 11.160 98.190 ;
        RECT 11.330 98.020 11.590 98.190 ;
        RECT 11.760 98.020 12.030 98.190 ;
        RECT 12.200 98.020 12.440 98.190 ;
        RECT 12.610 98.020 12.840 98.190 ;
        RECT 10.100 98.000 12.840 98.020 ;
        RECT 13.690 98.190 15.140 99.060 ;
        RECT 13.690 98.020 13.940 98.190 ;
        RECT 14.110 98.020 14.300 98.190 ;
        RECT 14.470 98.020 14.740 98.190 ;
        RECT 14.910 98.020 15.140 98.190 ;
        RECT 13.690 97.990 15.140 98.020 ;
      LAYER li1 ;
        RECT 16.440 97.990 16.870 99.570 ;
      LAYER li1 ;
        RECT 17.050 98.240 17.610 99.570 ;
      LAYER li1 ;
        RECT 17.790 98.490 18.120 100.280 ;
      LAYER li1 ;
        RECT 18.300 98.740 18.550 100.460 ;
        RECT 19.200 100.500 20.500 100.900 ;
        RECT 22.170 101.350 22.760 101.380 ;
        RECT 22.170 101.180 22.200 101.350 ;
        RECT 22.370 101.180 22.560 101.350 ;
        RECT 22.730 101.180 22.760 101.350 ;
        RECT 24.100 101.360 26.830 101.390 ;
        RECT 19.200 99.720 19.530 100.500 ;
        RECT 22.170 100.420 22.760 101.180 ;
        RECT 19.740 99.060 20.070 100.050 ;
      LAYER li1 ;
        RECT 22.210 99.810 22.920 100.200 ;
        RECT 23.100 99.570 23.430 101.250 ;
      LAYER li1 ;
        RECT 24.100 101.190 24.270 101.360 ;
        RECT 24.440 101.190 24.710 101.360 ;
        RECT 24.880 101.190 25.120 101.360 ;
        RECT 25.290 101.190 25.550 101.360 ;
        RECT 25.720 101.190 25.990 101.360 ;
        RECT 26.160 101.190 26.400 101.360 ;
        RECT 26.570 101.190 26.830 101.360 ;
        RECT 24.100 100.390 26.830 101.190 ;
        RECT 28.890 101.350 29.480 101.380 ;
        RECT 28.890 101.180 28.920 101.350 ;
        RECT 29.090 101.180 29.280 101.350 ;
        RECT 29.450 101.180 29.480 101.350 ;
        RECT 30.410 101.350 32.020 101.380 ;
        RECT 32.710 101.350 33.960 101.380 ;
        RECT 34.730 101.350 36.340 101.380 ;
        RECT 37.030 101.350 38.280 101.380 ;
        RECT 39.050 101.350 40.660 101.380 ;
        RECT 28.890 100.420 29.480 101.180 ;
        RECT 24.260 99.720 24.590 100.390 ;
        RECT 17.050 98.070 17.060 98.240 ;
        RECT 17.230 98.070 17.420 98.240 ;
        RECT 17.590 98.070 17.610 98.240 ;
        RECT 17.050 97.990 17.610 98.070 ;
        RECT 18.970 98.190 20.420 99.060 ;
        RECT 18.970 98.020 19.220 98.190 ;
        RECT 19.390 98.020 19.580 98.190 ;
        RECT 19.750 98.020 20.020 98.190 ;
        RECT 20.190 98.020 20.420 98.190 ;
        RECT 18.970 97.990 20.420 98.020 ;
        RECT 22.170 98.240 22.760 99.570 ;
        RECT 22.170 98.070 22.200 98.240 ;
        RECT 22.370 98.070 22.560 98.240 ;
        RECT 22.730 98.070 22.760 98.240 ;
        RECT 22.170 97.990 22.760 98.070 ;
      LAYER li1 ;
        RECT 23.040 97.990 23.430 99.570 ;
      LAYER li1 ;
        RECT 24.990 99.070 25.320 100.050 ;
        RECT 25.540 99.720 25.870 100.390 ;
        RECT 26.270 99.070 26.600 100.050 ;
      LAYER li1 ;
        RECT 28.930 99.810 29.640 100.200 ;
        RECT 29.820 99.570 30.150 101.250 ;
      LAYER li1 ;
        RECT 30.410 101.180 30.460 101.350 ;
        RECT 30.630 101.180 30.900 101.350 ;
        RECT 31.070 101.180 31.340 101.350 ;
        RECT 31.510 101.180 31.750 101.350 ;
        RECT 31.920 101.180 32.020 101.350 ;
        RECT 30.410 100.900 32.020 101.180 ;
        RECT 30.720 100.500 32.020 100.900 ;
        RECT 30.720 99.720 31.050 100.500 ;
        RECT 24.020 98.190 26.760 99.070 ;
        RECT 24.020 98.020 24.230 98.190 ;
        RECT 24.400 98.020 24.670 98.190 ;
        RECT 24.840 98.020 25.080 98.190 ;
        RECT 25.250 98.020 25.510 98.190 ;
        RECT 25.680 98.020 25.950 98.190 ;
        RECT 26.120 98.020 26.360 98.190 ;
        RECT 26.530 98.020 26.760 98.190 ;
        RECT 24.020 98.000 26.760 98.020 ;
        RECT 28.890 98.240 29.480 99.570 ;
        RECT 28.890 98.070 28.920 98.240 ;
        RECT 29.090 98.070 29.280 98.240 ;
        RECT 29.450 98.070 29.480 98.240 ;
        RECT 28.890 97.990 29.480 98.070 ;
      LAYER li1 ;
        RECT 29.760 97.990 30.150 99.570 ;
      LAYER li1 ;
        RECT 31.260 99.060 31.590 100.050 ;
      LAYER li1 ;
        RECT 32.280 99.570 32.530 101.250 ;
      LAYER li1 ;
        RECT 32.880 101.180 33.070 101.350 ;
        RECT 33.240 101.180 33.430 101.350 ;
        RECT 33.600 101.180 33.790 101.350 ;
        RECT 32.710 100.810 33.960 101.180 ;
        RECT 34.140 100.630 34.390 101.250 ;
        RECT 34.730 101.180 34.780 101.350 ;
        RECT 34.950 101.180 35.220 101.350 ;
        RECT 35.390 101.180 35.660 101.350 ;
        RECT 35.830 101.180 36.070 101.350 ;
        RECT 36.240 101.180 36.340 101.350 ;
        RECT 34.730 100.900 36.340 101.180 ;
        RECT 32.840 100.460 34.390 100.630 ;
        RECT 32.840 100.000 33.170 100.460 ;
        RECT 30.490 98.190 31.940 99.060 ;
        RECT 30.490 98.020 30.740 98.190 ;
        RECT 30.910 98.020 31.100 98.190 ;
        RECT 31.270 98.020 31.540 98.190 ;
        RECT 31.710 98.020 31.940 98.190 ;
        RECT 30.490 97.990 31.940 98.020 ;
      LAYER li1 ;
        RECT 32.280 97.990 32.710 99.570 ;
      LAYER li1 ;
        RECT 32.890 98.240 33.450 99.570 ;
      LAYER li1 ;
        RECT 33.630 98.490 33.960 100.280 ;
      LAYER li1 ;
        RECT 34.140 98.740 34.390 100.460 ;
        RECT 35.040 100.500 36.340 100.900 ;
        RECT 35.040 99.720 35.370 100.500 ;
        RECT 35.580 99.060 35.910 100.050 ;
      LAYER li1 ;
        RECT 36.600 99.570 36.850 101.250 ;
      LAYER li1 ;
        RECT 37.200 101.180 37.390 101.350 ;
        RECT 37.560 101.180 37.750 101.350 ;
        RECT 37.920 101.180 38.110 101.350 ;
        RECT 37.030 100.810 38.280 101.180 ;
        RECT 38.460 100.630 38.710 101.250 ;
        RECT 39.050 101.180 39.100 101.350 ;
        RECT 39.270 101.180 39.540 101.350 ;
        RECT 39.710 101.180 39.980 101.350 ;
        RECT 40.150 101.180 40.390 101.350 ;
        RECT 40.560 101.180 40.660 101.350 ;
        RECT 39.050 100.900 40.660 101.180 ;
        RECT 37.160 100.460 38.710 100.630 ;
        RECT 37.160 100.000 37.490 100.460 ;
        RECT 32.890 98.070 32.900 98.240 ;
        RECT 33.070 98.070 33.260 98.240 ;
        RECT 33.430 98.070 33.450 98.240 ;
        RECT 32.890 97.990 33.450 98.070 ;
        RECT 34.810 98.190 36.260 99.060 ;
        RECT 34.810 98.020 35.060 98.190 ;
        RECT 35.230 98.020 35.420 98.190 ;
        RECT 35.590 98.020 35.860 98.190 ;
        RECT 36.030 98.020 36.260 98.190 ;
        RECT 34.810 97.990 36.260 98.020 ;
      LAYER li1 ;
        RECT 36.600 97.990 37.030 99.570 ;
      LAYER li1 ;
        RECT 37.210 98.240 37.770 99.570 ;
      LAYER li1 ;
        RECT 37.950 98.490 38.280 100.280 ;
      LAYER li1 ;
        RECT 38.460 98.740 38.710 100.460 ;
        RECT 39.360 100.500 40.660 100.900 ;
        RECT 40.890 101.350 41.840 101.380 ;
        RECT 40.890 101.180 40.920 101.350 ;
        RECT 41.090 101.180 41.280 101.350 ;
        RECT 41.450 101.180 41.640 101.350 ;
        RECT 41.810 101.180 41.840 101.350 ;
        RECT 42.450 101.350 43.400 101.380 ;
        RECT 39.360 99.720 39.690 100.500 ;
        RECT 40.890 100.420 41.840 101.180 ;
      LAYER li1 ;
        RECT 42.020 100.540 42.270 101.250 ;
      LAYER li1 ;
        RECT 42.450 101.180 42.480 101.350 ;
        RECT 42.650 101.180 42.840 101.350 ;
        RECT 43.010 101.180 43.200 101.350 ;
        RECT 43.370 101.180 43.400 101.350 ;
        RECT 44.010 101.350 44.960 101.380 ;
        RECT 42.450 100.720 43.400 101.180 ;
      LAYER li1 ;
        RECT 43.580 100.540 43.830 101.250 ;
        RECT 42.020 100.370 43.830 100.540 ;
      LAYER li1 ;
        RECT 44.010 101.180 44.040 101.350 ;
        RECT 44.210 101.180 44.400 101.350 ;
        RECT 44.570 101.180 44.760 101.350 ;
        RECT 44.930 101.180 44.960 101.350 ;
        RECT 45.770 101.350 47.380 101.380 ;
        RECT 44.010 100.500 44.960 101.180 ;
      LAYER li1 ;
        RECT 42.020 100.200 42.190 100.370 ;
      LAYER li1 ;
        RECT 45.140 100.320 45.470 101.250 ;
        RECT 45.770 101.180 45.820 101.350 ;
        RECT 45.990 101.180 46.260 101.350 ;
        RECT 46.430 101.180 46.700 101.350 ;
        RECT 46.870 101.180 47.110 101.350 ;
        RECT 47.280 101.180 47.380 101.350 ;
        RECT 45.770 100.900 47.380 101.180 ;
        RECT 39.900 99.060 40.230 100.050 ;
      LAYER li1 ;
        RECT 40.930 99.970 42.190 100.200 ;
      LAYER li1 ;
        RECT 44.230 100.190 45.470 100.320 ;
        RECT 42.370 100.150 45.470 100.190 ;
        RECT 42.370 100.020 44.400 100.150 ;
      LAYER li1 ;
        RECT 42.020 99.840 42.190 99.970 ;
        RECT 42.020 99.670 43.910 99.840 ;
      LAYER li1 ;
        RECT 37.210 98.070 37.220 98.240 ;
        RECT 37.390 98.070 37.580 98.240 ;
        RECT 37.750 98.070 37.770 98.240 ;
        RECT 37.210 97.990 37.770 98.070 ;
        RECT 39.130 98.190 40.580 99.060 ;
        RECT 39.130 98.020 39.380 98.190 ;
        RECT 39.550 98.020 39.740 98.190 ;
        RECT 39.910 98.020 40.180 98.190 ;
        RECT 40.350 98.020 40.580 98.190 ;
        RECT 39.130 97.990 40.580 98.020 ;
        RECT 40.890 98.240 41.840 99.570 ;
        RECT 40.890 98.070 40.920 98.240 ;
        RECT 41.090 98.070 41.280 98.240 ;
        RECT 41.450 98.070 41.640 98.240 ;
        RECT 41.810 98.070 41.840 98.240 ;
        RECT 40.890 97.990 41.840 98.070 ;
      LAYER li1 ;
        RECT 42.020 97.990 42.270 99.670 ;
      LAYER li1 ;
        RECT 42.450 98.240 43.400 99.490 ;
        RECT 42.450 98.070 42.480 98.240 ;
        RECT 42.650 98.070 42.840 98.240 ;
        RECT 43.010 98.070 43.200 98.240 ;
        RECT 43.370 98.070 43.400 98.240 ;
        RECT 42.450 97.990 43.400 98.070 ;
      LAYER li1 ;
        RECT 43.580 97.990 43.910 99.670 ;
        RECT 44.690 99.630 45.020 99.970 ;
      LAYER li1 ;
        RECT 44.090 98.240 45.040 99.450 ;
        RECT 44.090 98.070 44.120 98.240 ;
        RECT 44.290 98.070 44.480 98.240 ;
        RECT 44.650 98.070 44.840 98.240 ;
        RECT 45.010 98.070 45.040 98.240 ;
        RECT 44.090 97.990 45.040 98.070 ;
        RECT 45.220 97.990 45.470 100.150 ;
        RECT 46.080 100.500 47.380 100.900 ;
        RECT 47.610 101.350 48.560 101.380 ;
        RECT 47.610 101.180 47.640 101.350 ;
        RECT 47.810 101.180 48.000 101.350 ;
        RECT 48.170 101.180 48.360 101.350 ;
        RECT 48.530 101.180 48.560 101.350 ;
        RECT 49.170 101.350 50.120 101.380 ;
        RECT 46.080 99.720 46.410 100.500 ;
        RECT 47.610 100.420 48.560 101.180 ;
      LAYER li1 ;
        RECT 48.740 100.540 48.990 101.250 ;
      LAYER li1 ;
        RECT 49.170 101.180 49.200 101.350 ;
        RECT 49.370 101.180 49.560 101.350 ;
        RECT 49.730 101.180 49.920 101.350 ;
        RECT 50.090 101.180 50.120 101.350 ;
        RECT 50.730 101.350 51.680 101.380 ;
        RECT 49.170 100.720 50.120 101.180 ;
      LAYER li1 ;
        RECT 50.300 100.540 50.550 101.250 ;
        RECT 48.740 100.370 50.550 100.540 ;
      LAYER li1 ;
        RECT 50.730 101.180 50.760 101.350 ;
        RECT 50.930 101.180 51.120 101.350 ;
        RECT 51.290 101.180 51.480 101.350 ;
        RECT 51.650 101.180 51.680 101.350 ;
        RECT 52.490 101.350 54.100 101.380 ;
        RECT 50.730 100.500 51.680 101.180 ;
      LAYER li1 ;
        RECT 48.740 100.200 48.910 100.370 ;
      LAYER li1 ;
        RECT 51.860 100.320 52.190 101.250 ;
        RECT 52.490 101.180 52.540 101.350 ;
        RECT 52.710 101.180 52.980 101.350 ;
        RECT 53.150 101.180 53.420 101.350 ;
        RECT 53.590 101.180 53.830 101.350 ;
        RECT 54.000 101.180 54.100 101.350 ;
        RECT 52.490 100.900 54.100 101.180 ;
        RECT 46.620 99.060 46.950 100.050 ;
      LAYER li1 ;
        RECT 47.650 99.970 48.910 100.200 ;
      LAYER li1 ;
        RECT 50.950 100.190 52.190 100.320 ;
        RECT 49.090 100.150 52.190 100.190 ;
        RECT 49.090 100.020 51.120 100.150 ;
      LAYER li1 ;
        RECT 48.740 99.840 48.910 99.970 ;
        RECT 48.740 99.670 50.630 99.840 ;
      LAYER li1 ;
        RECT 45.850 98.190 47.300 99.060 ;
        RECT 45.850 98.020 46.100 98.190 ;
        RECT 46.270 98.020 46.460 98.190 ;
        RECT 46.630 98.020 46.900 98.190 ;
        RECT 47.070 98.020 47.300 98.190 ;
        RECT 45.850 97.990 47.300 98.020 ;
        RECT 47.610 98.240 48.560 99.570 ;
        RECT 47.610 98.070 47.640 98.240 ;
        RECT 47.810 98.070 48.000 98.240 ;
        RECT 48.170 98.070 48.360 98.240 ;
        RECT 48.530 98.070 48.560 98.240 ;
        RECT 47.610 97.990 48.560 98.070 ;
      LAYER li1 ;
        RECT 48.740 97.990 48.990 99.670 ;
      LAYER li1 ;
        RECT 49.170 98.240 50.120 99.490 ;
        RECT 49.170 98.070 49.200 98.240 ;
        RECT 49.370 98.070 49.560 98.240 ;
        RECT 49.730 98.070 49.920 98.240 ;
        RECT 50.090 98.070 50.120 98.240 ;
        RECT 49.170 97.990 50.120 98.070 ;
      LAYER li1 ;
        RECT 50.300 97.990 50.630 99.670 ;
        RECT 51.410 99.630 51.740 99.970 ;
      LAYER li1 ;
        RECT 50.810 98.240 51.760 99.450 ;
        RECT 50.810 98.070 50.840 98.240 ;
        RECT 51.010 98.070 51.200 98.240 ;
        RECT 51.370 98.070 51.560 98.240 ;
        RECT 51.730 98.070 51.760 98.240 ;
        RECT 50.810 97.990 51.760 98.070 ;
        RECT 51.940 97.990 52.190 100.150 ;
        RECT 52.800 100.500 54.100 100.900 ;
        RECT 54.330 101.350 55.280 101.380 ;
        RECT 54.330 101.180 54.360 101.350 ;
        RECT 54.530 101.180 54.720 101.350 ;
        RECT 54.890 101.180 55.080 101.350 ;
        RECT 55.250 101.180 55.280 101.350 ;
        RECT 55.890 101.350 56.840 101.380 ;
        RECT 52.800 99.720 53.130 100.500 ;
        RECT 54.330 100.420 55.280 101.180 ;
      LAYER li1 ;
        RECT 55.460 100.540 55.710 101.250 ;
      LAYER li1 ;
        RECT 55.890 101.180 55.920 101.350 ;
        RECT 56.090 101.180 56.280 101.350 ;
        RECT 56.450 101.180 56.640 101.350 ;
        RECT 56.810 101.180 56.840 101.350 ;
        RECT 57.450 101.350 58.400 101.380 ;
        RECT 55.890 100.720 56.840 101.180 ;
      LAYER li1 ;
        RECT 57.020 100.540 57.270 101.250 ;
        RECT 55.460 100.370 57.270 100.540 ;
      LAYER li1 ;
        RECT 57.450 101.180 57.480 101.350 ;
        RECT 57.650 101.180 57.840 101.350 ;
        RECT 58.010 101.180 58.200 101.350 ;
        RECT 58.370 101.180 58.400 101.350 ;
        RECT 59.210 101.350 60.820 101.380 ;
        RECT 57.450 100.500 58.400 101.180 ;
      LAYER li1 ;
        RECT 55.460 100.200 55.630 100.370 ;
      LAYER li1 ;
        RECT 58.580 100.320 58.910 101.250 ;
        RECT 59.210 101.180 59.260 101.350 ;
        RECT 59.430 101.180 59.700 101.350 ;
        RECT 59.870 101.180 60.140 101.350 ;
        RECT 60.310 101.180 60.550 101.350 ;
        RECT 60.720 101.180 60.820 101.350 ;
        RECT 59.210 100.900 60.820 101.180 ;
        RECT 53.340 99.060 53.670 100.050 ;
      LAYER li1 ;
        RECT 54.370 99.970 55.630 100.200 ;
      LAYER li1 ;
        RECT 57.670 100.190 58.910 100.320 ;
        RECT 55.810 100.150 58.910 100.190 ;
        RECT 55.810 100.020 57.840 100.150 ;
      LAYER li1 ;
        RECT 55.460 99.840 55.630 99.970 ;
        RECT 55.460 99.670 57.350 99.840 ;
      LAYER li1 ;
        RECT 52.570 98.190 54.020 99.060 ;
        RECT 52.570 98.020 52.820 98.190 ;
        RECT 52.990 98.020 53.180 98.190 ;
        RECT 53.350 98.020 53.620 98.190 ;
        RECT 53.790 98.020 54.020 98.190 ;
        RECT 52.570 97.990 54.020 98.020 ;
        RECT 54.330 98.240 55.280 99.570 ;
        RECT 54.330 98.070 54.360 98.240 ;
        RECT 54.530 98.070 54.720 98.240 ;
        RECT 54.890 98.070 55.080 98.240 ;
        RECT 55.250 98.070 55.280 98.240 ;
        RECT 54.330 97.990 55.280 98.070 ;
      LAYER li1 ;
        RECT 55.460 97.990 55.710 99.670 ;
      LAYER li1 ;
        RECT 55.890 98.240 56.840 99.490 ;
        RECT 55.890 98.070 55.920 98.240 ;
        RECT 56.090 98.070 56.280 98.240 ;
        RECT 56.450 98.070 56.640 98.240 ;
        RECT 56.810 98.070 56.840 98.240 ;
        RECT 55.890 97.990 56.840 98.070 ;
      LAYER li1 ;
        RECT 57.020 97.990 57.350 99.670 ;
        RECT 58.130 99.630 58.460 99.970 ;
      LAYER li1 ;
        RECT 57.530 98.240 58.480 99.450 ;
        RECT 57.530 98.070 57.560 98.240 ;
        RECT 57.730 98.070 57.920 98.240 ;
        RECT 58.090 98.070 58.280 98.240 ;
        RECT 58.450 98.070 58.480 98.240 ;
        RECT 57.530 97.990 58.480 98.070 ;
        RECT 58.660 97.990 58.910 100.150 ;
        RECT 59.520 100.500 60.820 100.900 ;
        RECT 61.120 101.310 62.930 101.480 ;
        RECT 59.520 99.720 59.850 100.500 ;
        RECT 61.120 100.390 61.450 101.310 ;
      LAYER li1 ;
        RECT 61.700 100.390 62.230 101.130 ;
      LAYER li1 ;
        RECT 60.060 99.060 60.390 100.050 ;
      LAYER li1 ;
        RECT 61.090 99.880 61.510 100.210 ;
        RECT 61.700 99.820 61.870 100.390 ;
      LAYER li1 ;
        RECT 62.760 100.290 62.930 101.310 ;
        RECT 63.110 101.350 64.210 101.380 ;
        RECT 63.110 101.180 63.160 101.350 ;
        RECT 63.330 101.180 63.520 101.350 ;
        RECT 63.690 101.180 63.880 101.350 ;
        RECT 64.050 101.180 64.210 101.350 ;
        RECT 64.970 101.350 66.580 101.380 ;
        RECT 67.270 101.350 68.520 101.380 ;
        RECT 69.290 101.350 70.900 101.380 ;
        RECT 63.110 100.470 64.210 101.180 ;
        RECT 64.380 100.290 64.630 101.220 ;
        RECT 64.970 101.180 65.020 101.350 ;
        RECT 65.190 101.180 65.460 101.350 ;
        RECT 65.630 101.180 65.900 101.350 ;
        RECT 66.070 101.180 66.310 101.350 ;
        RECT 66.480 101.180 66.580 101.350 ;
        RECT 64.970 100.900 66.580 101.180 ;
      LAYER li1 ;
        RECT 62.050 100.000 62.560 100.210 ;
      LAYER li1 ;
        RECT 62.760 100.120 64.630 100.290 ;
        RECT 65.280 100.500 66.580 100.900 ;
      LAYER li1 ;
        RECT 61.700 99.650 62.760 99.820 ;
        RECT 62.490 99.570 62.760 99.650 ;
        RECT 63.210 99.630 63.720 99.940 ;
        RECT 63.970 99.630 64.680 99.940 ;
      LAYER li1 ;
        RECT 65.280 99.720 65.610 100.500 ;
        RECT 59.290 98.190 60.740 99.060 ;
        RECT 59.290 98.020 59.540 98.190 ;
        RECT 59.710 98.020 59.900 98.190 ;
        RECT 60.070 98.020 60.340 98.190 ;
        RECT 60.510 98.020 60.740 98.190 ;
        RECT 59.290 97.990 60.740 98.020 ;
        RECT 61.050 98.240 62.310 99.470 ;
      LAYER li1 ;
        RECT 62.490 98.490 63.010 99.570 ;
      LAYER li1 ;
        RECT 61.050 98.070 61.060 98.240 ;
        RECT 61.230 98.070 61.420 98.240 ;
        RECT 61.590 98.070 61.780 98.240 ;
        RECT 61.950 98.070 62.140 98.240 ;
        RECT 61.050 97.990 62.310 98.070 ;
      LAYER li1 ;
        RECT 62.840 97.990 63.010 98.490 ;
      LAYER li1 ;
        RECT 63.270 98.240 64.580 99.450 ;
        RECT 65.820 99.060 66.150 100.050 ;
      LAYER li1 ;
        RECT 66.840 99.570 67.090 101.250 ;
      LAYER li1 ;
        RECT 67.440 101.180 67.630 101.350 ;
        RECT 67.800 101.180 67.990 101.350 ;
        RECT 68.160 101.180 68.350 101.350 ;
        RECT 67.270 100.810 68.520 101.180 ;
        RECT 68.700 100.630 68.950 101.250 ;
        RECT 69.290 101.180 69.340 101.350 ;
        RECT 69.510 101.180 69.780 101.350 ;
        RECT 69.950 101.180 70.220 101.350 ;
        RECT 70.390 101.180 70.630 101.350 ;
        RECT 70.800 101.180 70.900 101.350 ;
        RECT 69.290 100.900 70.900 101.180 ;
        RECT 67.400 100.460 68.950 100.630 ;
        RECT 67.400 100.000 67.730 100.460 ;
        RECT 63.270 98.070 63.300 98.240 ;
        RECT 63.470 98.070 63.660 98.240 ;
        RECT 63.830 98.070 64.020 98.240 ;
        RECT 64.190 98.070 64.380 98.240 ;
        RECT 64.550 98.070 64.580 98.240 ;
        RECT 63.270 97.990 64.580 98.070 ;
        RECT 65.050 98.190 66.500 99.060 ;
        RECT 65.050 98.020 65.300 98.190 ;
        RECT 65.470 98.020 65.660 98.190 ;
        RECT 65.830 98.020 66.100 98.190 ;
        RECT 66.270 98.020 66.500 98.190 ;
        RECT 65.050 97.990 66.500 98.020 ;
      LAYER li1 ;
        RECT 66.840 97.990 67.270 99.570 ;
      LAYER li1 ;
        RECT 67.450 98.240 68.010 99.570 ;
      LAYER li1 ;
        RECT 68.190 98.490 68.520 100.280 ;
      LAYER li1 ;
        RECT 68.700 98.740 68.950 100.460 ;
        RECT 69.600 100.500 70.900 100.900 ;
        RECT 72.570 101.350 73.160 101.380 ;
        RECT 72.570 101.180 72.600 101.350 ;
        RECT 72.770 101.180 72.960 101.350 ;
        RECT 73.130 101.180 73.160 101.350 ;
        RECT 73.840 101.350 74.790 101.380 ;
        RECT 69.600 99.720 69.930 100.500 ;
        RECT 72.570 100.420 73.160 101.180 ;
      LAYER li1 ;
        RECT 73.410 100.320 73.660 101.250 ;
      LAYER li1 ;
        RECT 73.840 101.180 73.870 101.350 ;
        RECT 74.040 101.180 74.230 101.350 ;
        RECT 74.400 101.180 74.590 101.350 ;
        RECT 74.760 101.180 74.790 101.350 ;
        RECT 76.010 101.350 77.620 101.380 ;
        RECT 73.840 100.500 74.790 101.180 ;
      LAYER li1 ;
        RECT 74.970 100.320 75.240 101.250 ;
      LAYER li1 ;
        RECT 76.010 101.180 76.060 101.350 ;
        RECT 76.230 101.180 76.500 101.350 ;
        RECT 76.670 101.180 76.940 101.350 ;
        RECT 77.110 101.180 77.350 101.350 ;
        RECT 77.520 101.180 77.620 101.350 ;
        RECT 76.010 100.900 77.620 101.180 ;
        RECT 70.140 99.060 70.470 100.050 ;
      LAYER li1 ;
        RECT 72.610 99.630 72.910 100.220 ;
        RECT 73.410 100.150 75.240 100.320 ;
        RECT 73.090 99.630 74.280 99.970 ;
      LAYER li1 ;
        RECT 67.450 98.070 67.460 98.240 ;
        RECT 67.630 98.070 67.820 98.240 ;
        RECT 67.990 98.070 68.010 98.240 ;
        RECT 67.450 97.990 68.010 98.070 ;
        RECT 69.370 98.190 70.820 99.060 ;
        RECT 69.370 98.020 69.620 98.190 ;
        RECT 69.790 98.020 69.980 98.190 ;
        RECT 70.150 98.020 70.420 98.190 ;
        RECT 70.590 98.020 70.820 98.190 ;
        RECT 69.370 97.990 70.820 98.020 ;
        RECT 72.570 98.240 74.240 99.450 ;
      LAYER li1 ;
        RECT 74.460 98.490 74.790 99.970 ;
      LAYER li1 ;
        RECT 72.570 98.070 72.600 98.240 ;
        RECT 72.770 98.070 72.960 98.240 ;
        RECT 73.130 98.070 73.320 98.240 ;
        RECT 73.490 98.070 73.680 98.240 ;
        RECT 73.850 98.070 74.040 98.240 ;
        RECT 74.210 98.070 74.240 98.240 ;
        RECT 72.570 97.990 74.240 98.070 ;
      LAYER li1 ;
        RECT 74.970 97.990 75.240 100.150 ;
      LAYER li1 ;
        RECT 76.320 100.500 77.620 100.900 ;
        RECT 77.850 101.350 78.800 101.380 ;
        RECT 77.850 101.180 77.880 101.350 ;
        RECT 78.050 101.180 78.240 101.350 ;
        RECT 78.410 101.180 78.600 101.350 ;
        RECT 78.770 101.180 78.800 101.350 ;
        RECT 79.410 101.350 80.360 101.380 ;
        RECT 76.320 99.720 76.650 100.500 ;
        RECT 77.850 100.420 78.800 101.180 ;
      LAYER li1 ;
        RECT 78.980 100.540 79.230 101.250 ;
      LAYER li1 ;
        RECT 79.410 101.180 79.440 101.350 ;
        RECT 79.610 101.180 79.800 101.350 ;
        RECT 79.970 101.180 80.160 101.350 ;
        RECT 80.330 101.180 80.360 101.350 ;
        RECT 80.970 101.350 81.920 101.380 ;
        RECT 79.410 100.720 80.360 101.180 ;
      LAYER li1 ;
        RECT 80.540 100.540 80.790 101.250 ;
        RECT 78.980 100.370 80.790 100.540 ;
      LAYER li1 ;
        RECT 80.970 101.180 81.000 101.350 ;
        RECT 81.170 101.180 81.360 101.350 ;
        RECT 81.530 101.180 81.720 101.350 ;
        RECT 81.890 101.180 81.920 101.350 ;
        RECT 82.730 101.350 84.340 101.380 ;
        RECT 80.970 100.500 81.920 101.180 ;
      LAYER li1 ;
        RECT 78.980 100.200 79.150 100.370 ;
      LAYER li1 ;
        RECT 82.100 100.320 82.430 101.250 ;
        RECT 82.730 101.180 82.780 101.350 ;
        RECT 82.950 101.180 83.220 101.350 ;
        RECT 83.390 101.180 83.660 101.350 ;
        RECT 83.830 101.180 84.070 101.350 ;
        RECT 84.240 101.180 84.340 101.350 ;
        RECT 82.730 100.900 84.340 101.180 ;
        RECT 76.860 99.060 77.190 100.050 ;
      LAYER li1 ;
        RECT 77.890 99.970 79.150 100.200 ;
      LAYER li1 ;
        RECT 81.190 100.190 82.430 100.320 ;
        RECT 79.330 100.150 82.430 100.190 ;
        RECT 79.330 100.020 81.360 100.150 ;
      LAYER li1 ;
        RECT 78.980 99.840 79.150 99.970 ;
        RECT 78.980 99.670 80.870 99.840 ;
      LAYER li1 ;
        RECT 76.090 98.190 77.540 99.060 ;
        RECT 76.090 98.020 76.340 98.190 ;
        RECT 76.510 98.020 76.700 98.190 ;
        RECT 76.870 98.020 77.140 98.190 ;
        RECT 77.310 98.020 77.540 98.190 ;
        RECT 76.090 97.990 77.540 98.020 ;
        RECT 77.850 98.240 78.800 99.570 ;
        RECT 77.850 98.070 77.880 98.240 ;
        RECT 78.050 98.070 78.240 98.240 ;
        RECT 78.410 98.070 78.600 98.240 ;
        RECT 78.770 98.070 78.800 98.240 ;
        RECT 77.850 97.990 78.800 98.070 ;
      LAYER li1 ;
        RECT 78.980 97.990 79.230 99.670 ;
      LAYER li1 ;
        RECT 79.410 98.240 80.360 99.490 ;
        RECT 79.410 98.070 79.440 98.240 ;
        RECT 79.610 98.070 79.800 98.240 ;
        RECT 79.970 98.070 80.160 98.240 ;
        RECT 80.330 98.070 80.360 98.240 ;
        RECT 79.410 97.990 80.360 98.070 ;
      LAYER li1 ;
        RECT 80.540 97.990 80.870 99.670 ;
        RECT 81.650 99.630 81.980 99.970 ;
      LAYER li1 ;
        RECT 81.050 98.240 82.000 99.450 ;
        RECT 81.050 98.070 81.080 98.240 ;
        RECT 81.250 98.070 81.440 98.240 ;
        RECT 81.610 98.070 81.800 98.240 ;
        RECT 81.970 98.070 82.000 98.240 ;
        RECT 81.050 97.990 82.000 98.070 ;
        RECT 82.180 97.990 82.430 100.150 ;
        RECT 83.040 100.500 84.340 100.900 ;
        RECT 84.570 101.350 85.520 101.380 ;
        RECT 84.570 101.180 84.600 101.350 ;
        RECT 84.770 101.180 84.960 101.350 ;
        RECT 85.130 101.180 85.320 101.350 ;
        RECT 85.490 101.180 85.520 101.350 ;
        RECT 86.130 101.350 87.080 101.380 ;
        RECT 83.040 99.720 83.370 100.500 ;
        RECT 84.570 100.420 85.520 101.180 ;
      LAYER li1 ;
        RECT 85.700 100.540 85.950 101.250 ;
      LAYER li1 ;
        RECT 86.130 101.180 86.160 101.350 ;
        RECT 86.330 101.180 86.520 101.350 ;
        RECT 86.690 101.180 86.880 101.350 ;
        RECT 87.050 101.180 87.080 101.350 ;
        RECT 87.690 101.350 88.640 101.380 ;
        RECT 86.130 100.720 87.080 101.180 ;
      LAYER li1 ;
        RECT 87.260 100.540 87.510 101.250 ;
        RECT 85.700 100.370 87.510 100.540 ;
      LAYER li1 ;
        RECT 87.690 101.180 87.720 101.350 ;
        RECT 87.890 101.180 88.080 101.350 ;
        RECT 88.250 101.180 88.440 101.350 ;
        RECT 88.610 101.180 88.640 101.350 ;
        RECT 89.860 101.360 92.590 101.390 ;
        RECT 87.690 100.500 88.640 101.180 ;
      LAYER li1 ;
        RECT 85.700 100.200 85.870 100.370 ;
      LAYER li1 ;
        RECT 88.820 100.320 89.150 101.250 ;
        RECT 89.860 101.190 90.030 101.360 ;
        RECT 90.200 101.190 90.470 101.360 ;
        RECT 90.640 101.190 90.880 101.360 ;
        RECT 91.050 101.190 91.310 101.360 ;
        RECT 91.480 101.190 91.750 101.360 ;
        RECT 91.920 101.190 92.160 101.360 ;
        RECT 92.330 101.190 92.590 101.360 ;
        RECT 89.860 100.390 92.590 101.190 ;
        RECT 93.210 101.350 94.160 101.380 ;
        RECT 93.210 101.180 93.240 101.350 ;
        RECT 93.410 101.180 93.600 101.350 ;
        RECT 93.770 101.180 93.960 101.350 ;
        RECT 94.130 101.180 94.160 101.350 ;
        RECT 94.770 101.350 95.720 101.380 ;
        RECT 93.210 100.420 94.160 101.180 ;
      LAYER li1 ;
        RECT 94.340 100.540 94.590 101.250 ;
      LAYER li1 ;
        RECT 94.770 101.180 94.800 101.350 ;
        RECT 94.970 101.180 95.160 101.350 ;
        RECT 95.330 101.180 95.520 101.350 ;
        RECT 95.690 101.180 95.720 101.350 ;
        RECT 96.330 101.350 97.280 101.380 ;
        RECT 94.770 100.720 95.720 101.180 ;
      LAYER li1 ;
        RECT 95.900 100.540 96.150 101.250 ;
      LAYER li1 ;
        RECT 83.580 99.060 83.910 100.050 ;
      LAYER li1 ;
        RECT 84.610 99.970 85.870 100.200 ;
      LAYER li1 ;
        RECT 87.910 100.190 89.150 100.320 ;
        RECT 86.050 100.150 89.150 100.190 ;
        RECT 86.050 100.020 88.080 100.150 ;
      LAYER li1 ;
        RECT 85.700 99.840 85.870 99.970 ;
        RECT 85.700 99.670 87.590 99.840 ;
      LAYER li1 ;
        RECT 82.810 98.190 84.260 99.060 ;
        RECT 82.810 98.020 83.060 98.190 ;
        RECT 83.230 98.020 83.420 98.190 ;
        RECT 83.590 98.020 83.860 98.190 ;
        RECT 84.030 98.020 84.260 98.190 ;
        RECT 82.810 97.990 84.260 98.020 ;
        RECT 84.570 98.240 85.520 99.570 ;
        RECT 84.570 98.070 84.600 98.240 ;
        RECT 84.770 98.070 84.960 98.240 ;
        RECT 85.130 98.070 85.320 98.240 ;
        RECT 85.490 98.070 85.520 98.240 ;
        RECT 84.570 97.990 85.520 98.070 ;
      LAYER li1 ;
        RECT 85.700 97.990 85.950 99.670 ;
      LAYER li1 ;
        RECT 86.130 98.240 87.080 99.490 ;
        RECT 86.130 98.070 86.160 98.240 ;
        RECT 86.330 98.070 86.520 98.240 ;
        RECT 86.690 98.070 86.880 98.240 ;
        RECT 87.050 98.070 87.080 98.240 ;
        RECT 86.130 97.990 87.080 98.070 ;
      LAYER li1 ;
        RECT 87.260 97.990 87.590 99.670 ;
        RECT 88.370 99.630 88.700 99.970 ;
      LAYER li1 ;
        RECT 87.770 98.240 88.720 99.450 ;
        RECT 87.770 98.070 87.800 98.240 ;
        RECT 87.970 98.070 88.160 98.240 ;
        RECT 88.330 98.070 88.520 98.240 ;
        RECT 88.690 98.070 88.720 98.240 ;
        RECT 87.770 97.990 88.720 98.070 ;
        RECT 88.900 97.990 89.150 100.150 ;
        RECT 90.020 99.720 90.350 100.390 ;
        RECT 90.750 99.070 91.080 100.050 ;
        RECT 91.300 99.720 91.630 100.390 ;
      LAYER li1 ;
        RECT 94.340 100.370 96.150 100.540 ;
      LAYER li1 ;
        RECT 96.330 101.180 96.360 101.350 ;
        RECT 96.530 101.180 96.720 101.350 ;
        RECT 96.890 101.180 97.080 101.350 ;
        RECT 97.250 101.180 97.280 101.350 ;
        RECT 98.090 101.350 99.700 101.380 ;
        RECT 100.400 101.350 101.290 101.380 ;
        RECT 96.330 100.500 97.280 101.180 ;
      LAYER li1 ;
        RECT 94.340 100.200 94.510 100.370 ;
      LAYER li1 ;
        RECT 97.460 100.320 97.790 101.250 ;
        RECT 98.090 101.180 98.140 101.350 ;
        RECT 98.310 101.180 98.580 101.350 ;
        RECT 98.750 101.180 99.020 101.350 ;
        RECT 99.190 101.180 99.430 101.350 ;
        RECT 99.600 101.180 99.700 101.350 ;
        RECT 98.090 100.900 99.700 101.180 ;
        RECT 92.030 99.070 92.360 100.050 ;
      LAYER li1 ;
        RECT 93.250 99.970 94.510 100.200 ;
      LAYER li1 ;
        RECT 96.550 100.190 97.790 100.320 ;
        RECT 94.690 100.150 97.790 100.190 ;
        RECT 94.690 100.020 96.720 100.150 ;
      LAYER li1 ;
        RECT 94.340 99.840 94.510 99.970 ;
        RECT 94.340 99.670 96.230 99.840 ;
      LAYER li1 ;
        RECT 89.780 98.190 92.520 99.070 ;
        RECT 89.780 98.020 89.990 98.190 ;
        RECT 90.160 98.020 90.430 98.190 ;
        RECT 90.600 98.020 90.840 98.190 ;
        RECT 91.010 98.020 91.270 98.190 ;
        RECT 91.440 98.020 91.710 98.190 ;
        RECT 91.880 98.020 92.120 98.190 ;
        RECT 92.290 98.020 92.520 98.190 ;
        RECT 89.780 98.000 92.520 98.020 ;
        RECT 93.210 98.240 94.160 99.570 ;
        RECT 93.210 98.070 93.240 98.240 ;
        RECT 93.410 98.070 93.600 98.240 ;
        RECT 93.770 98.070 93.960 98.240 ;
        RECT 94.130 98.070 94.160 98.240 ;
        RECT 93.210 97.990 94.160 98.070 ;
      LAYER li1 ;
        RECT 94.340 97.990 94.590 99.670 ;
      LAYER li1 ;
        RECT 94.770 98.240 95.720 99.490 ;
        RECT 94.770 98.070 94.800 98.240 ;
        RECT 94.970 98.070 95.160 98.240 ;
        RECT 95.330 98.070 95.520 98.240 ;
        RECT 95.690 98.070 95.720 98.240 ;
        RECT 94.770 97.990 95.720 98.070 ;
      LAYER li1 ;
        RECT 95.900 97.990 96.230 99.670 ;
        RECT 97.010 99.630 97.340 99.970 ;
      LAYER li1 ;
        RECT 96.410 98.240 97.360 99.450 ;
        RECT 96.410 98.070 96.440 98.240 ;
        RECT 96.610 98.070 96.800 98.240 ;
        RECT 96.970 98.070 97.160 98.240 ;
        RECT 97.330 98.070 97.360 98.240 ;
        RECT 96.410 97.990 97.360 98.070 ;
        RECT 97.540 97.990 97.790 100.150 ;
        RECT 98.400 100.500 99.700 100.900 ;
        RECT 98.400 99.720 98.730 100.500 ;
        RECT 98.940 99.060 99.270 100.050 ;
        RECT 98.170 98.190 99.620 99.060 ;
        RECT 98.170 98.020 98.420 98.190 ;
        RECT 98.590 98.020 98.780 98.190 ;
        RECT 98.950 98.020 99.220 98.190 ;
        RECT 99.390 98.020 99.620 98.190 ;
        RECT 98.170 97.990 99.620 98.020 ;
      LAYER li1 ;
        RECT 99.970 97.990 100.220 101.250 ;
      LAYER li1 ;
        RECT 100.570 101.180 100.760 101.350 ;
        RECT 100.930 101.180 101.120 101.350 ;
        RECT 101.590 101.310 103.520 101.480 ;
        RECT 100.400 100.500 101.290 101.180 ;
        RECT 101.590 100.880 101.920 101.310 ;
        RECT 102.370 100.870 102.700 101.130 ;
        RECT 102.100 100.700 102.700 100.870 ;
        RECT 103.190 100.720 103.520 101.310 ;
        RECT 103.730 101.350 105.030 101.380 ;
        RECT 103.730 101.180 103.760 101.350 ;
        RECT 103.930 101.180 104.120 101.350 ;
        RECT 104.290 101.180 104.480 101.350 ;
        RECT 104.650 101.180 104.840 101.350 ;
        RECT 105.010 101.180 105.030 101.350 ;
        RECT 103.730 100.700 105.030 101.180 ;
        RECT 105.290 101.350 106.900 101.380 ;
        RECT 107.590 101.350 108.840 101.380 ;
        RECT 109.610 101.350 111.220 101.380 ;
        RECT 105.290 101.180 105.340 101.350 ;
        RECT 105.510 101.180 105.780 101.350 ;
        RECT 105.950 101.180 106.220 101.350 ;
        RECT 106.390 101.180 106.630 101.350 ;
        RECT 106.800 101.180 106.900 101.350 ;
        RECT 105.290 100.900 106.900 101.180 ;
        RECT 101.470 100.530 102.270 100.700 ;
        RECT 101.470 100.320 101.640 100.530 ;
      LAYER li1 ;
        RECT 102.880 100.520 103.550 100.540 ;
        RECT 102.450 100.350 104.720 100.520 ;
      LAYER li1 ;
        RECT 100.430 100.150 101.640 100.320 ;
      LAYER li1 ;
        RECT 101.820 100.180 102.620 100.350 ;
      LAYER li1 ;
        RECT 100.430 99.450 100.760 100.150 ;
      LAYER li1 ;
        RECT 101.820 99.970 101.990 100.180 ;
        RECT 104.390 100.170 104.720 100.350 ;
        RECT 101.260 99.690 101.990 99.970 ;
        RECT 102.800 99.630 103.090 100.170 ;
        RECT 103.330 99.840 104.040 100.170 ;
        RECT 104.310 100.000 104.720 100.170 ;
        RECT 104.390 99.730 104.720 100.000 ;
      LAYER li1 ;
        RECT 105.600 100.500 106.900 100.900 ;
        RECT 105.600 99.720 105.930 100.500 ;
        RECT 103.270 99.450 103.520 99.570 ;
        RECT 100.430 99.280 103.520 99.450 ;
        RECT 100.400 98.240 103.090 99.100 ;
        RECT 100.570 98.070 100.760 98.240 ;
        RECT 100.930 98.070 101.120 98.240 ;
        RECT 101.290 98.070 101.480 98.240 ;
        RECT 101.650 98.070 101.840 98.240 ;
        RECT 102.010 98.070 102.200 98.240 ;
        RECT 102.370 98.070 102.560 98.240 ;
        RECT 102.730 98.070 102.920 98.240 ;
        RECT 100.400 97.990 103.090 98.070 ;
        RECT 103.270 97.990 103.520 99.280 ;
        RECT 103.700 98.240 105.010 99.550 ;
        RECT 106.140 99.060 106.470 100.050 ;
      LAYER li1 ;
        RECT 107.160 99.570 107.410 101.250 ;
      LAYER li1 ;
        RECT 107.760 101.180 107.950 101.350 ;
        RECT 108.120 101.180 108.310 101.350 ;
        RECT 108.480 101.180 108.670 101.350 ;
        RECT 107.590 100.810 108.840 101.180 ;
        RECT 109.020 100.630 109.270 101.250 ;
        RECT 109.610 101.180 109.660 101.350 ;
        RECT 109.830 101.180 110.100 101.350 ;
        RECT 110.270 101.180 110.540 101.350 ;
        RECT 110.710 101.180 110.950 101.350 ;
        RECT 111.120 101.180 111.220 101.350 ;
        RECT 109.610 100.900 111.220 101.180 ;
        RECT 111.930 101.350 112.520 101.380 ;
        RECT 111.930 101.180 111.960 101.350 ;
        RECT 112.130 101.180 112.320 101.350 ;
        RECT 112.490 101.180 112.520 101.350 ;
        RECT 107.720 100.460 109.270 100.630 ;
        RECT 107.720 100.000 108.050 100.460 ;
        RECT 103.700 98.070 103.730 98.240 ;
        RECT 103.900 98.070 104.090 98.240 ;
        RECT 104.260 98.070 104.450 98.240 ;
        RECT 104.620 98.070 104.810 98.240 ;
        RECT 104.980 98.070 105.010 98.240 ;
        RECT 103.700 98.010 105.010 98.070 ;
        RECT 105.370 98.190 106.820 99.060 ;
        RECT 105.370 98.020 105.620 98.190 ;
        RECT 105.790 98.020 105.980 98.190 ;
        RECT 106.150 98.020 106.420 98.190 ;
        RECT 106.590 98.020 106.820 98.190 ;
        RECT 105.370 97.990 106.820 98.020 ;
      LAYER li1 ;
        RECT 107.160 97.990 107.590 99.570 ;
      LAYER li1 ;
        RECT 107.770 98.240 108.330 99.570 ;
      LAYER li1 ;
        RECT 108.510 98.490 108.840 100.280 ;
      LAYER li1 ;
        RECT 109.020 98.740 109.270 100.460 ;
        RECT 109.920 100.500 111.220 100.900 ;
        RECT 109.920 99.720 110.250 100.500 ;
        RECT 111.480 100.450 111.740 101.130 ;
        RECT 111.930 100.630 112.520 101.180 ;
        RECT 112.700 101.310 113.650 101.480 ;
        RECT 113.830 101.350 114.370 101.380 ;
        RECT 112.700 100.450 112.870 101.310 ;
        RECT 111.480 100.280 112.870 100.450 ;
        RECT 110.460 99.060 110.790 100.050 ;
        RECT 107.770 98.070 107.780 98.240 ;
        RECT 107.950 98.070 108.140 98.240 ;
        RECT 108.310 98.070 108.330 98.240 ;
        RECT 107.770 97.990 108.330 98.070 ;
        RECT 109.690 98.190 111.140 99.060 ;
        RECT 109.690 98.020 109.940 98.190 ;
        RECT 110.110 98.020 110.300 98.190 ;
        RECT 110.470 98.020 110.740 98.190 ;
        RECT 110.910 98.020 111.140 98.190 ;
        RECT 109.690 97.990 111.140 98.020 ;
        RECT 111.480 98.010 111.730 100.280 ;
        RECT 112.540 99.850 112.870 100.280 ;
      LAYER li1 ;
        RECT 111.910 99.000 112.240 99.670 ;
      LAYER li1 ;
        RECT 113.050 99.470 113.300 101.130 ;
        RECT 113.480 100.570 113.650 101.310 ;
        RECT 114.000 101.180 114.190 101.350 ;
        RECT 114.360 101.180 114.370 101.350 ;
        RECT 116.220 101.350 117.170 101.380 ;
        RECT 113.830 100.750 114.370 101.180 ;
        RECT 114.550 100.750 114.900 101.250 ;
        RECT 113.480 100.400 114.550 100.570 ;
      LAYER li1 ;
        RECT 113.870 99.650 114.200 100.220 ;
      LAYER li1 ;
        RECT 113.050 99.300 114.200 99.470 ;
        RECT 111.910 98.240 112.860 98.820 ;
        RECT 113.050 98.800 113.370 99.300 ;
        RECT 111.910 98.070 111.940 98.240 ;
        RECT 112.110 98.070 112.300 98.240 ;
        RECT 112.470 98.070 112.660 98.240 ;
        RECT 112.830 98.070 112.860 98.240 ;
        RECT 111.910 97.990 112.860 98.070 ;
        RECT 113.040 98.010 113.370 98.800 ;
        RECT 113.600 98.240 113.850 99.120 ;
        RECT 113.600 98.070 113.630 98.240 ;
        RECT 113.800 98.070 113.850 98.240 ;
        RECT 113.600 98.040 113.850 98.070 ;
        RECT 114.030 97.990 114.200 99.300 ;
        RECT 114.380 98.460 114.550 100.400 ;
        RECT 114.730 98.640 114.900 100.750 ;
        RECT 115.430 100.780 115.680 101.250 ;
        RECT 116.220 101.180 116.250 101.350 ;
        RECT 116.420 101.180 116.610 101.350 ;
        RECT 116.780 101.180 116.970 101.350 ;
        RECT 117.140 101.180 117.170 101.350 ;
        RECT 116.220 100.960 117.170 101.180 ;
        RECT 117.350 100.780 117.680 101.480 ;
        RECT 115.080 98.460 115.250 100.660 ;
        RECT 115.430 100.610 117.680 100.780 ;
        RECT 118.160 101.350 119.110 101.380 ;
        RECT 118.160 101.180 118.190 101.350 ;
        RECT 118.360 101.180 118.550 101.350 ;
        RECT 118.720 101.180 118.910 101.350 ;
        RECT 119.080 101.180 119.110 101.350 ;
        RECT 122.700 101.350 123.290 101.380 ;
        RECT 115.430 99.140 115.600 100.610 ;
        RECT 115.780 99.940 116.020 100.250 ;
        RECT 116.500 100.120 117.230 100.430 ;
        RECT 118.160 100.370 119.110 101.180 ;
      LAYER li1 ;
        RECT 119.650 100.910 122.520 101.190 ;
        RECT 119.290 100.740 122.520 100.910 ;
        RECT 119.290 100.190 119.460 100.740 ;
        RECT 122.250 100.710 122.520 100.740 ;
      LAYER li1 ;
        RECT 122.700 101.180 122.730 101.350 ;
        RECT 122.900 101.180 123.090 101.350 ;
        RECT 123.260 101.180 123.290 101.350 ;
        RECT 120.390 100.270 121.020 100.560 ;
        RECT 122.700 100.270 123.290 101.180 ;
        RECT 124.620 101.350 125.570 101.380 ;
        RECT 124.620 101.180 124.650 101.350 ;
        RECT 124.820 101.180 125.010 101.350 ;
        RECT 125.180 101.180 125.370 101.350 ;
        RECT 125.540 101.180 125.570 101.350 ;
      LAYER li1 ;
        RECT 118.530 99.950 119.460 100.190 ;
      LAYER li1 ;
        RECT 119.640 100.040 120.150 100.200 ;
        RECT 115.780 99.770 118.350 99.940 ;
        RECT 119.640 99.870 120.670 100.040 ;
        RECT 119.640 99.770 119.810 99.870 ;
        RECT 115.780 99.580 116.020 99.770 ;
        RECT 118.180 99.600 119.810 99.770 ;
        RECT 116.200 99.420 118.000 99.590 ;
        RECT 119.990 99.420 120.320 99.660 ;
        RECT 115.430 98.640 115.760 99.140 ;
        RECT 116.200 98.460 116.370 99.420 ;
        RECT 117.830 99.250 120.320 99.420 ;
        RECT 114.380 98.130 116.370 98.460 ;
        RECT 116.550 99.070 117.650 99.240 ;
        RECT 120.500 99.070 120.670 99.870 ;
        RECT 116.550 98.190 116.790 99.070 ;
        RECT 117.480 98.900 118.260 99.070 ;
        RECT 116.970 98.240 117.300 98.890 ;
        RECT 117.930 98.640 118.260 98.900 ;
        RECT 116.970 98.070 117.000 98.240 ;
        RECT 117.170 98.070 117.300 98.240 ;
        RECT 116.970 98.040 117.300 98.070 ;
        RECT 118.440 98.240 119.390 99.070 ;
        RECT 118.440 98.070 118.470 98.240 ;
        RECT 118.640 98.070 118.830 98.240 ;
        RECT 119.000 98.070 119.190 98.240 ;
        RECT 119.360 98.070 119.390 98.240 ;
        RECT 118.440 98.040 119.390 98.070 ;
        RECT 120.060 98.900 120.670 99.070 ;
        RECT 120.850 99.430 121.020 100.270 ;
        RECT 121.670 100.090 122.000 100.200 ;
        RECT 123.480 100.090 123.810 100.770 ;
        RECT 124.110 100.270 124.440 100.770 ;
        RECT 124.620 100.270 125.570 101.180 ;
        RECT 126.410 101.350 128.020 101.380 ;
        RECT 126.410 101.180 126.460 101.350 ;
        RECT 126.630 101.180 126.900 101.350 ;
        RECT 127.070 101.180 127.340 101.350 ;
        RECT 127.510 101.180 127.750 101.350 ;
        RECT 127.920 101.180 128.020 101.350 ;
        RECT 126.410 100.900 128.020 101.180 ;
        RECT 126.720 100.500 128.020 100.900 ;
        RECT 128.250 101.350 129.200 101.380 ;
        RECT 128.250 101.180 128.280 101.350 ;
        RECT 128.450 101.180 128.640 101.350 ;
        RECT 128.810 101.180 129.000 101.350 ;
        RECT 129.170 101.180 129.200 101.350 ;
        RECT 129.810 101.350 130.760 101.380 ;
        RECT 121.670 99.920 123.920 100.090 ;
        RECT 121.670 99.610 122.000 99.920 ;
        RECT 123.240 99.430 123.570 99.740 ;
        RECT 120.850 99.260 123.570 99.430 ;
        RECT 120.060 98.150 120.230 98.900 ;
        RECT 120.850 98.720 121.020 99.260 ;
        RECT 120.410 98.330 121.020 98.720 ;
        RECT 121.370 98.240 122.320 99.080 ;
        RECT 122.770 99.070 123.570 99.260 ;
        RECT 122.770 98.920 123.100 99.070 ;
        RECT 123.750 98.740 123.920 99.920 ;
        RECT 122.740 98.570 123.920 98.740 ;
        RECT 124.230 99.520 124.440 100.270 ;
        RECT 125.270 99.520 125.600 100.020 ;
        RECT 126.720 99.720 127.050 100.500 ;
        RECT 128.250 100.420 129.200 101.180 ;
      LAYER li1 ;
        RECT 129.380 100.540 129.630 101.250 ;
      LAYER li1 ;
        RECT 129.810 101.180 129.840 101.350 ;
        RECT 130.010 101.180 130.200 101.350 ;
        RECT 130.370 101.180 130.560 101.350 ;
        RECT 130.730 101.180 130.760 101.350 ;
        RECT 131.370 101.350 132.320 101.380 ;
        RECT 129.810 100.720 130.760 101.180 ;
      LAYER li1 ;
        RECT 130.940 100.540 131.190 101.250 ;
        RECT 129.380 100.370 131.190 100.540 ;
      LAYER li1 ;
        RECT 131.370 101.180 131.400 101.350 ;
        RECT 131.570 101.180 131.760 101.350 ;
        RECT 131.930 101.180 132.120 101.350 ;
        RECT 132.290 101.180 132.320 101.350 ;
        RECT 133.540 101.360 136.270 101.390 ;
        RECT 131.370 100.500 132.320 101.180 ;
      LAYER li1 ;
        RECT 129.380 100.200 129.550 100.370 ;
      LAYER li1 ;
        RECT 132.500 100.320 132.830 101.250 ;
        RECT 133.540 101.190 133.710 101.360 ;
        RECT 133.880 101.190 134.150 101.360 ;
        RECT 134.320 101.190 134.560 101.360 ;
        RECT 134.730 101.190 134.990 101.360 ;
        RECT 135.160 101.190 135.430 101.360 ;
        RECT 135.600 101.190 135.840 101.360 ;
        RECT 136.010 101.190 136.270 101.360 ;
        RECT 133.540 100.390 136.270 101.190 ;
        RECT 137.380 101.360 140.110 101.390 ;
        RECT 137.380 101.190 137.550 101.360 ;
        RECT 137.720 101.190 137.990 101.360 ;
        RECT 138.160 101.190 138.400 101.360 ;
        RECT 138.570 101.190 138.830 101.360 ;
        RECT 139.000 101.190 139.270 101.360 ;
        RECT 139.440 101.190 139.680 101.360 ;
        RECT 139.850 101.190 140.110 101.360 ;
        RECT 137.380 100.390 140.110 101.190 ;
        RECT 124.230 99.350 125.600 99.520 ;
        RECT 122.740 98.490 122.910 98.570 ;
        RECT 120.060 97.940 121.190 98.150 ;
        RECT 121.370 98.070 121.400 98.240 ;
        RECT 121.570 98.070 121.760 98.240 ;
        RECT 121.930 98.070 122.120 98.240 ;
        RECT 122.290 98.070 122.320 98.240 ;
        RECT 121.370 98.040 122.320 98.070 ;
        RECT 122.660 97.990 122.910 98.490 ;
        RECT 123.090 98.240 124.040 98.390 ;
        RECT 124.230 98.380 124.480 99.350 ;
        RECT 123.090 98.070 123.120 98.240 ;
        RECT 123.290 98.070 123.480 98.240 ;
        RECT 123.650 98.070 123.840 98.240 ;
        RECT 124.010 98.070 124.040 98.240 ;
        RECT 123.090 98.010 124.040 98.070 ;
        RECT 124.660 98.240 125.600 99.170 ;
        RECT 127.260 99.060 127.590 100.050 ;
      LAYER li1 ;
        RECT 128.290 99.970 129.550 100.200 ;
      LAYER li1 ;
        RECT 131.590 100.190 132.830 100.320 ;
        RECT 129.730 100.150 132.830 100.190 ;
        RECT 129.730 100.020 131.760 100.150 ;
      LAYER li1 ;
        RECT 129.380 99.840 129.550 99.970 ;
        RECT 129.380 99.670 131.270 99.840 ;
      LAYER li1 ;
        RECT 124.660 98.070 124.680 98.240 ;
        RECT 124.850 98.070 125.040 98.240 ;
        RECT 125.210 98.070 125.400 98.240 ;
        RECT 125.570 98.070 125.600 98.240 ;
        RECT 124.660 98.040 125.600 98.070 ;
        RECT 126.490 98.190 127.940 99.060 ;
        RECT 126.490 98.020 126.740 98.190 ;
        RECT 126.910 98.020 127.100 98.190 ;
        RECT 127.270 98.020 127.540 98.190 ;
        RECT 127.710 98.020 127.940 98.190 ;
        RECT 126.490 97.990 127.940 98.020 ;
        RECT 128.250 98.240 129.200 99.570 ;
        RECT 128.250 98.070 128.280 98.240 ;
        RECT 128.450 98.070 128.640 98.240 ;
        RECT 128.810 98.070 129.000 98.240 ;
        RECT 129.170 98.070 129.200 98.240 ;
        RECT 128.250 97.990 129.200 98.070 ;
      LAYER li1 ;
        RECT 129.380 97.990 129.630 99.670 ;
      LAYER li1 ;
        RECT 129.810 98.240 130.760 99.490 ;
        RECT 129.810 98.070 129.840 98.240 ;
        RECT 130.010 98.070 130.200 98.240 ;
        RECT 130.370 98.070 130.560 98.240 ;
        RECT 130.730 98.070 130.760 98.240 ;
        RECT 129.810 97.990 130.760 98.070 ;
      LAYER li1 ;
        RECT 130.940 97.990 131.270 99.670 ;
        RECT 132.050 99.630 132.380 99.970 ;
      LAYER li1 ;
        RECT 131.450 98.240 132.400 99.450 ;
        RECT 131.450 98.070 131.480 98.240 ;
        RECT 131.650 98.070 131.840 98.240 ;
        RECT 132.010 98.070 132.200 98.240 ;
        RECT 132.370 98.070 132.400 98.240 ;
        RECT 131.450 97.990 132.400 98.070 ;
        RECT 132.580 97.990 132.830 100.150 ;
        RECT 133.700 99.720 134.030 100.390 ;
        RECT 134.430 99.070 134.760 100.050 ;
        RECT 134.980 99.720 135.310 100.390 ;
        RECT 135.710 99.070 136.040 100.050 ;
        RECT 137.540 99.720 137.870 100.390 ;
        RECT 138.270 99.070 138.600 100.050 ;
        RECT 138.820 99.720 139.150 100.390 ;
        RECT 139.550 99.070 139.880 100.050 ;
        RECT 133.460 98.190 136.200 99.070 ;
        RECT 133.460 98.020 133.670 98.190 ;
        RECT 133.840 98.020 134.110 98.190 ;
        RECT 134.280 98.020 134.520 98.190 ;
        RECT 134.690 98.020 134.950 98.190 ;
        RECT 135.120 98.020 135.390 98.190 ;
        RECT 135.560 98.020 135.800 98.190 ;
        RECT 135.970 98.020 136.200 98.190 ;
        RECT 133.460 98.000 136.200 98.020 ;
        RECT 137.300 98.190 140.040 99.070 ;
        RECT 137.300 98.020 137.510 98.190 ;
        RECT 137.680 98.020 137.950 98.190 ;
        RECT 138.120 98.020 138.360 98.190 ;
        RECT 138.530 98.020 138.790 98.190 ;
        RECT 138.960 98.020 139.230 98.190 ;
        RECT 139.400 98.020 139.640 98.190 ;
        RECT 139.810 98.020 140.040 98.190 ;
        RECT 137.300 98.000 140.040 98.020 ;
        RECT 5.760 97.590 5.920 97.770 ;
        RECT 6.090 97.590 6.400 97.770 ;
        RECT 6.570 97.590 6.880 97.770 ;
        RECT 7.050 97.590 7.360 97.770 ;
        RECT 7.530 97.590 7.840 97.770 ;
        RECT 8.010 97.590 8.320 97.770 ;
        RECT 8.490 97.590 8.800 97.770 ;
        RECT 8.970 97.590 9.280 97.770 ;
        RECT 9.450 97.590 9.760 97.770 ;
        RECT 9.930 97.590 10.240 97.770 ;
        RECT 10.410 97.590 10.720 97.770 ;
        RECT 10.890 97.590 11.200 97.770 ;
        RECT 11.370 97.590 11.680 97.770 ;
        RECT 11.850 97.590 12.160 97.770 ;
        RECT 12.330 97.590 12.640 97.770 ;
        RECT 12.810 97.590 13.120 97.770 ;
        RECT 13.290 97.590 13.600 97.770 ;
        RECT 13.770 97.590 14.080 97.770 ;
        RECT 14.250 97.590 14.560 97.770 ;
        RECT 14.730 97.590 15.040 97.770 ;
        RECT 15.210 97.590 15.520 97.770 ;
        RECT 15.690 97.590 16.000 97.770 ;
        RECT 16.170 97.590 16.480 97.770 ;
        RECT 16.650 97.590 16.960 97.770 ;
        RECT 17.130 97.590 17.440 97.770 ;
        RECT 17.610 97.590 17.920 97.770 ;
        RECT 18.090 97.590 18.400 97.770 ;
        RECT 18.570 97.590 18.880 97.770 ;
        RECT 19.050 97.590 19.360 97.770 ;
        RECT 19.530 97.590 19.840 97.770 ;
        RECT 20.010 97.590 20.320 97.770 ;
        RECT 20.490 97.590 20.800 97.770 ;
        RECT 20.970 97.590 21.280 97.770 ;
        RECT 21.450 97.760 21.760 97.770 ;
        RECT 21.930 97.760 22.240 97.770 ;
        RECT 21.450 97.590 21.600 97.760 ;
        RECT 22.080 97.590 22.240 97.760 ;
        RECT 22.410 97.590 22.720 97.770 ;
        RECT 22.890 97.590 23.200 97.770 ;
        RECT 23.370 97.590 23.680 97.770 ;
        RECT 23.850 97.590 24.160 97.770 ;
        RECT 24.330 97.590 24.640 97.770 ;
        RECT 24.810 97.590 25.120 97.770 ;
        RECT 25.290 97.590 25.600 97.770 ;
        RECT 25.770 97.590 26.080 97.770 ;
        RECT 26.250 97.590 26.560 97.770 ;
        RECT 26.730 97.590 27.040 97.770 ;
        RECT 27.210 97.590 27.520 97.770 ;
        RECT 27.690 97.590 28.000 97.770 ;
        RECT 28.170 97.760 28.480 97.770 ;
        RECT 28.650 97.760 28.960 97.770 ;
        RECT 28.170 97.590 28.320 97.760 ;
        RECT 28.800 97.590 28.960 97.760 ;
        RECT 29.130 97.590 29.440 97.770 ;
        RECT 29.610 97.590 29.920 97.770 ;
        RECT 30.090 97.590 30.400 97.770 ;
        RECT 30.570 97.590 30.880 97.770 ;
        RECT 31.050 97.590 31.360 97.770 ;
        RECT 31.530 97.590 31.840 97.770 ;
        RECT 32.010 97.590 32.320 97.770 ;
        RECT 32.490 97.760 32.640 97.770 ;
        RECT 33.120 97.760 33.280 97.770 ;
        RECT 32.490 97.590 32.800 97.760 ;
        RECT 32.970 97.590 33.280 97.760 ;
        RECT 33.450 97.590 33.760 97.770 ;
        RECT 33.930 97.590 34.240 97.770 ;
        RECT 34.410 97.590 34.720 97.770 ;
        RECT 34.890 97.590 35.200 97.770 ;
        RECT 35.370 97.590 35.680 97.770 ;
        RECT 35.850 97.590 36.160 97.770 ;
        RECT 36.330 97.590 36.640 97.770 ;
        RECT 36.810 97.590 37.120 97.770 ;
        RECT 37.290 97.590 37.600 97.770 ;
        RECT 37.770 97.590 38.080 97.770 ;
        RECT 38.250 97.590 38.560 97.770 ;
        RECT 38.730 97.590 39.040 97.770 ;
        RECT 39.210 97.590 39.520 97.770 ;
        RECT 39.690 97.590 40.000 97.770 ;
        RECT 40.170 97.590 40.480 97.770 ;
        RECT 40.650 97.590 40.960 97.770 ;
        RECT 41.130 97.590 41.440 97.770 ;
        RECT 41.610 97.590 41.920 97.770 ;
        RECT 42.090 97.590 42.400 97.770 ;
        RECT 42.570 97.590 42.880 97.770 ;
        RECT 43.050 97.590 43.360 97.770 ;
        RECT 43.530 97.590 43.840 97.770 ;
        RECT 44.010 97.590 44.320 97.770 ;
        RECT 44.490 97.590 44.800 97.770 ;
        RECT 44.970 97.590 45.280 97.770 ;
        RECT 45.450 97.590 45.760 97.770 ;
        RECT 45.930 97.590 46.240 97.770 ;
        RECT 46.410 97.590 46.720 97.770 ;
        RECT 46.890 97.590 47.200 97.770 ;
        RECT 47.370 97.590 47.680 97.770 ;
        RECT 47.850 97.590 48.160 97.770 ;
        RECT 48.330 97.590 48.640 97.770 ;
        RECT 48.810 97.590 49.120 97.770 ;
        RECT 49.290 97.590 49.600 97.770 ;
        RECT 49.770 97.590 50.080 97.770 ;
        RECT 50.250 97.590 50.560 97.770 ;
        RECT 50.730 97.590 51.040 97.770 ;
        RECT 51.210 97.590 51.520 97.770 ;
        RECT 51.690 97.590 52.000 97.770 ;
        RECT 52.170 97.590 52.480 97.770 ;
        RECT 52.650 97.590 52.960 97.770 ;
        RECT 53.130 97.590 53.440 97.770 ;
        RECT 53.610 97.590 53.920 97.770 ;
        RECT 54.090 97.590 54.400 97.770 ;
        RECT 54.570 97.590 54.880 97.770 ;
        RECT 55.050 97.590 55.360 97.770 ;
        RECT 55.530 97.590 55.840 97.770 ;
        RECT 56.010 97.590 56.320 97.770 ;
        RECT 56.490 97.590 56.800 97.770 ;
        RECT 56.970 97.590 57.280 97.770 ;
        RECT 57.450 97.590 57.760 97.770 ;
        RECT 57.930 97.590 58.240 97.770 ;
        RECT 58.410 97.590 58.720 97.770 ;
        RECT 58.890 97.590 59.200 97.770 ;
        RECT 59.370 97.590 59.680 97.770 ;
        RECT 59.850 97.590 60.160 97.770 ;
        RECT 60.330 97.590 60.640 97.770 ;
        RECT 60.810 97.590 61.120 97.770 ;
        RECT 61.290 97.590 61.600 97.770 ;
        RECT 61.770 97.590 62.080 97.770 ;
        RECT 62.250 97.590 62.560 97.770 ;
        RECT 62.730 97.590 63.040 97.770 ;
        RECT 63.210 97.590 63.520 97.770 ;
        RECT 63.690 97.590 64.000 97.770 ;
        RECT 64.170 97.590 64.480 97.770 ;
        RECT 64.650 97.590 64.960 97.770 ;
        RECT 65.130 97.590 65.440 97.770 ;
        RECT 65.610 97.590 65.920 97.770 ;
        RECT 66.090 97.590 66.400 97.770 ;
        RECT 66.570 97.590 66.880 97.770 ;
        RECT 67.050 97.590 67.360 97.770 ;
        RECT 67.530 97.590 67.840 97.770 ;
        RECT 68.010 97.590 68.320 97.770 ;
        RECT 68.490 97.590 68.800 97.770 ;
        RECT 68.970 97.590 69.280 97.770 ;
        RECT 69.450 97.590 69.760 97.770 ;
        RECT 69.930 97.590 70.240 97.770 ;
        RECT 70.410 97.590 70.720 97.770 ;
        RECT 70.890 97.590 71.200 97.770 ;
        RECT 71.370 97.590 71.680 97.770 ;
        RECT 71.850 97.760 72.160 97.770 ;
        RECT 72.330 97.760 72.640 97.770 ;
        RECT 71.850 97.590 72.000 97.760 ;
        RECT 72.480 97.590 72.640 97.760 ;
        RECT 72.810 97.590 73.120 97.770 ;
        RECT 73.290 97.590 73.600 97.770 ;
        RECT 73.770 97.760 73.920 97.770 ;
        RECT 74.400 97.760 74.560 97.770 ;
        RECT 73.770 97.590 74.080 97.760 ;
        RECT 74.250 97.590 74.560 97.760 ;
        RECT 74.730 97.590 75.040 97.770 ;
        RECT 75.210 97.590 75.520 97.770 ;
        RECT 75.690 97.590 76.000 97.770 ;
        RECT 76.170 97.590 76.480 97.770 ;
        RECT 76.650 97.590 76.960 97.770 ;
        RECT 77.130 97.590 77.440 97.770 ;
        RECT 77.610 97.590 77.920 97.770 ;
        RECT 78.090 97.590 78.400 97.770 ;
        RECT 78.570 97.590 78.880 97.770 ;
        RECT 79.050 97.590 79.360 97.770 ;
        RECT 79.530 97.590 79.840 97.770 ;
        RECT 80.010 97.590 80.320 97.770 ;
        RECT 80.490 97.590 80.800 97.770 ;
        RECT 80.970 97.590 81.280 97.770 ;
        RECT 81.450 97.590 81.760 97.770 ;
        RECT 81.930 97.590 82.240 97.770 ;
        RECT 82.410 97.590 82.720 97.770 ;
        RECT 82.890 97.590 83.200 97.770 ;
        RECT 83.370 97.590 83.680 97.770 ;
        RECT 83.850 97.590 84.160 97.770 ;
        RECT 84.330 97.590 84.640 97.770 ;
        RECT 84.810 97.590 85.120 97.770 ;
        RECT 85.290 97.590 85.600 97.770 ;
        RECT 85.770 97.590 86.080 97.770 ;
        RECT 86.250 97.590 86.560 97.770 ;
        RECT 86.730 97.590 87.040 97.770 ;
        RECT 87.210 97.590 87.520 97.770 ;
        RECT 87.690 97.590 88.000 97.770 ;
        RECT 88.170 97.590 88.480 97.770 ;
        RECT 88.650 97.590 88.960 97.770 ;
        RECT 89.130 97.590 89.440 97.770 ;
        RECT 89.610 97.590 89.920 97.770 ;
        RECT 90.090 97.590 90.400 97.770 ;
        RECT 90.570 97.590 90.880 97.770 ;
        RECT 91.050 97.590 91.360 97.770 ;
        RECT 91.530 97.590 91.840 97.770 ;
        RECT 92.010 97.590 92.320 97.770 ;
        RECT 92.490 97.590 92.800 97.770 ;
        RECT 92.970 97.590 93.280 97.770 ;
        RECT 93.450 97.590 93.760 97.770 ;
        RECT 93.930 97.590 94.240 97.770 ;
        RECT 94.410 97.590 94.720 97.770 ;
        RECT 94.890 97.590 95.200 97.770 ;
        RECT 95.370 97.590 95.680 97.770 ;
        RECT 95.850 97.590 96.160 97.770 ;
        RECT 96.330 97.590 96.640 97.770 ;
        RECT 96.810 97.590 97.120 97.770 ;
        RECT 97.290 97.590 97.600 97.770 ;
        RECT 97.770 97.590 98.080 97.770 ;
        RECT 98.250 97.760 98.400 97.770 ;
        RECT 98.880 97.760 99.040 97.770 ;
        RECT 98.250 97.590 98.560 97.760 ;
        RECT 98.730 97.590 99.040 97.760 ;
        RECT 99.210 97.590 99.520 97.770 ;
        RECT 99.690 97.590 100.000 97.770 ;
        RECT 100.170 97.590 100.480 97.770 ;
        RECT 100.650 97.590 100.960 97.770 ;
        RECT 101.130 97.590 101.440 97.770 ;
        RECT 101.610 97.590 101.920 97.770 ;
        RECT 102.090 97.590 102.400 97.770 ;
        RECT 102.570 97.590 102.880 97.770 ;
        RECT 103.050 97.590 103.360 97.770 ;
        RECT 103.530 97.590 103.840 97.770 ;
        RECT 104.010 97.590 104.320 97.770 ;
        RECT 104.490 97.590 104.800 97.770 ;
        RECT 104.970 97.590 105.280 97.770 ;
        RECT 105.450 97.590 105.760 97.770 ;
        RECT 105.930 97.590 106.240 97.770 ;
        RECT 106.410 97.590 106.720 97.770 ;
        RECT 106.890 97.590 107.200 97.770 ;
        RECT 107.370 97.590 107.680 97.770 ;
        RECT 107.850 97.590 108.160 97.770 ;
        RECT 108.330 97.590 108.640 97.770 ;
        RECT 108.810 97.590 109.120 97.770 ;
        RECT 109.290 97.590 109.600 97.770 ;
        RECT 109.770 97.590 110.080 97.770 ;
        RECT 110.250 97.590 110.560 97.770 ;
        RECT 110.730 97.590 111.040 97.770 ;
        RECT 111.210 97.590 111.520 97.770 ;
        RECT 111.690 97.590 112.000 97.770 ;
        RECT 112.170 97.590 112.480 97.770 ;
        RECT 112.650 97.590 112.960 97.770 ;
        RECT 113.130 97.590 113.440 97.770 ;
        RECT 113.610 97.590 113.920 97.770 ;
        RECT 114.090 97.590 114.400 97.770 ;
        RECT 114.570 97.590 114.880 97.770 ;
        RECT 115.050 97.590 115.360 97.770 ;
        RECT 115.530 97.590 115.840 97.770 ;
        RECT 116.010 97.590 116.320 97.770 ;
        RECT 116.490 97.590 116.800 97.770 ;
        RECT 116.970 97.590 117.280 97.770 ;
        RECT 117.450 97.590 117.760 97.770 ;
        RECT 117.930 97.590 118.240 97.770 ;
        RECT 118.410 97.590 118.720 97.770 ;
        RECT 118.890 97.590 119.200 97.770 ;
        RECT 119.370 97.590 119.680 97.770 ;
        RECT 119.850 97.590 120.160 97.770 ;
        RECT 120.330 97.590 120.640 97.770 ;
        RECT 120.810 97.760 120.960 97.770 ;
        RECT 121.440 97.760 121.600 97.770 ;
        RECT 120.810 97.590 121.120 97.760 ;
        RECT 121.290 97.590 121.600 97.760 ;
        RECT 121.770 97.590 122.080 97.770 ;
        RECT 122.250 97.590 122.560 97.770 ;
        RECT 122.730 97.590 123.040 97.770 ;
        RECT 123.210 97.590 123.520 97.770 ;
        RECT 123.690 97.590 124.000 97.770 ;
        RECT 124.170 97.590 124.480 97.770 ;
        RECT 124.650 97.590 124.960 97.770 ;
        RECT 125.130 97.590 125.440 97.770 ;
        RECT 125.610 97.590 125.920 97.770 ;
        RECT 126.090 97.590 126.400 97.770 ;
        RECT 126.570 97.590 126.880 97.770 ;
        RECT 127.050 97.590 127.360 97.770 ;
        RECT 127.530 97.590 127.840 97.770 ;
        RECT 128.010 97.590 128.320 97.770 ;
        RECT 128.490 97.590 128.800 97.770 ;
        RECT 128.970 97.590 129.280 97.770 ;
        RECT 129.450 97.590 129.760 97.770 ;
        RECT 129.930 97.590 130.240 97.770 ;
        RECT 130.410 97.590 130.720 97.770 ;
        RECT 130.890 97.590 131.200 97.770 ;
        RECT 131.370 97.590 131.680 97.770 ;
        RECT 131.850 97.590 132.160 97.770 ;
        RECT 132.330 97.590 132.640 97.770 ;
        RECT 132.810 97.590 133.120 97.770 ;
        RECT 133.290 97.590 133.600 97.770 ;
        RECT 133.770 97.590 134.080 97.770 ;
        RECT 134.250 97.590 134.560 97.770 ;
        RECT 134.730 97.590 135.040 97.770 ;
        RECT 135.210 97.590 135.520 97.770 ;
        RECT 135.690 97.590 136.000 97.770 ;
        RECT 136.170 97.590 136.480 97.770 ;
        RECT 136.650 97.590 136.960 97.770 ;
        RECT 137.130 97.590 137.440 97.770 ;
        RECT 137.610 97.590 137.920 97.770 ;
        RECT 138.090 97.590 138.400 97.770 ;
        RECT 138.570 97.590 138.880 97.770 ;
        RECT 139.050 97.590 139.360 97.770 ;
        RECT 139.530 97.590 139.840 97.770 ;
        RECT 140.010 97.590 140.320 97.770 ;
        RECT 140.490 97.590 140.800 97.770 ;
        RECT 140.970 97.590 141.280 97.770 ;
        RECT 141.450 97.760 141.760 97.770 ;
        RECT 141.930 97.760 142.080 97.770 ;
        RECT 141.450 97.590 141.600 97.760 ;
        RECT 6.390 97.290 6.980 97.320 ;
        RECT 6.390 97.120 6.420 97.290 ;
        RECT 6.590 97.120 6.780 97.290 ;
        RECT 6.950 97.120 6.980 97.290 ;
        RECT 5.870 96.140 6.200 97.070 ;
        RECT 6.390 96.340 6.980 97.120 ;
        RECT 7.160 97.250 8.600 97.420 ;
        RECT 7.160 96.140 7.330 97.250 ;
        RECT 5.870 95.970 7.330 96.140 ;
        RECT 5.870 94.110 6.140 95.970 ;
        RECT 7.000 95.470 7.330 95.970 ;
        RECT 7.510 95.760 7.760 97.070 ;
        RECT 8.000 96.450 8.250 97.070 ;
        RECT 8.430 96.800 8.600 97.250 ;
        RECT 8.780 97.290 9.110 97.320 ;
        RECT 8.780 97.120 8.810 97.290 ;
        RECT 8.980 97.120 9.110 97.290 ;
        RECT 8.780 96.980 9.110 97.120 ;
        RECT 9.290 97.250 11.030 97.420 ;
        RECT 9.290 96.800 9.460 97.250 ;
        RECT 8.430 96.630 9.460 96.800 ;
        RECT 9.640 96.450 9.810 97.070 ;
        RECT 10.340 96.810 10.670 97.070 ;
        RECT 8.000 96.280 9.810 96.450 ;
        RECT 9.990 96.280 10.210 96.610 ;
        RECT 9.640 96.100 9.810 96.280 ;
        RECT 7.510 95.530 8.040 95.760 ;
        RECT 7.510 94.610 7.780 95.530 ;
      LAYER li1 ;
        RECT 8.460 95.230 9.000 96.100 ;
      LAYER li1 ;
        RECT 9.640 95.930 9.860 96.100 ;
        RECT 6.320 93.980 7.270 94.610 ;
        RECT 7.450 94.110 7.780 94.610 ;
        RECT 7.960 93.980 8.550 94.860 ;
      LAYER li1 ;
        RECT 8.830 94.620 9.000 95.230 ;
        RECT 8.790 94.450 9.000 94.620 ;
        RECT 8.830 94.240 9.000 94.450 ;
        RECT 9.180 94.420 9.510 95.720 ;
      LAYER li1 ;
        RECT 9.690 94.940 9.860 95.930 ;
        RECT 10.040 95.760 10.210 96.280 ;
        RECT 10.390 96.110 10.560 96.810 ;
        RECT 10.860 96.660 11.030 97.250 ;
        RECT 11.210 97.290 12.160 97.320 ;
        RECT 11.210 97.120 11.240 97.290 ;
        RECT 11.410 97.120 11.600 97.290 ;
        RECT 11.770 97.120 11.960 97.290 ;
        RECT 12.130 97.120 12.160 97.290 ;
        RECT 11.210 96.840 12.160 97.120 ;
        RECT 12.340 97.250 13.370 97.420 ;
        RECT 12.340 96.660 12.510 97.250 ;
        RECT 10.860 96.610 12.510 96.660 ;
        RECT 10.740 96.490 12.510 96.610 ;
        RECT 10.740 96.290 11.070 96.490 ;
        RECT 12.690 96.310 13.020 97.070 ;
        RECT 13.200 96.890 13.370 97.250 ;
        RECT 13.550 97.290 14.500 97.370 ;
        RECT 13.550 97.120 13.580 97.290 ;
        RECT 13.750 97.120 13.940 97.290 ;
        RECT 14.110 97.120 14.300 97.290 ;
        RECT 14.470 97.120 14.500 97.290 ;
        RECT 13.550 97.070 14.500 97.120 ;
        RECT 13.200 96.720 15.010 96.890 ;
        RECT 11.250 96.140 13.020 96.310 ;
        RECT 11.250 96.110 11.420 96.140 ;
        RECT 10.390 95.940 11.420 96.110 ;
        RECT 14.330 95.960 14.660 96.540 ;
        RECT 10.040 95.530 11.070 95.760 ;
        RECT 10.740 95.040 11.070 95.530 ;
        RECT 11.250 95.260 11.420 95.940 ;
        RECT 11.600 95.790 14.660 95.960 ;
        RECT 11.600 95.440 11.930 95.790 ;
      LAYER li1 ;
        RECT 12.370 95.440 14.220 95.610 ;
      LAYER li1 ;
        RECT 11.250 95.090 13.870 95.260 ;
        RECT 9.690 94.440 9.960 94.940 ;
        RECT 11.250 94.860 11.420 95.090 ;
      LAYER li1 ;
        RECT 14.050 94.910 14.220 95.440 ;
      LAYER li1 ;
        RECT 10.410 94.690 11.420 94.860 ;
      LAYER li1 ;
        RECT 11.600 94.740 14.220 94.910 ;
      LAYER li1 ;
        RECT 10.410 94.440 10.740 94.690 ;
      LAYER li1 ;
        RECT 11.600 94.240 11.770 94.740 ;
        RECT 8.830 94.070 11.770 94.240 ;
      LAYER li1 ;
        RECT 12.920 93.980 13.870 94.560 ;
      LAYER li1 ;
        RECT 14.050 94.050 14.220 94.740 ;
      LAYER li1 ;
        RECT 14.400 94.940 14.660 95.790 ;
        RECT 14.840 95.370 15.010 96.720 ;
        RECT 15.190 96.460 15.440 97.370 ;
        RECT 16.250 97.290 17.200 97.320 ;
        RECT 18.030 97.290 18.930 97.320 ;
        RECT 16.250 97.120 16.280 97.290 ;
        RECT 16.450 97.120 16.640 97.290 ;
        RECT 16.810 97.120 17.000 97.290 ;
        RECT 17.170 97.120 17.200 97.290 ;
        RECT 18.200 97.120 18.390 97.290 ;
        RECT 18.560 97.120 18.750 97.290 ;
        RECT 18.920 97.120 18.930 97.290 ;
        RECT 15.190 96.290 16.070 96.460 ;
        RECT 16.250 96.290 17.200 97.120 ;
        RECT 17.600 96.320 17.850 96.790 ;
        RECT 18.030 96.500 18.930 97.120 ;
        RECT 19.540 97.290 20.480 97.350 ;
        RECT 19.540 97.120 19.560 97.290 ;
        RECT 19.730 97.120 19.920 97.290 ;
        RECT 20.090 97.120 20.280 97.290 ;
        RECT 20.450 97.120 20.480 97.290 ;
        RECT 15.390 95.550 15.720 96.050 ;
        RECT 15.900 95.970 16.070 96.290 ;
        RECT 17.600 96.150 18.610 96.320 ;
        RECT 15.900 95.800 18.260 95.970 ;
        RECT 14.840 95.200 16.010 95.370 ;
        RECT 14.400 94.230 14.730 94.940 ;
        RECT 15.190 94.400 15.520 94.940 ;
        RECT 15.730 94.700 16.010 95.200 ;
        RECT 16.190 94.400 16.360 95.800 ;
        RECT 18.440 95.620 18.610 96.150 ;
        RECT 16.570 95.450 18.610 95.620 ;
        RECT 16.570 95.060 16.900 95.450 ;
      LAYER li1 ;
        RECT 17.220 94.880 17.550 95.270 ;
      LAYER li1 ;
        RECT 15.190 94.230 16.360 94.400 ;
      LAYER li1 ;
        RECT 16.540 94.710 17.550 94.880 ;
        RECT 16.540 94.050 16.710 94.710 ;
      LAYER li1 ;
        RECT 18.380 94.610 18.610 95.450 ;
        RECT 19.110 95.620 19.360 96.620 ;
        RECT 19.540 95.810 20.480 97.120 ;
        RECT 19.110 95.290 20.480 95.620 ;
        RECT 19.110 95.110 19.320 95.290 ;
        RECT 18.990 94.610 19.320 95.110 ;
      LAYER li1 ;
        RECT 14.050 93.880 16.710 94.050 ;
      LAYER li1 ;
        RECT 16.890 93.980 17.840 94.530 ;
        RECT 18.380 94.110 18.710 94.610 ;
        RECT 19.500 93.980 20.450 95.110 ;
      LAYER li1 ;
        RECT 20.660 94.280 21.000 97.350 ;
      LAYER li1 ;
        RECT 21.620 97.340 24.360 97.360 ;
        RECT 21.620 97.170 21.830 97.340 ;
        RECT 22.000 97.170 22.270 97.340 ;
        RECT 22.440 97.170 22.680 97.340 ;
        RECT 22.850 97.170 23.110 97.340 ;
        RECT 23.280 97.170 23.550 97.340 ;
        RECT 23.720 97.170 23.960 97.340 ;
        RECT 24.130 97.170 24.360 97.340 ;
        RECT 21.620 96.290 24.360 97.170 ;
        RECT 25.050 97.290 26.310 97.370 ;
        RECT 25.050 97.120 25.060 97.290 ;
        RECT 25.230 97.120 25.420 97.290 ;
        RECT 25.590 97.120 25.780 97.290 ;
        RECT 25.950 97.120 26.140 97.290 ;
        RECT 21.860 94.970 22.190 95.640 ;
        RECT 22.590 95.310 22.920 96.290 ;
        RECT 23.140 94.970 23.470 95.640 ;
        RECT 23.870 95.310 24.200 96.290 ;
        RECT 25.050 95.890 26.310 97.120 ;
      LAYER li1 ;
        RECT 26.840 96.870 27.010 97.370 ;
        RECT 26.490 95.790 27.010 96.870 ;
      LAYER li1 ;
        RECT 27.270 97.290 28.580 97.370 ;
        RECT 27.270 97.120 27.300 97.290 ;
        RECT 27.470 97.120 27.660 97.290 ;
        RECT 27.830 97.120 28.020 97.290 ;
        RECT 28.190 97.120 28.380 97.290 ;
        RECT 28.550 97.120 28.580 97.290 ;
        RECT 27.270 95.910 28.580 97.120 ;
        RECT 29.300 97.340 32.040 97.360 ;
        RECT 29.300 97.170 29.510 97.340 ;
        RECT 29.680 97.170 29.950 97.340 ;
        RECT 30.120 97.170 30.360 97.340 ;
        RECT 30.530 97.170 30.790 97.340 ;
        RECT 30.960 97.170 31.230 97.340 ;
        RECT 31.400 97.170 31.640 97.340 ;
        RECT 31.810 97.170 32.040 97.340 ;
        RECT 29.300 96.290 32.040 97.170 ;
      LAYER li1 ;
        RECT 26.490 95.710 26.760 95.790 ;
        RECT 25.700 95.540 26.760 95.710 ;
        RECT 25.090 95.150 25.510 95.480 ;
        RECT 25.700 94.970 25.870 95.540 ;
        RECT 27.210 95.420 27.720 95.730 ;
        RECT 27.970 95.420 28.680 95.730 ;
        RECT 26.050 95.150 26.560 95.360 ;
      LAYER li1 ;
        RECT 26.760 95.070 28.630 95.240 ;
        RECT 21.700 93.970 24.430 94.970 ;
        RECT 25.120 94.050 25.450 94.970 ;
      LAYER li1 ;
        RECT 25.700 94.620 26.230 94.970 ;
        RECT 25.700 94.450 26.240 94.620 ;
        RECT 25.700 94.230 26.230 94.450 ;
      LAYER li1 ;
        RECT 26.760 94.050 26.930 95.070 ;
        RECT 25.120 93.880 26.930 94.050 ;
        RECT 27.110 93.980 28.210 94.890 ;
        RECT 28.380 94.140 28.630 95.070 ;
        RECT 29.540 94.970 29.870 95.640 ;
        RECT 30.270 95.310 30.600 96.290 ;
        RECT 30.820 94.970 31.150 95.640 ;
        RECT 31.550 95.310 31.880 96.290 ;
      LAYER li1 ;
        RECT 33.240 95.790 33.670 97.370 ;
      LAYER li1 ;
        RECT 33.850 97.290 34.410 97.370 ;
        RECT 33.850 97.120 33.860 97.290 ;
        RECT 34.030 97.120 34.220 97.290 ;
        RECT 34.390 97.120 34.410 97.290 ;
        RECT 33.850 95.790 34.410 97.120 ;
        RECT 35.770 97.340 37.220 97.370 ;
        RECT 35.770 97.170 36.020 97.340 ;
        RECT 36.190 97.170 36.380 97.340 ;
        RECT 36.550 97.170 36.820 97.340 ;
        RECT 36.990 97.170 37.220 97.340 ;
        RECT 29.380 93.970 32.110 94.970 ;
      LAYER li1 ;
        RECT 33.240 94.110 33.490 95.790 ;
      LAYER li1 ;
        RECT 33.800 94.900 34.130 95.360 ;
      LAYER li1 ;
        RECT 34.590 95.080 34.920 96.870 ;
      LAYER li1 ;
        RECT 35.100 94.900 35.350 96.620 ;
        RECT 35.770 96.300 37.220 97.170 ;
        RECT 33.800 94.730 35.350 94.900 ;
        RECT 33.670 93.980 34.920 94.550 ;
        RECT 35.100 94.110 35.350 94.730 ;
        RECT 36.000 94.860 36.330 95.640 ;
        RECT 36.540 95.310 36.870 96.300 ;
      LAYER li1 ;
        RECT 37.560 95.790 37.990 97.370 ;
      LAYER li1 ;
        RECT 38.170 97.290 38.730 97.370 ;
        RECT 38.170 97.120 38.180 97.290 ;
        RECT 38.350 97.120 38.540 97.290 ;
        RECT 38.710 97.120 38.730 97.290 ;
        RECT 38.170 95.790 38.730 97.120 ;
        RECT 40.090 97.340 41.540 97.370 ;
        RECT 40.090 97.170 40.340 97.340 ;
        RECT 40.510 97.170 40.700 97.340 ;
        RECT 40.870 97.170 41.140 97.340 ;
        RECT 41.310 97.170 41.540 97.340 ;
        RECT 36.000 94.460 37.300 94.860 ;
        RECT 35.690 93.980 37.300 94.460 ;
      LAYER li1 ;
        RECT 37.560 94.110 37.810 95.790 ;
      LAYER li1 ;
        RECT 38.120 94.900 38.450 95.360 ;
      LAYER li1 ;
        RECT 38.910 95.080 39.240 96.870 ;
      LAYER li1 ;
        RECT 39.420 94.900 39.670 96.620 ;
        RECT 40.090 96.300 41.540 97.170 ;
        RECT 41.850 97.290 42.800 97.370 ;
        RECT 41.850 97.120 41.880 97.290 ;
        RECT 42.050 97.120 42.240 97.290 ;
        RECT 42.410 97.120 42.600 97.290 ;
        RECT 42.770 97.120 42.800 97.290 ;
        RECT 38.120 94.730 39.670 94.900 ;
        RECT 37.990 93.980 39.240 94.550 ;
        RECT 39.420 94.110 39.670 94.730 ;
        RECT 40.320 94.860 40.650 95.640 ;
        RECT 40.860 95.310 41.190 96.300 ;
        RECT 41.850 95.790 42.800 97.120 ;
      LAYER li1 ;
        RECT 42.980 95.690 43.230 97.370 ;
      LAYER li1 ;
        RECT 43.410 97.290 44.360 97.370 ;
        RECT 43.410 97.120 43.440 97.290 ;
        RECT 43.610 97.120 43.800 97.290 ;
        RECT 43.970 97.120 44.160 97.290 ;
        RECT 44.330 97.120 44.360 97.290 ;
        RECT 43.410 95.870 44.360 97.120 ;
      LAYER li1 ;
        RECT 44.540 95.690 44.870 97.370 ;
      LAYER li1 ;
        RECT 45.050 97.290 46.000 97.370 ;
        RECT 45.050 97.120 45.080 97.290 ;
        RECT 45.250 97.120 45.440 97.290 ;
        RECT 45.610 97.120 45.800 97.290 ;
        RECT 45.970 97.120 46.000 97.290 ;
        RECT 45.050 95.910 46.000 97.120 ;
      LAYER li1 ;
        RECT 42.980 95.520 44.870 95.690 ;
        RECT 42.980 95.390 43.150 95.520 ;
        RECT 45.650 95.390 45.980 95.730 ;
        RECT 41.890 95.160 43.150 95.390 ;
      LAYER li1 ;
        RECT 43.330 95.210 45.360 95.340 ;
        RECT 46.180 95.210 46.430 97.370 ;
        RECT 46.810 97.340 48.260 97.370 ;
        RECT 46.810 97.170 47.060 97.340 ;
        RECT 47.230 97.170 47.420 97.340 ;
        RECT 47.590 97.170 47.860 97.340 ;
        RECT 48.030 97.170 48.260 97.340 ;
        RECT 46.810 96.300 48.260 97.170 ;
        RECT 48.570 97.290 49.520 97.370 ;
        RECT 48.570 97.120 48.600 97.290 ;
        RECT 48.770 97.120 48.960 97.290 ;
        RECT 49.130 97.120 49.320 97.290 ;
        RECT 49.490 97.120 49.520 97.290 ;
        RECT 43.330 95.170 46.430 95.210 ;
      LAYER li1 ;
        RECT 42.980 94.990 43.150 95.160 ;
      LAYER li1 ;
        RECT 45.190 95.040 46.430 95.170 ;
        RECT 40.320 94.460 41.620 94.860 ;
        RECT 40.010 93.980 41.620 94.460 ;
        RECT 41.850 93.980 42.800 94.940 ;
      LAYER li1 ;
        RECT 42.980 94.820 44.790 94.990 ;
        RECT 42.980 94.110 43.230 94.820 ;
      LAYER li1 ;
        RECT 43.410 93.980 44.360 94.640 ;
      LAYER li1 ;
        RECT 44.540 94.110 44.790 94.820 ;
      LAYER li1 ;
        RECT 44.970 93.980 45.920 94.860 ;
        RECT 46.100 94.110 46.430 95.040 ;
        RECT 47.040 94.860 47.370 95.640 ;
        RECT 47.580 95.310 47.910 96.300 ;
        RECT 48.570 95.790 49.520 97.120 ;
      LAYER li1 ;
        RECT 49.700 95.690 49.950 97.370 ;
      LAYER li1 ;
        RECT 50.130 97.290 51.080 97.370 ;
        RECT 50.130 97.120 50.160 97.290 ;
        RECT 50.330 97.120 50.520 97.290 ;
        RECT 50.690 97.120 50.880 97.290 ;
        RECT 51.050 97.120 51.080 97.290 ;
        RECT 50.130 95.870 51.080 97.120 ;
      LAYER li1 ;
        RECT 51.260 95.690 51.590 97.370 ;
      LAYER li1 ;
        RECT 51.770 97.290 52.720 97.370 ;
        RECT 51.770 97.120 51.800 97.290 ;
        RECT 51.970 97.120 52.160 97.290 ;
        RECT 52.330 97.120 52.520 97.290 ;
        RECT 52.690 97.120 52.720 97.290 ;
        RECT 51.770 95.910 52.720 97.120 ;
      LAYER li1 ;
        RECT 49.700 95.520 51.590 95.690 ;
        RECT 49.700 95.390 49.870 95.520 ;
        RECT 52.370 95.390 52.700 95.730 ;
        RECT 48.610 95.160 49.870 95.390 ;
      LAYER li1 ;
        RECT 50.050 95.210 52.080 95.340 ;
        RECT 52.900 95.210 53.150 97.370 ;
        RECT 53.530 97.340 54.980 97.370 ;
        RECT 53.530 97.170 53.780 97.340 ;
        RECT 53.950 97.170 54.140 97.340 ;
        RECT 54.310 97.170 54.580 97.340 ;
        RECT 54.750 97.170 54.980 97.340 ;
        RECT 53.530 96.300 54.980 97.170 ;
        RECT 55.290 97.290 56.240 97.370 ;
        RECT 55.290 97.120 55.320 97.290 ;
        RECT 55.490 97.120 55.680 97.290 ;
        RECT 55.850 97.120 56.040 97.290 ;
        RECT 56.210 97.120 56.240 97.290 ;
        RECT 50.050 95.170 53.150 95.210 ;
      LAYER li1 ;
        RECT 49.700 94.990 49.870 95.160 ;
      LAYER li1 ;
        RECT 51.910 95.040 53.150 95.170 ;
        RECT 47.040 94.460 48.340 94.860 ;
        RECT 46.730 93.980 48.340 94.460 ;
        RECT 48.570 93.980 49.520 94.940 ;
      LAYER li1 ;
        RECT 49.700 94.820 51.510 94.990 ;
        RECT 49.700 94.110 49.950 94.820 ;
      LAYER li1 ;
        RECT 50.130 93.980 51.080 94.640 ;
      LAYER li1 ;
        RECT 51.260 94.110 51.510 94.820 ;
      LAYER li1 ;
        RECT 51.690 93.980 52.640 94.860 ;
        RECT 52.820 94.110 53.150 95.040 ;
        RECT 53.760 94.860 54.090 95.640 ;
        RECT 54.300 95.310 54.630 96.300 ;
        RECT 55.290 95.790 56.240 97.120 ;
      LAYER li1 ;
        RECT 56.420 95.690 56.670 97.370 ;
      LAYER li1 ;
        RECT 56.850 97.290 57.800 97.370 ;
        RECT 56.850 97.120 56.880 97.290 ;
        RECT 57.050 97.120 57.240 97.290 ;
        RECT 57.410 97.120 57.600 97.290 ;
        RECT 57.770 97.120 57.800 97.290 ;
        RECT 56.850 95.870 57.800 97.120 ;
      LAYER li1 ;
        RECT 57.980 95.690 58.310 97.370 ;
      LAYER li1 ;
        RECT 58.490 97.290 59.440 97.370 ;
        RECT 58.490 97.120 58.520 97.290 ;
        RECT 58.690 97.120 58.880 97.290 ;
        RECT 59.050 97.120 59.240 97.290 ;
        RECT 59.410 97.120 59.440 97.290 ;
        RECT 58.490 95.910 59.440 97.120 ;
      LAYER li1 ;
        RECT 56.420 95.520 58.310 95.690 ;
        RECT 56.420 95.390 56.590 95.520 ;
        RECT 59.090 95.390 59.420 95.730 ;
        RECT 55.330 95.160 56.590 95.390 ;
      LAYER li1 ;
        RECT 56.770 95.210 58.800 95.340 ;
        RECT 59.620 95.210 59.870 97.370 ;
        RECT 60.250 97.340 61.700 97.370 ;
        RECT 60.250 97.170 60.500 97.340 ;
        RECT 60.670 97.170 60.860 97.340 ;
        RECT 61.030 97.170 61.300 97.340 ;
        RECT 61.470 97.170 61.700 97.340 ;
        RECT 60.250 96.300 61.700 97.170 ;
        RECT 56.770 95.170 59.870 95.210 ;
      LAYER li1 ;
        RECT 56.420 94.990 56.590 95.160 ;
      LAYER li1 ;
        RECT 58.630 95.040 59.870 95.170 ;
        RECT 53.760 94.460 55.060 94.860 ;
        RECT 53.450 93.980 55.060 94.460 ;
        RECT 55.290 93.980 56.240 94.940 ;
      LAYER li1 ;
        RECT 56.420 94.820 58.230 94.990 ;
        RECT 56.420 94.110 56.670 94.820 ;
      LAYER li1 ;
        RECT 56.850 93.980 57.800 94.640 ;
      LAYER li1 ;
        RECT 57.980 94.110 58.230 94.820 ;
      LAYER li1 ;
        RECT 58.410 93.980 59.360 94.860 ;
        RECT 59.540 94.110 59.870 95.040 ;
        RECT 60.480 94.860 60.810 95.640 ;
        RECT 61.020 95.310 61.350 96.300 ;
      LAYER li1 ;
        RECT 62.040 95.790 62.470 97.370 ;
      LAYER li1 ;
        RECT 62.650 97.290 63.210 97.370 ;
        RECT 62.650 97.120 62.660 97.290 ;
        RECT 62.830 97.120 63.020 97.290 ;
        RECT 63.190 97.120 63.210 97.290 ;
        RECT 62.650 95.790 63.210 97.120 ;
        RECT 64.570 97.340 66.020 97.370 ;
        RECT 64.570 97.170 64.820 97.340 ;
        RECT 64.990 97.170 65.180 97.340 ;
        RECT 65.350 97.170 65.620 97.340 ;
        RECT 65.790 97.170 66.020 97.340 ;
        RECT 60.480 94.460 61.780 94.860 ;
        RECT 60.170 93.980 61.780 94.460 ;
      LAYER li1 ;
        RECT 62.040 94.110 62.290 95.790 ;
      LAYER li1 ;
        RECT 62.600 94.900 62.930 95.360 ;
      LAYER li1 ;
        RECT 63.390 95.080 63.720 96.870 ;
      LAYER li1 ;
        RECT 63.900 94.900 64.150 96.620 ;
        RECT 64.570 96.300 66.020 97.170 ;
        RECT 66.330 97.290 66.920 97.370 ;
        RECT 66.330 97.120 66.360 97.290 ;
        RECT 66.530 97.120 66.720 97.290 ;
        RECT 66.890 97.120 66.920 97.290 ;
        RECT 62.600 94.730 64.150 94.900 ;
        RECT 62.470 93.980 63.720 94.550 ;
        RECT 63.900 94.110 64.150 94.730 ;
        RECT 64.800 94.860 65.130 95.640 ;
        RECT 65.340 95.310 65.670 96.300 ;
        RECT 66.330 95.790 66.920 97.120 ;
      LAYER li1 ;
        RECT 67.200 95.790 67.590 97.370 ;
      LAYER li1 ;
        RECT 67.930 97.340 69.380 97.370 ;
        RECT 67.930 97.170 68.180 97.340 ;
        RECT 68.350 97.170 68.540 97.340 ;
        RECT 68.710 97.170 68.980 97.340 ;
        RECT 69.150 97.170 69.380 97.340 ;
        RECT 67.930 96.300 69.380 97.170 ;
      LAYER li1 ;
        RECT 66.370 95.160 67.080 95.550 ;
      LAYER li1 ;
        RECT 64.800 94.460 66.100 94.860 ;
        RECT 64.490 93.980 66.100 94.460 ;
        RECT 66.330 93.980 66.920 94.940 ;
      LAYER li1 ;
        RECT 67.260 94.110 67.590 95.790 ;
      LAYER li1 ;
        RECT 68.160 94.860 68.490 95.640 ;
        RECT 68.700 95.310 69.030 96.300 ;
      LAYER li1 ;
        RECT 69.720 95.790 70.150 97.370 ;
      LAYER li1 ;
        RECT 70.330 97.290 70.890 97.370 ;
        RECT 70.330 97.120 70.340 97.290 ;
        RECT 70.510 97.120 70.700 97.290 ;
        RECT 70.870 97.120 70.890 97.290 ;
        RECT 70.330 95.790 70.890 97.120 ;
        RECT 72.250 97.340 73.700 97.370 ;
        RECT 72.250 97.170 72.500 97.340 ;
        RECT 72.670 97.170 72.860 97.340 ;
        RECT 73.030 97.170 73.300 97.340 ;
        RECT 73.470 97.170 73.700 97.340 ;
        RECT 68.160 94.460 69.460 94.860 ;
        RECT 67.850 93.980 69.460 94.460 ;
      LAYER li1 ;
        RECT 69.720 94.110 69.970 95.790 ;
      LAYER li1 ;
        RECT 70.280 94.900 70.610 95.360 ;
      LAYER li1 ;
        RECT 71.070 95.080 71.400 96.870 ;
      LAYER li1 ;
        RECT 71.580 94.900 71.830 96.620 ;
        RECT 72.250 96.300 73.700 97.170 ;
        RECT 74.490 97.290 75.440 97.370 ;
        RECT 74.490 97.120 74.520 97.290 ;
        RECT 74.690 97.120 74.880 97.290 ;
        RECT 75.050 97.120 75.240 97.290 ;
        RECT 75.410 97.120 75.440 97.290 ;
        RECT 70.280 94.730 71.830 94.900 ;
        RECT 70.150 93.980 71.400 94.550 ;
        RECT 71.580 94.110 71.830 94.730 ;
        RECT 72.480 94.860 72.810 95.640 ;
        RECT 73.020 95.310 73.350 96.300 ;
        RECT 72.480 94.460 73.780 94.860 ;
      LAYER li1 ;
        RECT 74.070 94.820 74.240 96.100 ;
      LAYER li1 ;
        RECT 74.490 95.790 75.440 97.120 ;
      LAYER li1 ;
        RECT 75.970 95.720 76.440 97.370 ;
      LAYER li1 ;
        RECT 76.620 97.290 77.570 97.370 ;
        RECT 76.620 97.120 76.650 97.290 ;
        RECT 76.820 97.120 77.010 97.290 ;
        RECT 77.180 97.120 77.370 97.290 ;
        RECT 77.540 97.120 77.570 97.290 ;
        RECT 76.620 95.910 77.570 97.120 ;
        RECT 78.010 97.340 79.460 97.370 ;
        RECT 78.010 97.170 78.260 97.340 ;
        RECT 78.430 97.170 78.620 97.340 ;
        RECT 78.790 97.170 79.060 97.340 ;
        RECT 79.230 97.170 79.460 97.340 ;
        RECT 78.010 96.300 79.460 97.170 ;
        RECT 79.770 97.290 80.720 97.370 ;
        RECT 79.770 97.120 79.800 97.290 ;
        RECT 79.970 97.120 80.160 97.290 ;
        RECT 80.330 97.120 80.520 97.290 ;
        RECT 80.690 97.120 80.720 97.290 ;
      LAYER li1 ;
        RECT 75.970 95.550 76.550 95.720 ;
        RECT 74.530 95.120 75.260 95.450 ;
        RECT 75.470 95.120 76.200 95.370 ;
        RECT 76.380 95.240 76.550 95.550 ;
        RECT 76.730 95.420 77.640 95.730 ;
        RECT 76.380 95.070 77.220 95.240 ;
      LAYER li1 ;
        RECT 74.530 94.890 74.860 94.940 ;
        RECT 72.170 93.980 73.780 94.460 ;
        RECT 74.530 94.720 76.440 94.890 ;
        RECT 74.530 94.110 74.860 94.720 ;
        RECT 75.040 93.980 75.930 94.540 ;
        RECT 76.110 94.110 76.440 94.720 ;
      LAYER li1 ;
        RECT 76.890 94.110 77.220 95.070 ;
      LAYER li1 ;
        RECT 78.240 94.860 78.570 95.640 ;
        RECT 78.780 95.310 79.110 96.300 ;
        RECT 79.770 95.790 80.720 97.120 ;
      LAYER li1 ;
        RECT 80.900 95.690 81.150 97.370 ;
      LAYER li1 ;
        RECT 81.330 97.290 82.280 97.370 ;
        RECT 81.330 97.120 81.360 97.290 ;
        RECT 81.530 97.120 81.720 97.290 ;
        RECT 81.890 97.120 82.080 97.290 ;
        RECT 82.250 97.120 82.280 97.290 ;
        RECT 81.330 95.870 82.280 97.120 ;
      LAYER li1 ;
        RECT 82.460 95.690 82.790 97.370 ;
      LAYER li1 ;
        RECT 82.970 97.290 83.920 97.370 ;
        RECT 82.970 97.120 83.000 97.290 ;
        RECT 83.170 97.120 83.360 97.290 ;
        RECT 83.530 97.120 83.720 97.290 ;
        RECT 83.890 97.120 83.920 97.290 ;
        RECT 82.970 95.910 83.920 97.120 ;
      LAYER li1 ;
        RECT 80.900 95.520 82.790 95.690 ;
        RECT 80.900 95.390 81.070 95.520 ;
        RECT 83.570 95.390 83.900 95.730 ;
        RECT 79.810 95.160 81.070 95.390 ;
      LAYER li1 ;
        RECT 81.250 95.210 83.280 95.340 ;
        RECT 84.100 95.210 84.350 97.370 ;
        RECT 84.730 97.340 86.180 97.370 ;
        RECT 84.730 97.170 84.980 97.340 ;
        RECT 85.150 97.170 85.340 97.340 ;
        RECT 85.510 97.170 85.780 97.340 ;
        RECT 85.950 97.170 86.180 97.340 ;
        RECT 84.730 96.300 86.180 97.170 ;
        RECT 86.490 97.290 87.440 97.370 ;
        RECT 86.490 97.120 86.520 97.290 ;
        RECT 86.690 97.120 86.880 97.290 ;
        RECT 87.050 97.120 87.240 97.290 ;
        RECT 87.410 97.120 87.440 97.290 ;
        RECT 81.250 95.170 84.350 95.210 ;
      LAYER li1 ;
        RECT 80.900 94.990 81.070 95.160 ;
      LAYER li1 ;
        RECT 83.110 95.040 84.350 95.170 ;
        RECT 78.240 94.460 79.540 94.860 ;
        RECT 77.930 93.980 79.540 94.460 ;
        RECT 79.770 93.980 80.720 94.940 ;
      LAYER li1 ;
        RECT 80.900 94.820 82.710 94.990 ;
        RECT 80.900 94.110 81.150 94.820 ;
      LAYER li1 ;
        RECT 81.330 93.980 82.280 94.640 ;
      LAYER li1 ;
        RECT 82.460 94.110 82.710 94.820 ;
      LAYER li1 ;
        RECT 82.890 93.980 83.840 94.860 ;
        RECT 84.020 94.110 84.350 95.040 ;
        RECT 84.960 94.860 85.290 95.640 ;
        RECT 85.500 95.310 85.830 96.300 ;
        RECT 86.490 95.790 87.440 97.120 ;
      LAYER li1 ;
        RECT 87.620 95.690 87.870 97.370 ;
      LAYER li1 ;
        RECT 88.050 97.290 89.000 97.370 ;
        RECT 88.050 97.120 88.080 97.290 ;
        RECT 88.250 97.120 88.440 97.290 ;
        RECT 88.610 97.120 88.800 97.290 ;
        RECT 88.970 97.120 89.000 97.290 ;
        RECT 88.050 95.870 89.000 97.120 ;
      LAYER li1 ;
        RECT 89.180 95.690 89.510 97.370 ;
      LAYER li1 ;
        RECT 89.690 97.290 90.640 97.370 ;
        RECT 89.690 97.120 89.720 97.290 ;
        RECT 89.890 97.120 90.080 97.290 ;
        RECT 90.250 97.120 90.440 97.290 ;
        RECT 90.610 97.120 90.640 97.290 ;
        RECT 89.690 95.910 90.640 97.120 ;
      LAYER li1 ;
        RECT 87.620 95.520 89.510 95.690 ;
        RECT 87.620 95.390 87.790 95.520 ;
        RECT 90.290 95.390 90.620 95.730 ;
        RECT 86.530 95.160 87.790 95.390 ;
      LAYER li1 ;
        RECT 87.970 95.210 90.000 95.340 ;
        RECT 90.820 95.210 91.070 97.370 ;
        RECT 91.450 97.340 92.900 97.370 ;
        RECT 91.450 97.170 91.700 97.340 ;
        RECT 91.870 97.170 92.060 97.340 ;
        RECT 92.230 97.170 92.500 97.340 ;
        RECT 92.670 97.170 92.900 97.340 ;
        RECT 91.450 96.300 92.900 97.170 ;
        RECT 93.210 97.290 94.880 97.370 ;
        RECT 93.210 97.120 93.240 97.290 ;
        RECT 93.410 97.120 93.600 97.290 ;
        RECT 93.770 97.120 93.960 97.290 ;
        RECT 94.130 97.120 94.320 97.290 ;
        RECT 94.490 97.120 94.680 97.290 ;
        RECT 94.850 97.120 94.880 97.290 ;
        RECT 87.970 95.170 91.070 95.210 ;
      LAYER li1 ;
        RECT 87.620 94.990 87.790 95.160 ;
      LAYER li1 ;
        RECT 89.830 95.040 91.070 95.170 ;
        RECT 84.960 94.460 86.260 94.860 ;
        RECT 84.650 93.980 86.260 94.460 ;
        RECT 86.490 93.980 87.440 94.940 ;
      LAYER li1 ;
        RECT 87.620 94.820 89.430 94.990 ;
        RECT 87.620 94.110 87.870 94.820 ;
      LAYER li1 ;
        RECT 88.050 93.980 89.000 94.640 ;
      LAYER li1 ;
        RECT 89.180 94.110 89.430 94.820 ;
      LAYER li1 ;
        RECT 89.610 93.980 90.560 94.860 ;
        RECT 90.740 94.110 91.070 95.040 ;
        RECT 91.680 94.860 92.010 95.640 ;
        RECT 92.220 95.310 92.550 96.300 ;
        RECT 93.210 95.910 94.880 97.120 ;
      LAYER li1 ;
        RECT 93.250 95.140 93.550 95.730 ;
        RECT 93.730 95.390 94.920 95.730 ;
        RECT 95.100 95.390 95.430 96.870 ;
        RECT 95.610 95.210 95.880 97.370 ;
      LAYER li1 ;
        RECT 96.730 97.340 98.180 97.370 ;
        RECT 96.730 97.170 96.980 97.340 ;
        RECT 97.150 97.170 97.340 97.340 ;
        RECT 97.510 97.170 97.780 97.340 ;
        RECT 97.950 97.170 98.180 97.340 ;
        RECT 96.730 96.300 98.180 97.170 ;
        RECT 98.970 97.290 99.920 97.370 ;
        RECT 98.970 97.120 99.000 97.290 ;
        RECT 99.170 97.120 99.360 97.290 ;
        RECT 99.530 97.120 99.720 97.290 ;
        RECT 99.890 97.120 99.920 97.290 ;
      LAYER li1 ;
        RECT 94.050 95.040 95.880 95.210 ;
      LAYER li1 ;
        RECT 91.680 94.460 92.980 94.860 ;
        RECT 91.370 93.980 92.980 94.460 ;
        RECT 93.210 93.980 93.800 94.940 ;
      LAYER li1 ;
        RECT 94.050 94.110 94.300 95.040 ;
      LAYER li1 ;
        RECT 94.480 93.980 95.430 94.860 ;
      LAYER li1 ;
        RECT 95.610 94.110 95.880 95.040 ;
      LAYER li1 ;
        RECT 96.960 94.860 97.290 95.640 ;
        RECT 97.500 95.310 97.830 96.300 ;
        RECT 98.970 95.790 99.920 97.120 ;
      LAYER li1 ;
        RECT 100.100 95.690 100.350 97.370 ;
      LAYER li1 ;
        RECT 100.530 97.290 101.480 97.370 ;
        RECT 100.530 97.120 100.560 97.290 ;
        RECT 100.730 97.120 100.920 97.290 ;
        RECT 101.090 97.120 101.280 97.290 ;
        RECT 101.450 97.120 101.480 97.290 ;
        RECT 100.530 95.870 101.480 97.120 ;
      LAYER li1 ;
        RECT 101.660 95.690 101.990 97.370 ;
      LAYER li1 ;
        RECT 102.170 97.290 103.120 97.370 ;
        RECT 102.170 97.120 102.200 97.290 ;
        RECT 102.370 97.120 102.560 97.290 ;
        RECT 102.730 97.120 102.920 97.290 ;
        RECT 103.090 97.120 103.120 97.290 ;
        RECT 102.170 95.910 103.120 97.120 ;
      LAYER li1 ;
        RECT 100.100 95.520 101.990 95.690 ;
        RECT 100.100 95.390 100.270 95.520 ;
        RECT 102.770 95.390 103.100 95.730 ;
        RECT 99.010 95.160 100.270 95.390 ;
      LAYER li1 ;
        RECT 100.450 95.210 102.480 95.340 ;
        RECT 103.300 95.210 103.550 97.370 ;
        RECT 103.930 97.340 105.380 97.370 ;
        RECT 103.930 97.170 104.180 97.340 ;
        RECT 104.350 97.170 104.540 97.340 ;
        RECT 104.710 97.170 104.980 97.340 ;
        RECT 105.150 97.170 105.380 97.340 ;
        RECT 103.930 96.300 105.380 97.170 ;
        RECT 105.690 97.290 106.640 97.370 ;
        RECT 105.690 97.120 105.720 97.290 ;
        RECT 105.890 97.120 106.080 97.290 ;
        RECT 106.250 97.120 106.440 97.290 ;
        RECT 106.610 97.120 106.640 97.290 ;
        RECT 100.450 95.170 103.550 95.210 ;
      LAYER li1 ;
        RECT 100.100 94.990 100.270 95.160 ;
      LAYER li1 ;
        RECT 102.310 95.040 103.550 95.170 ;
        RECT 96.960 94.460 98.260 94.860 ;
        RECT 96.650 93.980 98.260 94.460 ;
        RECT 98.970 93.980 99.920 94.940 ;
      LAYER li1 ;
        RECT 100.100 94.820 101.910 94.990 ;
        RECT 100.100 94.110 100.350 94.820 ;
      LAYER li1 ;
        RECT 100.530 93.980 101.480 94.640 ;
      LAYER li1 ;
        RECT 101.660 94.110 101.910 94.820 ;
      LAYER li1 ;
        RECT 102.090 93.980 103.040 94.860 ;
        RECT 103.220 94.110 103.550 95.040 ;
        RECT 104.160 94.860 104.490 95.640 ;
        RECT 104.700 95.310 105.030 96.300 ;
        RECT 105.690 95.790 106.640 97.120 ;
      LAYER li1 ;
        RECT 106.820 95.690 107.070 97.370 ;
      LAYER li1 ;
        RECT 107.250 97.290 108.200 97.370 ;
        RECT 107.250 97.120 107.280 97.290 ;
        RECT 107.450 97.120 107.640 97.290 ;
        RECT 107.810 97.120 108.000 97.290 ;
        RECT 108.170 97.120 108.200 97.290 ;
        RECT 107.250 95.870 108.200 97.120 ;
      LAYER li1 ;
        RECT 108.380 95.690 108.710 97.370 ;
      LAYER li1 ;
        RECT 108.890 97.290 109.840 97.370 ;
        RECT 108.890 97.120 108.920 97.290 ;
        RECT 109.090 97.120 109.280 97.290 ;
        RECT 109.450 97.120 109.640 97.290 ;
        RECT 109.810 97.120 109.840 97.290 ;
        RECT 108.890 95.910 109.840 97.120 ;
      LAYER li1 ;
        RECT 106.820 95.520 108.710 95.690 ;
        RECT 106.820 95.390 106.990 95.520 ;
        RECT 109.490 95.390 109.820 95.730 ;
        RECT 105.730 95.160 106.990 95.390 ;
      LAYER li1 ;
        RECT 107.170 95.210 109.200 95.340 ;
        RECT 110.020 95.210 110.270 97.370 ;
        RECT 110.650 97.340 112.100 97.370 ;
        RECT 110.650 97.170 110.900 97.340 ;
        RECT 111.070 97.170 111.260 97.340 ;
        RECT 111.430 97.170 111.700 97.340 ;
        RECT 111.870 97.170 112.100 97.340 ;
        RECT 110.650 96.300 112.100 97.170 ;
        RECT 112.410 97.290 114.080 97.370 ;
        RECT 112.410 97.120 112.440 97.290 ;
        RECT 112.610 97.120 112.800 97.290 ;
        RECT 112.970 97.120 113.160 97.290 ;
        RECT 113.330 97.120 113.520 97.290 ;
        RECT 113.690 97.120 113.880 97.290 ;
        RECT 114.050 97.120 114.080 97.290 ;
        RECT 107.170 95.170 110.270 95.210 ;
      LAYER li1 ;
        RECT 106.820 94.990 106.990 95.160 ;
      LAYER li1 ;
        RECT 109.030 95.040 110.270 95.170 ;
        RECT 104.160 94.460 105.460 94.860 ;
        RECT 103.850 93.980 105.460 94.460 ;
        RECT 105.690 93.980 106.640 94.940 ;
      LAYER li1 ;
        RECT 106.820 94.820 108.630 94.990 ;
        RECT 106.820 94.110 107.070 94.820 ;
      LAYER li1 ;
        RECT 107.250 93.980 108.200 94.640 ;
      LAYER li1 ;
        RECT 108.380 94.110 108.630 94.820 ;
      LAYER li1 ;
        RECT 108.810 93.980 109.760 94.860 ;
        RECT 109.940 94.110 110.270 95.040 ;
        RECT 110.880 94.860 111.210 95.640 ;
        RECT 111.420 95.310 111.750 96.300 ;
        RECT 112.410 95.910 114.080 97.120 ;
      LAYER li1 ;
        RECT 112.450 95.390 113.640 95.730 ;
        RECT 113.820 95.390 114.150 95.730 ;
        RECT 114.340 95.210 114.600 97.370 ;
      LAYER li1 ;
        RECT 114.970 97.340 116.420 97.370 ;
        RECT 114.970 97.170 115.220 97.340 ;
        RECT 115.390 97.170 115.580 97.340 ;
        RECT 115.750 97.170 116.020 97.340 ;
        RECT 116.190 97.170 116.420 97.340 ;
        RECT 114.970 96.300 116.420 97.170 ;
      LAYER li1 ;
        RECT 113.520 95.040 114.600 95.210 ;
      LAYER li1 ;
        RECT 110.880 94.460 112.180 94.860 ;
        RECT 110.570 93.980 112.180 94.460 ;
        RECT 112.410 93.980 113.340 94.940 ;
      LAYER li1 ;
        RECT 113.520 94.110 113.850 95.040 ;
      LAYER li1 ;
        RECT 115.200 94.860 115.530 95.640 ;
        RECT 115.740 95.310 116.070 96.300 ;
      LAYER li1 ;
        RECT 116.760 95.790 117.190 97.370 ;
      LAYER li1 ;
        RECT 117.370 97.290 117.930 97.370 ;
        RECT 117.370 97.120 117.380 97.290 ;
        RECT 117.550 97.120 117.740 97.290 ;
        RECT 117.910 97.120 117.930 97.290 ;
        RECT 117.370 95.790 117.930 97.120 ;
        RECT 119.290 97.340 120.740 97.370 ;
        RECT 119.290 97.170 119.540 97.340 ;
        RECT 119.710 97.170 119.900 97.340 ;
        RECT 120.070 97.170 120.340 97.340 ;
        RECT 120.510 97.170 120.740 97.340 ;
        RECT 114.040 93.980 114.630 94.860 ;
        RECT 115.200 94.460 116.500 94.860 ;
        RECT 114.890 93.980 116.500 94.460 ;
      LAYER li1 ;
        RECT 116.760 94.110 117.010 95.790 ;
      LAYER li1 ;
        RECT 117.320 94.900 117.650 95.360 ;
      LAYER li1 ;
        RECT 118.110 95.080 118.440 96.870 ;
      LAYER li1 ;
        RECT 118.620 94.900 118.870 96.620 ;
        RECT 119.290 96.300 120.740 97.170 ;
        RECT 121.530 97.290 122.480 97.370 ;
        RECT 121.530 97.120 121.560 97.290 ;
        RECT 121.730 97.120 121.920 97.290 ;
        RECT 122.090 97.120 122.280 97.290 ;
        RECT 122.450 97.120 122.480 97.290 ;
        RECT 117.320 94.730 118.870 94.900 ;
        RECT 117.190 93.980 118.440 94.550 ;
        RECT 118.620 94.110 118.870 94.730 ;
        RECT 119.520 94.860 119.850 95.640 ;
        RECT 120.060 95.310 120.390 96.300 ;
        RECT 121.530 95.790 122.480 97.120 ;
      LAYER li1 ;
        RECT 122.660 95.690 122.910 97.370 ;
      LAYER li1 ;
        RECT 123.090 97.290 124.040 97.370 ;
        RECT 123.090 97.120 123.120 97.290 ;
        RECT 123.290 97.120 123.480 97.290 ;
        RECT 123.650 97.120 123.840 97.290 ;
        RECT 124.010 97.120 124.040 97.290 ;
        RECT 123.090 95.870 124.040 97.120 ;
      LAYER li1 ;
        RECT 124.220 95.690 124.550 97.370 ;
      LAYER li1 ;
        RECT 124.730 97.290 125.680 97.370 ;
        RECT 124.730 97.120 124.760 97.290 ;
        RECT 124.930 97.120 125.120 97.290 ;
        RECT 125.290 97.120 125.480 97.290 ;
        RECT 125.650 97.120 125.680 97.290 ;
        RECT 124.730 95.910 125.680 97.120 ;
      LAYER li1 ;
        RECT 122.660 95.520 124.550 95.690 ;
        RECT 122.660 95.390 122.830 95.520 ;
        RECT 125.330 95.390 125.660 95.730 ;
        RECT 121.570 95.160 122.830 95.390 ;
      LAYER li1 ;
        RECT 123.010 95.210 125.040 95.340 ;
        RECT 125.860 95.210 126.110 97.370 ;
        RECT 126.490 97.340 127.940 97.370 ;
        RECT 126.490 97.170 126.740 97.340 ;
        RECT 126.910 97.170 127.100 97.340 ;
        RECT 127.270 97.170 127.540 97.340 ;
        RECT 127.710 97.170 127.940 97.340 ;
        RECT 126.490 96.300 127.940 97.170 ;
        RECT 128.890 97.290 129.450 97.370 ;
        RECT 128.890 97.120 128.900 97.290 ;
        RECT 129.070 97.120 129.260 97.290 ;
        RECT 129.430 97.120 129.450 97.290 ;
        RECT 123.010 95.170 126.110 95.210 ;
      LAYER li1 ;
        RECT 122.660 94.990 122.830 95.160 ;
      LAYER li1 ;
        RECT 124.870 95.040 126.110 95.170 ;
        RECT 119.520 94.460 120.820 94.860 ;
        RECT 119.210 93.980 120.820 94.460 ;
        RECT 121.530 93.980 122.480 94.940 ;
      LAYER li1 ;
        RECT 122.660 94.820 124.470 94.990 ;
        RECT 122.660 94.110 122.910 94.820 ;
      LAYER li1 ;
        RECT 123.090 93.980 124.040 94.640 ;
      LAYER li1 ;
        RECT 124.220 94.110 124.470 94.820 ;
      LAYER li1 ;
        RECT 124.650 93.980 125.600 94.860 ;
        RECT 125.780 94.110 126.110 95.040 ;
        RECT 126.720 94.860 127.050 95.640 ;
        RECT 127.260 95.310 127.590 96.300 ;
        RECT 128.890 95.790 129.450 97.120 ;
        RECT 131.060 97.340 133.800 97.360 ;
        RECT 131.060 97.170 131.270 97.340 ;
        RECT 131.440 97.170 131.710 97.340 ;
        RECT 131.880 97.170 132.120 97.340 ;
        RECT 132.290 97.170 132.550 97.340 ;
        RECT 132.720 97.170 132.990 97.340 ;
        RECT 133.160 97.170 133.400 97.340 ;
        RECT 133.570 97.170 133.800 97.340 ;
        RECT 128.840 94.900 129.170 95.360 ;
        RECT 130.140 94.900 130.390 96.620 ;
        RECT 131.060 96.290 133.800 97.170 ;
        RECT 134.900 97.340 137.640 97.360 ;
        RECT 134.900 97.170 135.110 97.340 ;
        RECT 135.280 97.170 135.550 97.340 ;
        RECT 135.720 97.170 135.960 97.340 ;
        RECT 136.130 97.170 136.390 97.340 ;
        RECT 136.560 97.170 136.830 97.340 ;
        RECT 137.000 97.170 137.240 97.340 ;
        RECT 137.410 97.170 137.640 97.340 ;
        RECT 134.900 96.290 137.640 97.170 ;
        RECT 138.740 97.340 141.480 97.360 ;
        RECT 138.740 97.170 138.950 97.340 ;
        RECT 139.120 97.170 139.390 97.340 ;
        RECT 139.560 97.170 139.800 97.340 ;
        RECT 139.970 97.170 140.230 97.340 ;
        RECT 140.400 97.170 140.670 97.340 ;
        RECT 140.840 97.170 141.080 97.340 ;
        RECT 141.250 97.170 141.480 97.340 ;
        RECT 138.740 96.290 141.480 97.170 ;
        RECT 131.300 94.970 131.630 95.640 ;
        RECT 132.030 95.310 132.360 96.290 ;
        RECT 132.580 94.970 132.910 95.640 ;
        RECT 133.310 95.310 133.640 96.290 ;
        RECT 135.140 94.970 135.470 95.640 ;
        RECT 135.870 95.310 136.200 96.290 ;
        RECT 136.420 94.970 136.750 95.640 ;
        RECT 137.150 95.310 137.480 96.290 ;
        RECT 138.980 94.970 139.310 95.640 ;
        RECT 139.710 95.310 140.040 96.290 ;
        RECT 140.260 94.970 140.590 95.640 ;
        RECT 140.990 95.310 141.320 96.290 ;
        RECT 126.720 94.460 128.020 94.860 ;
        RECT 128.840 94.730 130.390 94.900 ;
        RECT 126.410 93.980 128.020 94.460 ;
        RECT 128.710 93.980 129.960 94.550 ;
        RECT 130.140 94.110 130.390 94.730 ;
        RECT 131.140 93.970 133.870 94.970 ;
        RECT 134.980 93.970 137.710 94.970 ;
        RECT 138.820 93.970 141.550 94.970 ;
        RECT 5.760 93.520 5.920 93.700 ;
        RECT 6.090 93.520 6.400 93.700 ;
        RECT 6.570 93.520 6.880 93.700 ;
        RECT 7.050 93.520 7.360 93.700 ;
        RECT 7.530 93.520 7.840 93.700 ;
        RECT 8.010 93.520 8.320 93.700 ;
        RECT 8.490 93.520 8.800 93.700 ;
        RECT 8.970 93.520 9.280 93.700 ;
        RECT 9.450 93.520 9.760 93.700 ;
        RECT 9.930 93.520 10.240 93.700 ;
        RECT 10.410 93.520 10.720 93.700 ;
        RECT 10.890 93.520 11.200 93.700 ;
        RECT 11.370 93.520 11.680 93.700 ;
        RECT 11.850 93.520 12.160 93.700 ;
        RECT 12.330 93.520 12.640 93.700 ;
        RECT 12.810 93.520 13.120 93.700 ;
        RECT 13.290 93.520 13.600 93.700 ;
        RECT 13.770 93.520 14.080 93.700 ;
        RECT 14.250 93.520 14.560 93.700 ;
        RECT 14.730 93.520 15.040 93.700 ;
        RECT 15.210 93.520 15.520 93.700 ;
        RECT 15.690 93.520 16.000 93.700 ;
        RECT 16.170 93.520 16.480 93.700 ;
        RECT 16.650 93.520 16.960 93.700 ;
        RECT 17.130 93.520 17.440 93.700 ;
        RECT 17.610 93.520 17.920 93.700 ;
        RECT 18.090 93.520 18.400 93.700 ;
        RECT 18.570 93.520 18.880 93.700 ;
        RECT 19.050 93.520 19.360 93.700 ;
        RECT 19.530 93.520 19.840 93.700 ;
        RECT 20.010 93.520 20.320 93.700 ;
        RECT 20.490 93.520 20.800 93.700 ;
        RECT 20.970 93.520 21.280 93.700 ;
        RECT 21.450 93.520 21.760 93.700 ;
        RECT 21.930 93.520 22.240 93.700 ;
        RECT 22.410 93.520 22.720 93.700 ;
        RECT 22.890 93.520 23.200 93.700 ;
        RECT 23.370 93.520 23.680 93.700 ;
        RECT 23.850 93.520 24.160 93.700 ;
        RECT 24.330 93.520 24.640 93.700 ;
        RECT 24.810 93.520 25.120 93.700 ;
        RECT 25.290 93.520 25.600 93.700 ;
        RECT 25.770 93.520 26.080 93.700 ;
        RECT 26.250 93.520 26.560 93.700 ;
        RECT 26.730 93.520 27.040 93.700 ;
        RECT 27.210 93.520 27.520 93.700 ;
        RECT 27.690 93.520 28.000 93.700 ;
        RECT 28.170 93.520 28.480 93.700 ;
        RECT 28.650 93.520 28.960 93.700 ;
        RECT 29.130 93.520 29.440 93.700 ;
        RECT 29.610 93.520 29.920 93.700 ;
        RECT 30.090 93.520 30.400 93.700 ;
        RECT 30.570 93.520 30.880 93.700 ;
        RECT 31.050 93.520 31.360 93.700 ;
        RECT 31.530 93.520 31.840 93.700 ;
        RECT 32.010 93.520 32.320 93.700 ;
        RECT 32.490 93.520 32.640 93.700 ;
        RECT 33.120 93.520 33.280 93.700 ;
        RECT 33.450 93.520 33.760 93.700 ;
        RECT 33.930 93.520 34.240 93.700 ;
        RECT 34.410 93.520 34.720 93.700 ;
        RECT 34.890 93.520 35.200 93.700 ;
        RECT 35.370 93.520 35.680 93.700 ;
        RECT 35.850 93.520 36.160 93.700 ;
        RECT 36.330 93.520 36.640 93.700 ;
        RECT 36.810 93.520 37.120 93.700 ;
        RECT 37.290 93.520 37.600 93.700 ;
        RECT 37.770 93.520 38.080 93.700 ;
        RECT 38.250 93.520 38.560 93.700 ;
        RECT 38.730 93.520 39.040 93.700 ;
        RECT 39.210 93.520 39.520 93.700 ;
        RECT 39.690 93.520 40.000 93.700 ;
        RECT 40.170 93.520 40.480 93.700 ;
        RECT 40.650 93.520 40.960 93.700 ;
        RECT 41.130 93.520 41.440 93.700 ;
        RECT 41.610 93.520 41.920 93.700 ;
        RECT 42.090 93.520 42.400 93.700 ;
        RECT 42.570 93.520 42.880 93.700 ;
        RECT 43.050 93.520 43.360 93.700 ;
        RECT 43.530 93.520 43.840 93.700 ;
        RECT 44.010 93.520 44.320 93.700 ;
        RECT 44.490 93.520 44.800 93.700 ;
        RECT 44.970 93.520 45.280 93.700 ;
        RECT 45.450 93.520 45.760 93.700 ;
        RECT 45.930 93.520 46.240 93.700 ;
        RECT 46.410 93.520 46.720 93.700 ;
        RECT 46.890 93.520 47.200 93.700 ;
        RECT 47.370 93.520 47.680 93.700 ;
        RECT 47.850 93.520 48.160 93.700 ;
        RECT 48.330 93.520 48.640 93.700 ;
        RECT 48.810 93.520 49.120 93.700 ;
        RECT 49.290 93.520 49.600 93.700 ;
        RECT 49.770 93.520 50.080 93.700 ;
        RECT 50.250 93.520 50.560 93.700 ;
        RECT 50.730 93.520 51.040 93.700 ;
        RECT 51.210 93.520 51.520 93.700 ;
        RECT 51.690 93.520 52.000 93.700 ;
        RECT 52.170 93.520 52.480 93.700 ;
        RECT 52.650 93.520 52.960 93.700 ;
        RECT 53.130 93.520 53.440 93.700 ;
        RECT 53.610 93.520 53.920 93.700 ;
        RECT 54.090 93.520 54.400 93.700 ;
        RECT 54.570 93.520 54.880 93.700 ;
        RECT 55.050 93.520 55.360 93.700 ;
        RECT 55.530 93.520 55.840 93.700 ;
        RECT 56.010 93.520 56.320 93.700 ;
        RECT 56.490 93.520 56.800 93.700 ;
        RECT 56.970 93.520 57.280 93.700 ;
        RECT 57.450 93.520 57.760 93.700 ;
        RECT 57.930 93.520 58.240 93.700 ;
        RECT 58.410 93.520 58.720 93.700 ;
        RECT 58.890 93.520 59.200 93.700 ;
        RECT 59.370 93.520 59.680 93.700 ;
        RECT 59.850 93.520 60.160 93.700 ;
        RECT 60.330 93.520 60.640 93.700 ;
        RECT 60.810 93.520 61.120 93.700 ;
        RECT 61.290 93.520 61.600 93.700 ;
        RECT 61.770 93.520 62.080 93.700 ;
        RECT 62.250 93.520 62.560 93.700 ;
        RECT 62.730 93.520 63.040 93.700 ;
        RECT 63.210 93.520 63.520 93.700 ;
        RECT 63.690 93.520 64.000 93.700 ;
        RECT 64.170 93.520 64.480 93.700 ;
        RECT 64.650 93.520 64.960 93.700 ;
        RECT 65.130 93.520 65.440 93.700 ;
        RECT 65.610 93.520 65.920 93.700 ;
        RECT 66.090 93.520 66.400 93.700 ;
        RECT 66.570 93.520 66.880 93.700 ;
        RECT 67.050 93.520 67.360 93.700 ;
        RECT 67.530 93.520 67.840 93.700 ;
        RECT 68.010 93.520 68.320 93.700 ;
        RECT 68.490 93.520 68.800 93.700 ;
        RECT 68.970 93.520 69.280 93.700 ;
        RECT 69.450 93.520 69.760 93.700 ;
        RECT 69.930 93.520 70.240 93.700 ;
        RECT 70.410 93.520 70.720 93.700 ;
        RECT 70.890 93.520 71.200 93.700 ;
        RECT 71.370 93.520 71.680 93.700 ;
        RECT 71.850 93.520 72.160 93.700 ;
        RECT 72.330 93.520 72.640 93.700 ;
        RECT 72.810 93.520 73.120 93.700 ;
        RECT 73.290 93.520 73.600 93.700 ;
        RECT 73.770 93.520 73.920 93.700 ;
        RECT 74.400 93.520 74.560 93.700 ;
        RECT 74.730 93.520 75.040 93.700 ;
        RECT 75.210 93.520 75.520 93.700 ;
        RECT 75.690 93.520 76.000 93.700 ;
        RECT 76.170 93.520 76.480 93.700 ;
        RECT 76.650 93.520 76.960 93.700 ;
        RECT 77.130 93.520 77.440 93.700 ;
        RECT 77.610 93.520 77.920 93.700 ;
        RECT 78.090 93.520 78.400 93.700 ;
        RECT 78.570 93.520 78.880 93.700 ;
        RECT 79.050 93.520 79.360 93.700 ;
        RECT 79.530 93.520 79.840 93.700 ;
        RECT 80.010 93.520 80.320 93.700 ;
        RECT 80.490 93.520 80.800 93.700 ;
        RECT 80.970 93.520 81.280 93.700 ;
        RECT 81.450 93.520 81.760 93.700 ;
        RECT 81.930 93.520 82.240 93.700 ;
        RECT 82.410 93.520 82.720 93.700 ;
        RECT 82.890 93.520 83.200 93.700 ;
        RECT 83.370 93.520 83.680 93.700 ;
        RECT 83.850 93.520 84.160 93.700 ;
        RECT 84.330 93.520 84.640 93.700 ;
        RECT 84.810 93.520 85.120 93.700 ;
        RECT 85.290 93.520 85.600 93.700 ;
        RECT 85.770 93.520 86.080 93.700 ;
        RECT 86.250 93.520 86.560 93.700 ;
        RECT 86.730 93.520 87.040 93.700 ;
        RECT 87.210 93.520 87.520 93.700 ;
        RECT 87.690 93.520 88.000 93.700 ;
        RECT 88.170 93.520 88.480 93.700 ;
        RECT 88.650 93.520 88.960 93.700 ;
        RECT 89.130 93.520 89.440 93.700 ;
        RECT 89.610 93.520 89.920 93.700 ;
        RECT 90.090 93.520 90.400 93.700 ;
        RECT 90.570 93.520 90.880 93.700 ;
        RECT 91.050 93.520 91.360 93.700 ;
        RECT 91.530 93.520 91.840 93.700 ;
        RECT 92.010 93.520 92.320 93.700 ;
        RECT 92.490 93.520 92.800 93.700 ;
        RECT 92.970 93.520 93.280 93.700 ;
        RECT 93.450 93.520 93.760 93.700 ;
        RECT 93.930 93.520 94.240 93.700 ;
        RECT 94.410 93.520 94.720 93.700 ;
        RECT 94.890 93.520 95.200 93.700 ;
        RECT 95.370 93.520 95.680 93.700 ;
        RECT 95.850 93.520 96.160 93.700 ;
        RECT 96.330 93.520 96.640 93.700 ;
        RECT 96.810 93.520 97.120 93.700 ;
        RECT 97.290 93.520 97.600 93.700 ;
        RECT 97.770 93.520 98.080 93.700 ;
        RECT 98.250 93.520 98.400 93.700 ;
        RECT 98.880 93.520 99.040 93.700 ;
        RECT 99.210 93.520 99.520 93.700 ;
        RECT 99.690 93.520 100.000 93.700 ;
        RECT 100.170 93.520 100.480 93.700 ;
        RECT 100.650 93.520 100.960 93.700 ;
        RECT 101.130 93.520 101.440 93.700 ;
        RECT 101.610 93.520 101.920 93.700 ;
        RECT 102.090 93.520 102.400 93.700 ;
        RECT 102.570 93.520 102.880 93.700 ;
        RECT 103.050 93.520 103.360 93.700 ;
        RECT 103.530 93.520 103.840 93.700 ;
        RECT 104.010 93.520 104.320 93.700 ;
        RECT 104.490 93.520 104.800 93.700 ;
        RECT 104.970 93.520 105.280 93.700 ;
        RECT 105.450 93.520 105.760 93.700 ;
        RECT 105.930 93.520 106.240 93.700 ;
        RECT 106.410 93.520 106.720 93.700 ;
        RECT 106.890 93.520 107.200 93.700 ;
        RECT 107.370 93.520 107.680 93.700 ;
        RECT 107.850 93.520 108.160 93.700 ;
        RECT 108.330 93.520 108.640 93.700 ;
        RECT 108.810 93.520 109.120 93.700 ;
        RECT 109.290 93.520 109.600 93.700 ;
        RECT 109.770 93.520 110.080 93.700 ;
        RECT 110.250 93.520 110.560 93.700 ;
        RECT 110.730 93.520 111.040 93.700 ;
        RECT 111.210 93.520 111.520 93.700 ;
        RECT 111.690 93.520 112.000 93.700 ;
        RECT 112.170 93.520 112.480 93.700 ;
        RECT 112.650 93.520 112.960 93.700 ;
        RECT 113.130 93.520 113.440 93.700 ;
        RECT 113.610 93.520 113.920 93.700 ;
        RECT 114.090 93.520 114.400 93.700 ;
        RECT 114.570 93.520 114.880 93.700 ;
        RECT 115.050 93.520 115.360 93.700 ;
        RECT 115.530 93.520 115.840 93.700 ;
        RECT 116.010 93.520 116.320 93.700 ;
        RECT 116.490 93.520 116.800 93.700 ;
        RECT 116.970 93.520 117.280 93.700 ;
        RECT 117.450 93.520 117.760 93.700 ;
        RECT 117.930 93.520 118.240 93.700 ;
        RECT 118.410 93.520 118.720 93.700 ;
        RECT 118.890 93.520 119.200 93.700 ;
        RECT 119.370 93.520 119.680 93.700 ;
        RECT 119.850 93.520 120.160 93.700 ;
        RECT 120.330 93.520 120.640 93.700 ;
        RECT 120.810 93.520 120.960 93.700 ;
        RECT 121.440 93.520 121.600 93.700 ;
        RECT 121.770 93.520 122.080 93.700 ;
        RECT 122.250 93.520 122.560 93.700 ;
        RECT 122.730 93.520 123.040 93.700 ;
        RECT 123.210 93.520 123.520 93.700 ;
        RECT 123.690 93.520 124.000 93.700 ;
        RECT 124.170 93.520 124.480 93.700 ;
        RECT 124.650 93.520 124.960 93.700 ;
        RECT 125.130 93.520 125.440 93.700 ;
        RECT 125.610 93.520 125.920 93.700 ;
        RECT 126.090 93.520 126.400 93.700 ;
        RECT 126.570 93.520 126.880 93.700 ;
        RECT 127.050 93.520 127.360 93.700 ;
        RECT 127.530 93.520 127.840 93.700 ;
        RECT 128.010 93.520 128.320 93.700 ;
        RECT 128.490 93.520 128.800 93.700 ;
        RECT 128.970 93.520 129.280 93.700 ;
        RECT 129.450 93.520 129.760 93.700 ;
        RECT 129.930 93.520 130.240 93.700 ;
        RECT 130.410 93.520 130.720 93.700 ;
        RECT 130.890 93.520 131.200 93.700 ;
        RECT 131.370 93.520 131.680 93.700 ;
        RECT 131.850 93.520 132.160 93.700 ;
        RECT 132.330 93.520 132.640 93.700 ;
        RECT 132.810 93.520 133.120 93.700 ;
        RECT 133.290 93.520 133.600 93.700 ;
        RECT 133.770 93.520 134.080 93.700 ;
        RECT 134.250 93.520 134.560 93.700 ;
        RECT 134.730 93.520 135.040 93.700 ;
        RECT 135.210 93.520 135.520 93.700 ;
        RECT 135.690 93.520 136.000 93.700 ;
        RECT 136.170 93.520 136.480 93.700 ;
        RECT 136.650 93.520 136.960 93.700 ;
        RECT 137.130 93.520 137.440 93.700 ;
        RECT 137.610 93.520 137.920 93.700 ;
        RECT 138.090 93.520 138.400 93.700 ;
        RECT 138.570 93.520 138.880 93.700 ;
        RECT 139.050 93.520 139.360 93.700 ;
        RECT 139.530 93.520 139.840 93.700 ;
        RECT 140.010 93.520 140.320 93.700 ;
        RECT 140.490 93.520 140.800 93.700 ;
        RECT 140.970 93.520 141.280 93.700 ;
        RECT 141.450 93.520 141.760 93.700 ;
        RECT 141.930 93.520 142.080 93.700 ;
        RECT 6.340 93.220 9.070 93.250 ;
        RECT 6.340 93.050 6.510 93.220 ;
        RECT 6.680 93.050 6.950 93.220 ;
        RECT 7.120 93.050 7.360 93.220 ;
        RECT 7.530 93.050 7.790 93.220 ;
        RECT 7.960 93.050 8.230 93.220 ;
        RECT 8.400 93.050 8.640 93.220 ;
        RECT 8.810 93.050 9.070 93.220 ;
        RECT 6.340 92.250 9.070 93.050 ;
        RECT 9.770 93.210 11.380 93.240 ;
        RECT 13.510 93.210 14.760 93.240 ;
        RECT 15.940 93.220 18.670 93.250 ;
        RECT 9.770 93.040 9.820 93.210 ;
        RECT 9.990 93.040 10.260 93.210 ;
        RECT 10.430 93.040 10.700 93.210 ;
        RECT 10.870 93.040 11.110 93.210 ;
        RECT 11.280 93.040 11.380 93.210 ;
        RECT 9.770 92.760 11.380 93.040 ;
        RECT 10.080 92.360 11.380 92.760 ;
        RECT 6.500 91.580 6.830 92.250 ;
        RECT 7.230 90.930 7.560 91.910 ;
        RECT 7.780 91.580 8.110 92.250 ;
        RECT 8.510 90.930 8.840 91.910 ;
        RECT 10.080 91.580 10.410 92.360 ;
        RECT 6.260 90.050 9.000 90.930 ;
        RECT 10.620 90.920 10.950 91.910 ;
      LAYER li1 ;
        RECT 13.080 91.430 13.330 93.110 ;
      LAYER li1 ;
        RECT 13.680 93.040 13.870 93.210 ;
        RECT 14.040 93.040 14.230 93.210 ;
        RECT 14.400 93.040 14.590 93.210 ;
        RECT 13.510 92.670 14.760 93.040 ;
        RECT 14.940 92.490 15.190 93.110 ;
        RECT 13.640 92.320 15.190 92.490 ;
        RECT 13.640 91.860 13.970 92.320 ;
        RECT 6.260 89.880 6.470 90.050 ;
        RECT 6.640 89.880 6.910 90.050 ;
        RECT 7.080 89.880 7.320 90.050 ;
        RECT 7.490 89.880 7.750 90.050 ;
        RECT 7.920 89.880 8.190 90.050 ;
        RECT 8.360 89.880 8.600 90.050 ;
        RECT 8.770 89.880 9.000 90.050 ;
        RECT 6.260 89.860 9.000 89.880 ;
        RECT 9.850 90.050 11.300 90.920 ;
        RECT 9.850 89.880 10.100 90.050 ;
        RECT 10.270 89.880 10.460 90.050 ;
        RECT 10.630 89.880 10.900 90.050 ;
        RECT 11.070 89.880 11.300 90.050 ;
        RECT 9.850 89.850 11.300 89.880 ;
      LAYER li1 ;
        RECT 13.080 89.850 13.510 91.430 ;
      LAYER li1 ;
        RECT 13.690 90.100 14.250 91.430 ;
      LAYER li1 ;
        RECT 14.430 90.350 14.760 92.140 ;
      LAYER li1 ;
        RECT 14.940 90.600 15.190 92.320 ;
        RECT 15.940 93.050 16.110 93.220 ;
        RECT 16.280 93.050 16.550 93.220 ;
        RECT 16.720 93.050 16.960 93.220 ;
        RECT 17.130 93.050 17.390 93.220 ;
        RECT 17.560 93.050 17.830 93.220 ;
        RECT 18.000 93.050 18.240 93.220 ;
        RECT 18.410 93.050 18.670 93.220 ;
        RECT 15.940 92.250 18.670 93.050 ;
        RECT 19.780 93.220 22.510 93.250 ;
        RECT 19.780 93.050 19.950 93.220 ;
        RECT 20.120 93.050 20.390 93.220 ;
        RECT 20.560 93.050 20.800 93.220 ;
        RECT 20.970 93.050 21.230 93.220 ;
        RECT 21.400 93.050 21.670 93.220 ;
        RECT 21.840 93.050 22.080 93.220 ;
        RECT 22.250 93.050 22.510 93.220 ;
        RECT 19.780 92.250 22.510 93.050 ;
        RECT 24.090 93.210 24.680 93.240 ;
        RECT 24.090 93.040 24.120 93.210 ;
        RECT 24.290 93.040 24.480 93.210 ;
        RECT 24.650 93.040 24.680 93.210 ;
        RECT 25.610 93.210 27.220 93.240 ;
        RECT 24.090 92.280 24.680 93.040 ;
        RECT 16.100 91.580 16.430 92.250 ;
        RECT 16.830 90.930 17.160 91.910 ;
        RECT 17.380 91.580 17.710 92.250 ;
        RECT 18.110 90.930 18.440 91.910 ;
        RECT 19.940 91.580 20.270 92.250 ;
        RECT 20.670 90.930 21.000 91.910 ;
        RECT 21.220 91.580 21.550 92.250 ;
        RECT 21.950 90.930 22.280 91.910 ;
      LAYER li1 ;
        RECT 24.130 91.670 24.840 92.060 ;
        RECT 25.020 91.430 25.350 93.110 ;
      LAYER li1 ;
        RECT 25.610 93.040 25.660 93.210 ;
        RECT 25.830 93.040 26.100 93.210 ;
        RECT 26.270 93.040 26.540 93.210 ;
        RECT 26.710 93.040 26.950 93.210 ;
        RECT 27.120 93.040 27.220 93.210 ;
        RECT 25.610 92.760 27.220 93.040 ;
        RECT 25.920 92.360 27.220 92.760 ;
        RECT 27.520 93.170 29.330 93.340 ;
        RECT 25.920 91.580 26.250 92.360 ;
        RECT 27.520 92.250 27.850 93.170 ;
      LAYER li1 ;
        RECT 28.100 92.770 28.630 92.990 ;
        RECT 28.100 92.600 28.640 92.770 ;
        RECT 28.100 92.250 28.630 92.600 ;
      LAYER li1 ;
        RECT 13.690 89.930 13.700 90.100 ;
        RECT 13.870 89.930 14.060 90.100 ;
        RECT 14.230 89.930 14.250 90.100 ;
        RECT 13.690 89.850 14.250 89.930 ;
        RECT 15.860 90.050 18.600 90.930 ;
        RECT 15.860 89.880 16.070 90.050 ;
        RECT 16.240 89.880 16.510 90.050 ;
        RECT 16.680 89.880 16.920 90.050 ;
        RECT 17.090 89.880 17.350 90.050 ;
        RECT 17.520 89.880 17.790 90.050 ;
        RECT 17.960 89.880 18.200 90.050 ;
        RECT 18.370 89.880 18.600 90.050 ;
        RECT 15.860 89.860 18.600 89.880 ;
        RECT 19.700 90.050 22.440 90.930 ;
        RECT 19.700 89.880 19.910 90.050 ;
        RECT 20.080 89.880 20.350 90.050 ;
        RECT 20.520 89.880 20.760 90.050 ;
        RECT 20.930 89.880 21.190 90.050 ;
        RECT 21.360 89.880 21.630 90.050 ;
        RECT 21.800 89.880 22.040 90.050 ;
        RECT 22.210 89.880 22.440 90.050 ;
        RECT 19.700 89.860 22.440 89.880 ;
        RECT 24.090 90.100 24.680 91.430 ;
        RECT 24.090 89.930 24.120 90.100 ;
        RECT 24.290 89.930 24.480 90.100 ;
        RECT 24.650 89.930 24.680 90.100 ;
        RECT 24.090 89.850 24.680 89.930 ;
      LAYER li1 ;
        RECT 24.960 89.850 25.350 91.430 ;
      LAYER li1 ;
        RECT 26.460 90.920 26.790 91.910 ;
      LAYER li1 ;
        RECT 27.490 91.740 27.910 92.070 ;
        RECT 28.100 91.680 28.270 92.250 ;
      LAYER li1 ;
        RECT 29.160 92.150 29.330 93.170 ;
        RECT 29.510 93.210 30.610 93.240 ;
        RECT 29.510 93.040 29.560 93.210 ;
        RECT 29.730 93.040 29.920 93.210 ;
        RECT 30.090 93.040 30.280 93.210 ;
        RECT 30.450 93.040 30.610 93.210 ;
        RECT 31.370 93.210 32.980 93.240 ;
        RECT 33.670 93.210 34.920 93.240 ;
        RECT 35.690 93.210 37.300 93.240 ;
        RECT 29.510 92.330 30.610 93.040 ;
        RECT 30.780 92.150 31.030 93.080 ;
        RECT 31.370 93.040 31.420 93.210 ;
        RECT 31.590 93.040 31.860 93.210 ;
        RECT 32.030 93.040 32.300 93.210 ;
        RECT 32.470 93.040 32.710 93.210 ;
        RECT 32.880 93.040 32.980 93.210 ;
        RECT 31.370 92.760 32.980 93.040 ;
      LAYER li1 ;
        RECT 28.450 91.860 28.960 92.070 ;
      LAYER li1 ;
        RECT 29.160 91.980 31.030 92.150 ;
        RECT 31.680 92.360 32.980 92.760 ;
      LAYER li1 ;
        RECT 28.100 91.510 29.160 91.680 ;
        RECT 28.890 91.430 29.160 91.510 ;
        RECT 29.610 91.490 30.120 91.800 ;
        RECT 30.370 91.490 31.080 91.800 ;
      LAYER li1 ;
        RECT 31.680 91.580 32.010 92.360 ;
        RECT 25.690 90.050 27.140 90.920 ;
        RECT 25.690 89.880 25.940 90.050 ;
        RECT 26.110 89.880 26.300 90.050 ;
        RECT 26.470 89.880 26.740 90.050 ;
        RECT 26.910 89.880 27.140 90.050 ;
        RECT 25.690 89.850 27.140 89.880 ;
        RECT 27.450 90.100 28.710 91.330 ;
      LAYER li1 ;
        RECT 28.890 90.350 29.410 91.430 ;
      LAYER li1 ;
        RECT 27.450 89.930 27.460 90.100 ;
        RECT 27.630 89.930 27.820 90.100 ;
        RECT 27.990 89.930 28.180 90.100 ;
        RECT 28.350 89.930 28.540 90.100 ;
        RECT 27.450 89.850 28.710 89.930 ;
      LAYER li1 ;
        RECT 29.240 89.850 29.410 90.350 ;
      LAYER li1 ;
        RECT 29.670 90.100 30.980 91.310 ;
        RECT 32.220 90.920 32.550 91.910 ;
      LAYER li1 ;
        RECT 33.240 91.430 33.490 93.110 ;
      LAYER li1 ;
        RECT 33.840 93.040 34.030 93.210 ;
        RECT 34.200 93.040 34.390 93.210 ;
        RECT 34.560 93.040 34.750 93.210 ;
        RECT 33.670 92.670 34.920 93.040 ;
        RECT 35.100 92.490 35.350 93.110 ;
        RECT 35.690 93.040 35.740 93.210 ;
        RECT 35.910 93.040 36.180 93.210 ;
        RECT 36.350 93.040 36.620 93.210 ;
        RECT 36.790 93.040 37.030 93.210 ;
        RECT 37.200 93.040 37.300 93.210 ;
        RECT 35.690 92.760 37.300 93.040 ;
        RECT 38.010 93.210 38.600 93.240 ;
        RECT 38.010 93.040 38.040 93.210 ;
        RECT 38.210 93.040 38.400 93.210 ;
        RECT 38.570 93.040 38.600 93.210 ;
        RECT 33.800 92.320 35.350 92.490 ;
        RECT 33.800 91.860 34.130 92.320 ;
        RECT 29.670 89.930 29.700 90.100 ;
        RECT 29.870 89.930 30.060 90.100 ;
        RECT 30.230 89.930 30.420 90.100 ;
        RECT 30.590 89.930 30.780 90.100 ;
        RECT 30.950 89.930 30.980 90.100 ;
        RECT 29.670 89.850 30.980 89.930 ;
        RECT 31.450 90.050 32.900 90.920 ;
        RECT 31.450 89.880 31.700 90.050 ;
        RECT 31.870 89.880 32.060 90.050 ;
        RECT 32.230 89.880 32.500 90.050 ;
        RECT 32.670 89.880 32.900 90.050 ;
        RECT 31.450 89.850 32.900 89.880 ;
      LAYER li1 ;
        RECT 33.240 89.850 33.670 91.430 ;
      LAYER li1 ;
        RECT 33.850 90.100 34.410 91.430 ;
      LAYER li1 ;
        RECT 34.590 90.350 34.920 92.140 ;
      LAYER li1 ;
        RECT 35.100 90.600 35.350 92.320 ;
        RECT 36.000 92.360 37.300 92.760 ;
        RECT 36.000 91.580 36.330 92.360 ;
        RECT 37.560 92.310 37.820 92.990 ;
        RECT 38.010 92.490 38.600 93.040 ;
        RECT 38.780 93.170 39.730 93.340 ;
        RECT 39.910 93.210 40.450 93.240 ;
        RECT 38.780 92.310 38.950 93.170 ;
        RECT 37.560 92.140 38.950 92.310 ;
        RECT 36.540 90.920 36.870 91.910 ;
        RECT 33.850 89.930 33.860 90.100 ;
        RECT 34.030 89.930 34.220 90.100 ;
        RECT 34.390 89.930 34.410 90.100 ;
        RECT 33.850 89.850 34.410 89.930 ;
        RECT 35.770 90.050 37.220 90.920 ;
        RECT 35.770 89.880 36.020 90.050 ;
        RECT 36.190 89.880 36.380 90.050 ;
        RECT 36.550 89.880 36.820 90.050 ;
        RECT 36.990 89.880 37.220 90.050 ;
        RECT 35.770 89.850 37.220 89.880 ;
        RECT 37.560 89.870 37.810 92.140 ;
        RECT 38.620 91.710 38.950 92.140 ;
        RECT 39.130 91.330 39.380 92.990 ;
        RECT 39.560 92.430 39.730 93.170 ;
        RECT 40.080 93.040 40.270 93.210 ;
        RECT 40.440 93.040 40.450 93.210 ;
        RECT 42.300 93.210 43.250 93.240 ;
        RECT 39.910 92.610 40.450 93.040 ;
        RECT 40.630 92.610 40.980 93.110 ;
        RECT 39.560 92.260 40.630 92.430 ;
      LAYER li1 ;
        RECT 39.950 91.510 40.280 92.080 ;
      LAYER li1 ;
        RECT 39.130 91.160 40.280 91.330 ;
        RECT 37.990 90.100 38.940 90.680 ;
        RECT 39.130 90.660 39.450 91.160 ;
        RECT 37.990 89.930 38.020 90.100 ;
        RECT 38.190 89.930 38.380 90.100 ;
        RECT 38.550 89.930 38.740 90.100 ;
        RECT 38.910 89.930 38.940 90.100 ;
        RECT 37.990 89.850 38.940 89.930 ;
        RECT 39.120 89.870 39.450 90.660 ;
        RECT 39.680 90.100 39.930 90.980 ;
        RECT 39.680 89.930 39.710 90.100 ;
        RECT 39.880 89.930 39.930 90.100 ;
        RECT 39.680 89.900 39.930 89.930 ;
        RECT 40.110 89.850 40.280 91.160 ;
        RECT 40.460 90.320 40.630 92.260 ;
        RECT 40.810 90.500 40.980 92.610 ;
        RECT 41.510 92.640 41.760 93.110 ;
        RECT 42.300 93.040 42.330 93.210 ;
        RECT 42.500 93.040 42.690 93.210 ;
        RECT 42.860 93.040 43.050 93.210 ;
        RECT 43.220 93.040 43.250 93.210 ;
        RECT 42.300 92.820 43.250 93.040 ;
        RECT 43.430 92.640 43.760 93.340 ;
        RECT 41.160 90.320 41.330 92.520 ;
        RECT 41.510 92.470 43.760 92.640 ;
        RECT 44.240 93.210 45.190 93.240 ;
        RECT 44.240 93.040 44.270 93.210 ;
        RECT 44.440 93.040 44.630 93.210 ;
        RECT 44.800 93.040 44.990 93.210 ;
        RECT 45.160 93.040 45.190 93.210 ;
        RECT 48.780 93.210 49.370 93.240 ;
        RECT 41.510 91.000 41.680 92.470 ;
        RECT 41.860 91.800 42.100 92.110 ;
        RECT 42.580 91.980 43.310 92.290 ;
        RECT 44.240 92.230 45.190 93.040 ;
      LAYER li1 ;
        RECT 45.730 92.770 48.600 93.050 ;
        RECT 45.370 92.600 48.600 92.770 ;
        RECT 45.370 92.050 45.540 92.600 ;
        RECT 48.330 92.570 48.600 92.600 ;
      LAYER li1 ;
        RECT 48.780 93.040 48.810 93.210 ;
        RECT 48.980 93.040 49.170 93.210 ;
        RECT 49.340 93.040 49.370 93.210 ;
        RECT 46.470 92.130 47.100 92.420 ;
        RECT 48.780 92.130 49.370 93.040 ;
        RECT 50.700 93.210 51.650 93.240 ;
        RECT 50.700 93.040 50.730 93.210 ;
        RECT 50.900 93.040 51.090 93.210 ;
        RECT 51.260 93.040 51.450 93.210 ;
        RECT 51.620 93.040 51.650 93.210 ;
      LAYER li1 ;
        RECT 44.610 91.810 45.540 92.050 ;
      LAYER li1 ;
        RECT 45.720 91.900 46.230 92.060 ;
        RECT 41.860 91.630 44.430 91.800 ;
        RECT 45.720 91.730 46.750 91.900 ;
        RECT 45.720 91.630 45.890 91.730 ;
        RECT 41.860 91.440 42.100 91.630 ;
        RECT 44.260 91.460 45.890 91.630 ;
        RECT 42.280 91.280 44.080 91.450 ;
        RECT 46.070 91.280 46.400 91.520 ;
        RECT 41.510 90.500 41.840 91.000 ;
        RECT 42.280 90.320 42.450 91.280 ;
        RECT 43.910 91.110 46.400 91.280 ;
        RECT 40.460 89.990 42.450 90.320 ;
        RECT 42.630 90.930 43.730 91.100 ;
        RECT 46.580 90.930 46.750 91.730 ;
        RECT 42.630 90.050 42.870 90.930 ;
        RECT 43.560 90.760 44.340 90.930 ;
        RECT 43.050 90.100 43.380 90.750 ;
        RECT 44.010 90.500 44.340 90.760 ;
        RECT 43.050 89.930 43.080 90.100 ;
        RECT 43.250 89.930 43.380 90.100 ;
        RECT 43.050 89.900 43.380 89.930 ;
        RECT 44.520 90.100 45.470 90.930 ;
        RECT 44.520 89.930 44.550 90.100 ;
        RECT 44.720 89.930 44.910 90.100 ;
        RECT 45.080 89.930 45.270 90.100 ;
        RECT 45.440 89.930 45.470 90.100 ;
        RECT 44.520 89.900 45.470 89.930 ;
        RECT 46.140 90.760 46.750 90.930 ;
        RECT 46.930 91.290 47.100 92.130 ;
        RECT 47.750 91.950 48.080 92.060 ;
        RECT 49.560 91.950 49.890 92.630 ;
        RECT 50.190 92.130 50.520 92.630 ;
        RECT 50.700 92.130 51.650 93.040 ;
        RECT 52.900 93.220 55.630 93.250 ;
        RECT 52.900 93.050 53.070 93.220 ;
        RECT 53.240 93.050 53.510 93.220 ;
        RECT 53.680 93.050 53.920 93.220 ;
        RECT 54.090 93.050 54.350 93.220 ;
        RECT 54.520 93.050 54.790 93.220 ;
        RECT 54.960 93.050 55.200 93.220 ;
        RECT 55.370 93.050 55.630 93.220 ;
        RECT 57.200 93.210 58.150 93.240 ;
        RECT 52.900 92.250 55.630 93.050 ;
        RECT 47.750 91.780 50.000 91.950 ;
        RECT 47.750 91.470 48.080 91.780 ;
        RECT 49.320 91.290 49.650 91.600 ;
        RECT 46.930 91.120 49.650 91.290 ;
        RECT 46.140 90.010 46.310 90.760 ;
        RECT 46.930 90.580 47.100 91.120 ;
        RECT 46.490 90.190 47.100 90.580 ;
        RECT 47.450 90.100 48.400 90.940 ;
        RECT 48.850 90.930 49.650 91.120 ;
        RECT 48.850 90.780 49.180 90.930 ;
        RECT 49.830 90.600 50.000 91.780 ;
        RECT 48.820 90.430 50.000 90.600 ;
        RECT 50.310 91.380 50.520 92.130 ;
        RECT 51.350 91.380 51.680 91.880 ;
        RECT 53.060 91.580 53.390 92.250 ;
        RECT 50.310 91.210 51.680 91.380 ;
        RECT 48.820 90.350 48.990 90.430 ;
        RECT 46.140 89.800 47.270 90.010 ;
        RECT 47.450 89.930 47.480 90.100 ;
        RECT 47.650 89.930 47.840 90.100 ;
        RECT 48.010 89.930 48.200 90.100 ;
        RECT 48.370 89.930 48.400 90.100 ;
        RECT 47.450 89.900 48.400 89.930 ;
        RECT 48.740 89.850 48.990 90.350 ;
        RECT 49.170 90.100 50.120 90.250 ;
        RECT 50.310 90.240 50.560 91.210 ;
        RECT 49.170 89.930 49.200 90.100 ;
        RECT 49.370 89.930 49.560 90.100 ;
        RECT 49.730 89.930 49.920 90.100 ;
        RECT 50.090 89.930 50.120 90.100 ;
        RECT 49.170 89.870 50.120 89.930 ;
        RECT 50.740 90.100 51.680 91.030 ;
        RECT 53.790 90.930 54.120 91.910 ;
        RECT 54.340 91.580 54.670 92.250 ;
        RECT 55.070 90.930 55.400 91.910 ;
        RECT 56.750 91.250 57.020 93.110 ;
        RECT 57.200 93.040 57.230 93.210 ;
        RECT 57.400 93.040 57.590 93.210 ;
        RECT 57.760 93.040 57.950 93.210 ;
        RECT 58.120 93.040 58.150 93.210 ;
        RECT 58.840 93.210 59.430 93.240 ;
        RECT 57.200 92.610 58.150 93.040 ;
        RECT 58.330 92.610 58.660 93.110 ;
      LAYER li1 ;
        RECT 57.200 91.460 57.530 92.430 ;
      LAYER li1 ;
        RECT 57.880 91.250 58.210 91.750 ;
        RECT 56.750 91.080 58.210 91.250 ;
        RECT 50.740 89.930 50.760 90.100 ;
        RECT 50.930 89.930 51.120 90.100 ;
        RECT 51.290 89.930 51.480 90.100 ;
        RECT 51.650 89.930 51.680 90.100 ;
        RECT 50.740 89.900 51.680 89.930 ;
        RECT 52.820 90.050 55.560 90.930 ;
        RECT 56.750 90.150 57.080 91.080 ;
        RECT 52.820 89.880 53.030 90.050 ;
        RECT 53.200 89.880 53.470 90.050 ;
        RECT 53.640 89.880 53.880 90.050 ;
        RECT 54.050 89.880 54.310 90.050 ;
        RECT 54.480 89.880 54.750 90.050 ;
        RECT 54.920 89.880 55.160 90.050 ;
        RECT 55.330 89.880 55.560 90.050 ;
        RECT 57.270 90.100 57.860 90.880 ;
        RECT 57.270 89.930 57.300 90.100 ;
        RECT 57.470 89.930 57.660 90.100 ;
        RECT 57.830 89.930 57.860 90.100 ;
        RECT 57.270 89.900 57.860 89.930 ;
        RECT 58.040 89.970 58.210 91.080 ;
        RECT 58.390 91.690 58.660 92.610 ;
        RECT 58.840 93.040 58.870 93.210 ;
        RECT 59.040 93.040 59.230 93.210 ;
        RECT 59.400 93.040 59.430 93.210 ;
        RECT 63.800 93.210 64.750 93.240 ;
        RECT 58.840 92.360 59.430 93.040 ;
      LAYER li1 ;
        RECT 59.710 92.980 62.650 93.150 ;
        RECT 59.710 91.990 59.880 92.980 ;
      LAYER li1 ;
        RECT 58.390 91.460 58.920 91.690 ;
        RECT 58.390 90.150 58.640 91.460 ;
      LAYER li1 ;
        RECT 59.340 91.120 59.880 91.990 ;
        RECT 60.060 91.500 60.390 92.800 ;
      LAYER li1 ;
        RECT 60.570 92.280 60.840 92.780 ;
        RECT 61.290 92.530 61.620 92.780 ;
        RECT 61.290 92.360 62.300 92.530 ;
        RECT 60.570 91.290 60.740 92.280 ;
        RECT 61.620 91.690 61.950 92.180 ;
        RECT 60.520 91.120 60.740 91.290 ;
        RECT 60.920 91.460 61.950 91.690 ;
        RECT 62.130 92.130 62.300 92.360 ;
      LAYER li1 ;
        RECT 62.480 92.480 62.650 92.980 ;
      LAYER li1 ;
        RECT 63.800 93.040 63.830 93.210 ;
        RECT 64.000 93.040 64.190 93.210 ;
        RECT 64.360 93.040 64.550 93.210 ;
        RECT 64.720 93.040 64.750 93.210 ;
        RECT 63.800 92.660 64.750 93.040 ;
      LAYER li1 ;
        RECT 64.930 93.170 67.590 93.340 ;
        RECT 64.930 92.480 65.100 93.170 ;
        RECT 62.480 92.310 65.100 92.480 ;
      LAYER li1 ;
        RECT 62.130 91.960 64.750 92.130 ;
        RECT 60.520 90.940 60.690 91.120 ;
        RECT 60.920 90.940 61.090 91.460 ;
        RECT 62.130 91.280 62.300 91.960 ;
      LAYER li1 ;
        RECT 64.930 91.780 65.100 92.310 ;
      LAYER li1 ;
        RECT 58.880 90.770 60.690 90.940 ;
        RECT 58.880 90.150 59.130 90.770 ;
        RECT 59.310 90.420 60.340 90.590 ;
        RECT 59.310 89.970 59.480 90.420 ;
        RECT 52.820 89.860 55.560 89.880 ;
        RECT 58.040 89.800 59.480 89.970 ;
        RECT 59.660 90.100 59.990 90.240 ;
        RECT 59.660 89.930 59.690 90.100 ;
        RECT 59.860 89.930 59.990 90.100 ;
        RECT 59.660 89.900 59.990 89.930 ;
        RECT 60.170 89.970 60.340 90.420 ;
        RECT 60.520 90.150 60.690 90.770 ;
        RECT 60.870 90.610 61.090 90.940 ;
        RECT 61.270 91.110 62.300 91.280 ;
        RECT 62.480 91.430 62.810 91.780 ;
      LAYER li1 ;
        RECT 63.250 91.610 65.100 91.780 ;
      LAYER li1 ;
        RECT 65.280 92.280 65.610 92.990 ;
        RECT 66.070 92.820 67.240 92.990 ;
        RECT 66.070 92.280 66.400 92.820 ;
        RECT 65.280 91.430 65.540 92.280 ;
        RECT 66.610 92.020 66.890 92.520 ;
        RECT 62.480 91.260 65.540 91.430 ;
        RECT 61.270 90.410 61.440 91.110 ;
        RECT 62.130 91.080 62.300 91.110 ;
        RECT 61.620 90.730 61.950 90.930 ;
        RECT 62.130 90.910 63.900 91.080 ;
        RECT 61.620 90.610 63.390 90.730 ;
        RECT 61.740 90.560 63.390 90.610 ;
        RECT 61.220 90.150 61.550 90.410 ;
        RECT 61.740 89.970 61.910 90.560 ;
        RECT 60.170 89.800 61.910 89.970 ;
        RECT 62.090 90.100 63.040 90.380 ;
        RECT 62.090 89.930 62.120 90.100 ;
        RECT 62.290 89.930 62.480 90.100 ;
        RECT 62.650 89.930 62.840 90.100 ;
        RECT 63.010 89.930 63.040 90.100 ;
        RECT 62.090 89.900 63.040 89.930 ;
        RECT 63.220 89.970 63.390 90.560 ;
        RECT 63.570 90.150 63.900 90.910 ;
        RECT 65.210 90.680 65.540 91.260 ;
        RECT 65.720 91.850 66.890 92.020 ;
        RECT 65.720 90.500 65.890 91.850 ;
        RECT 66.270 91.170 66.600 91.670 ;
        RECT 67.070 91.420 67.240 92.820 ;
      LAYER li1 ;
        RECT 67.420 92.510 67.590 93.170 ;
      LAYER li1 ;
        RECT 67.770 93.210 68.720 93.240 ;
        RECT 67.770 93.040 67.800 93.210 ;
        RECT 67.970 93.040 68.160 93.210 ;
        RECT 68.330 93.040 68.520 93.210 ;
        RECT 68.690 93.040 68.720 93.210 ;
        RECT 70.380 93.210 71.330 93.240 ;
        RECT 67.770 92.690 68.720 93.040 ;
        RECT 69.260 92.610 69.590 93.110 ;
        RECT 70.380 93.040 70.410 93.210 ;
        RECT 70.580 93.040 70.770 93.210 ;
        RECT 70.940 93.040 71.130 93.210 ;
        RECT 71.300 93.040 71.330 93.210 ;
      LAYER li1 ;
        RECT 67.420 92.340 68.430 92.510 ;
      LAYER li1 ;
        RECT 67.450 91.770 67.780 92.160 ;
      LAYER li1 ;
        RECT 68.100 91.950 68.430 92.340 ;
      LAYER li1 ;
        RECT 69.260 91.770 69.490 92.610 ;
        RECT 69.870 92.110 70.200 92.610 ;
        RECT 70.380 92.110 71.330 93.040 ;
        RECT 72.170 93.210 73.780 93.240 ;
        RECT 72.170 93.040 72.220 93.210 ;
        RECT 72.390 93.040 72.660 93.210 ;
        RECT 72.830 93.040 73.100 93.210 ;
        RECT 73.270 93.040 73.510 93.210 ;
        RECT 73.680 93.040 73.780 93.210 ;
        RECT 67.450 91.600 69.490 91.770 ;
        RECT 66.780 91.250 69.140 91.420 ;
        RECT 66.780 90.930 66.950 91.250 ;
        RECT 69.320 91.070 69.490 91.600 ;
        RECT 64.080 90.330 65.890 90.500 ;
        RECT 66.070 90.760 66.950 90.930 ;
        RECT 64.080 89.970 64.250 90.330 ;
        RECT 63.220 89.800 64.250 89.970 ;
        RECT 64.430 90.100 65.380 90.150 ;
        RECT 64.430 89.930 64.460 90.100 ;
        RECT 64.630 89.930 64.820 90.100 ;
        RECT 64.990 89.930 65.180 90.100 ;
        RECT 65.350 89.930 65.380 90.100 ;
        RECT 64.430 89.850 65.380 89.930 ;
        RECT 66.070 89.850 66.320 90.760 ;
        RECT 67.130 90.100 68.080 90.930 ;
        RECT 68.480 90.900 69.490 91.070 ;
        RECT 69.990 91.930 70.200 92.110 ;
        RECT 69.990 91.600 71.360 91.930 ;
        RECT 68.480 90.430 68.730 90.900 ;
        RECT 68.910 90.100 69.810 90.720 ;
        RECT 69.990 90.600 70.240 91.600 ;
        RECT 67.130 89.930 67.160 90.100 ;
        RECT 67.330 89.930 67.520 90.100 ;
        RECT 67.690 89.930 67.880 90.100 ;
        RECT 68.050 89.930 68.080 90.100 ;
        RECT 69.080 89.930 69.270 90.100 ;
        RECT 69.440 89.930 69.630 90.100 ;
        RECT 69.800 89.930 69.810 90.100 ;
        RECT 67.130 89.900 68.080 89.930 ;
        RECT 68.910 89.900 69.810 89.930 ;
        RECT 70.420 90.100 71.360 91.410 ;
        RECT 70.420 89.930 70.440 90.100 ;
        RECT 70.610 89.930 70.800 90.100 ;
        RECT 70.970 89.930 71.160 90.100 ;
        RECT 71.330 89.930 71.360 90.100 ;
        RECT 70.420 89.870 71.360 89.930 ;
      LAYER li1 ;
        RECT 71.540 89.870 71.880 92.940 ;
      LAYER li1 ;
        RECT 72.170 92.760 73.780 93.040 ;
        RECT 72.480 92.360 73.780 92.760 ;
        RECT 74.970 93.210 75.920 93.240 ;
        RECT 74.970 93.040 75.000 93.210 ;
        RECT 75.170 93.040 75.360 93.210 ;
        RECT 75.530 93.040 75.720 93.210 ;
        RECT 75.890 93.040 75.920 93.210 ;
        RECT 76.530 93.210 77.480 93.240 ;
        RECT 72.480 91.580 72.810 92.360 ;
        RECT 74.970 92.280 75.920 93.040 ;
      LAYER li1 ;
        RECT 76.100 92.400 76.350 93.110 ;
      LAYER li1 ;
        RECT 76.530 93.040 76.560 93.210 ;
        RECT 76.730 93.040 76.920 93.210 ;
        RECT 77.090 93.040 77.280 93.210 ;
        RECT 77.450 93.040 77.480 93.210 ;
        RECT 78.090 93.210 79.040 93.240 ;
        RECT 76.530 92.580 77.480 93.040 ;
      LAYER li1 ;
        RECT 77.660 92.400 77.910 93.110 ;
        RECT 76.100 92.230 77.910 92.400 ;
      LAYER li1 ;
        RECT 78.090 93.040 78.120 93.210 ;
        RECT 78.290 93.040 78.480 93.210 ;
        RECT 78.650 93.040 78.840 93.210 ;
        RECT 79.010 93.040 79.040 93.210 ;
        RECT 79.850 93.210 81.460 93.240 ;
        RECT 78.090 92.360 79.040 93.040 ;
      LAYER li1 ;
        RECT 76.100 92.060 76.270 92.230 ;
      LAYER li1 ;
        RECT 79.220 92.180 79.550 93.110 ;
        RECT 79.850 93.040 79.900 93.210 ;
        RECT 80.070 93.040 80.340 93.210 ;
        RECT 80.510 93.040 80.780 93.210 ;
        RECT 80.950 93.040 81.190 93.210 ;
        RECT 81.360 93.040 81.460 93.210 ;
        RECT 79.850 92.760 81.460 93.040 ;
        RECT 73.020 90.920 73.350 91.910 ;
      LAYER li1 ;
        RECT 75.010 91.830 76.270 92.060 ;
      LAYER li1 ;
        RECT 78.310 92.050 79.550 92.180 ;
        RECT 76.450 92.010 79.550 92.050 ;
        RECT 76.450 91.880 78.480 92.010 ;
      LAYER li1 ;
        RECT 76.100 91.700 76.270 91.830 ;
        RECT 76.100 91.530 77.990 91.700 ;
      LAYER li1 ;
        RECT 72.250 90.050 73.700 90.920 ;
        RECT 72.250 89.880 72.500 90.050 ;
        RECT 72.670 89.880 72.860 90.050 ;
        RECT 73.030 89.880 73.300 90.050 ;
        RECT 73.470 89.880 73.700 90.050 ;
        RECT 72.250 89.850 73.700 89.880 ;
        RECT 74.970 90.100 75.920 91.430 ;
        RECT 74.970 89.930 75.000 90.100 ;
        RECT 75.170 89.930 75.360 90.100 ;
        RECT 75.530 89.930 75.720 90.100 ;
        RECT 75.890 89.930 75.920 90.100 ;
        RECT 74.970 89.850 75.920 89.930 ;
      LAYER li1 ;
        RECT 76.100 89.850 76.350 91.530 ;
      LAYER li1 ;
        RECT 76.530 90.100 77.480 91.350 ;
        RECT 76.530 89.930 76.560 90.100 ;
        RECT 76.730 89.930 76.920 90.100 ;
        RECT 77.090 89.930 77.280 90.100 ;
        RECT 77.450 89.930 77.480 90.100 ;
        RECT 76.530 89.850 77.480 89.930 ;
      LAYER li1 ;
        RECT 77.660 89.850 77.990 91.530 ;
        RECT 78.770 91.490 79.100 91.830 ;
      LAYER li1 ;
        RECT 78.170 90.100 79.120 91.310 ;
        RECT 78.170 89.930 78.200 90.100 ;
        RECT 78.370 89.930 78.560 90.100 ;
        RECT 78.730 89.930 78.920 90.100 ;
        RECT 79.090 89.930 79.120 90.100 ;
        RECT 78.170 89.850 79.120 89.930 ;
        RECT 79.300 89.850 79.550 92.010 ;
        RECT 80.160 92.360 81.460 92.760 ;
        RECT 81.690 93.210 82.640 93.240 ;
        RECT 81.690 93.040 81.720 93.210 ;
        RECT 81.890 93.040 82.080 93.210 ;
        RECT 82.250 93.040 82.440 93.210 ;
        RECT 82.610 93.040 82.640 93.210 ;
        RECT 83.250 93.210 84.200 93.240 ;
        RECT 80.160 91.580 80.490 92.360 ;
        RECT 81.690 92.280 82.640 93.040 ;
      LAYER li1 ;
        RECT 82.820 92.400 83.070 93.110 ;
      LAYER li1 ;
        RECT 83.250 93.040 83.280 93.210 ;
        RECT 83.450 93.040 83.640 93.210 ;
        RECT 83.810 93.040 84.000 93.210 ;
        RECT 84.170 93.040 84.200 93.210 ;
        RECT 84.810 93.210 85.760 93.240 ;
        RECT 83.250 92.580 84.200 93.040 ;
      LAYER li1 ;
        RECT 84.380 92.400 84.630 93.110 ;
        RECT 82.820 92.230 84.630 92.400 ;
      LAYER li1 ;
        RECT 84.810 93.040 84.840 93.210 ;
        RECT 85.010 93.040 85.200 93.210 ;
        RECT 85.370 93.040 85.560 93.210 ;
        RECT 85.730 93.040 85.760 93.210 ;
        RECT 86.570 93.210 88.180 93.240 ;
        RECT 84.810 92.360 85.760 93.040 ;
      LAYER li1 ;
        RECT 82.820 92.060 82.990 92.230 ;
      LAYER li1 ;
        RECT 85.940 92.180 86.270 93.110 ;
        RECT 86.570 93.040 86.620 93.210 ;
        RECT 86.790 93.040 87.060 93.210 ;
        RECT 87.230 93.040 87.500 93.210 ;
        RECT 87.670 93.040 87.910 93.210 ;
        RECT 88.080 93.040 88.180 93.210 ;
        RECT 86.570 92.760 88.180 93.040 ;
        RECT 80.700 90.920 81.030 91.910 ;
      LAYER li1 ;
        RECT 81.730 91.830 82.990 92.060 ;
      LAYER li1 ;
        RECT 85.030 92.050 86.270 92.180 ;
        RECT 83.170 92.010 86.270 92.050 ;
        RECT 83.170 91.880 85.200 92.010 ;
      LAYER li1 ;
        RECT 82.820 91.700 82.990 91.830 ;
        RECT 82.820 91.530 84.710 91.700 ;
      LAYER li1 ;
        RECT 79.930 90.050 81.380 90.920 ;
        RECT 79.930 89.880 80.180 90.050 ;
        RECT 80.350 89.880 80.540 90.050 ;
        RECT 80.710 89.880 80.980 90.050 ;
        RECT 81.150 89.880 81.380 90.050 ;
        RECT 79.930 89.850 81.380 89.880 ;
        RECT 81.690 90.100 82.640 91.430 ;
        RECT 81.690 89.930 81.720 90.100 ;
        RECT 81.890 89.930 82.080 90.100 ;
        RECT 82.250 89.930 82.440 90.100 ;
        RECT 82.610 89.930 82.640 90.100 ;
        RECT 81.690 89.850 82.640 89.930 ;
      LAYER li1 ;
        RECT 82.820 89.850 83.070 91.530 ;
      LAYER li1 ;
        RECT 83.250 90.100 84.200 91.350 ;
        RECT 83.250 89.930 83.280 90.100 ;
        RECT 83.450 89.930 83.640 90.100 ;
        RECT 83.810 89.930 84.000 90.100 ;
        RECT 84.170 89.930 84.200 90.100 ;
        RECT 83.250 89.850 84.200 89.930 ;
      LAYER li1 ;
        RECT 84.380 89.850 84.710 91.530 ;
        RECT 85.490 91.490 85.820 91.830 ;
      LAYER li1 ;
        RECT 84.890 90.100 85.840 91.310 ;
        RECT 84.890 89.930 84.920 90.100 ;
        RECT 85.090 89.930 85.280 90.100 ;
        RECT 85.450 89.930 85.640 90.100 ;
        RECT 85.810 89.930 85.840 90.100 ;
        RECT 84.890 89.850 85.840 89.930 ;
        RECT 86.020 89.850 86.270 92.010 ;
        RECT 86.880 92.360 88.180 92.760 ;
        RECT 88.410 93.210 89.360 93.240 ;
        RECT 88.410 93.040 88.440 93.210 ;
        RECT 88.610 93.040 88.800 93.210 ;
        RECT 88.970 93.040 89.160 93.210 ;
        RECT 89.330 93.040 89.360 93.210 ;
        RECT 89.970 93.210 90.920 93.240 ;
        RECT 86.880 91.580 87.210 92.360 ;
        RECT 88.410 92.280 89.360 93.040 ;
      LAYER li1 ;
        RECT 89.540 92.400 89.790 93.110 ;
      LAYER li1 ;
        RECT 89.970 93.040 90.000 93.210 ;
        RECT 90.170 93.040 90.360 93.210 ;
        RECT 90.530 93.040 90.720 93.210 ;
        RECT 90.890 93.040 90.920 93.210 ;
        RECT 91.530 93.210 92.480 93.240 ;
        RECT 89.970 92.580 90.920 93.040 ;
      LAYER li1 ;
        RECT 91.100 92.400 91.350 93.110 ;
        RECT 89.540 92.230 91.350 92.400 ;
      LAYER li1 ;
        RECT 91.530 93.040 91.560 93.210 ;
        RECT 91.730 93.040 91.920 93.210 ;
        RECT 92.090 93.040 92.280 93.210 ;
        RECT 92.450 93.040 92.480 93.210 ;
        RECT 93.290 93.210 94.900 93.240 ;
        RECT 91.530 92.360 92.480 93.040 ;
      LAYER li1 ;
        RECT 89.540 92.060 89.710 92.230 ;
      LAYER li1 ;
        RECT 92.660 92.180 92.990 93.110 ;
        RECT 93.290 93.040 93.340 93.210 ;
        RECT 93.510 93.040 93.780 93.210 ;
        RECT 93.950 93.040 94.220 93.210 ;
        RECT 94.390 93.040 94.630 93.210 ;
        RECT 94.800 93.040 94.900 93.210 ;
        RECT 93.290 92.760 94.900 93.040 ;
        RECT 87.420 90.920 87.750 91.910 ;
      LAYER li1 ;
        RECT 88.450 91.830 89.710 92.060 ;
      LAYER li1 ;
        RECT 91.750 92.050 92.990 92.180 ;
        RECT 89.890 92.010 92.990 92.050 ;
        RECT 89.890 91.880 91.920 92.010 ;
      LAYER li1 ;
        RECT 89.540 91.700 89.710 91.830 ;
        RECT 89.540 91.530 91.430 91.700 ;
      LAYER li1 ;
        RECT 86.650 90.050 88.100 90.920 ;
        RECT 86.650 89.880 86.900 90.050 ;
        RECT 87.070 89.880 87.260 90.050 ;
        RECT 87.430 89.880 87.700 90.050 ;
        RECT 87.870 89.880 88.100 90.050 ;
        RECT 86.650 89.850 88.100 89.880 ;
        RECT 88.410 90.100 89.360 91.430 ;
        RECT 88.410 89.930 88.440 90.100 ;
        RECT 88.610 89.930 88.800 90.100 ;
        RECT 88.970 89.930 89.160 90.100 ;
        RECT 89.330 89.930 89.360 90.100 ;
        RECT 88.410 89.850 89.360 89.930 ;
      LAYER li1 ;
        RECT 89.540 89.850 89.790 91.530 ;
      LAYER li1 ;
        RECT 89.970 90.100 90.920 91.350 ;
        RECT 89.970 89.930 90.000 90.100 ;
        RECT 90.170 89.930 90.360 90.100 ;
        RECT 90.530 89.930 90.720 90.100 ;
        RECT 90.890 89.930 90.920 90.100 ;
        RECT 89.970 89.850 90.920 89.930 ;
      LAYER li1 ;
        RECT 91.100 89.850 91.430 91.530 ;
        RECT 92.210 91.490 92.540 91.830 ;
      LAYER li1 ;
        RECT 91.610 90.100 92.560 91.310 ;
        RECT 91.610 89.930 91.640 90.100 ;
        RECT 91.810 89.930 92.000 90.100 ;
        RECT 92.170 89.930 92.360 90.100 ;
        RECT 92.530 89.930 92.560 90.100 ;
        RECT 91.610 89.850 92.560 89.930 ;
        RECT 92.740 89.850 92.990 92.010 ;
        RECT 93.600 92.360 94.900 92.760 ;
        RECT 95.130 93.210 96.080 93.240 ;
        RECT 95.130 93.040 95.160 93.210 ;
        RECT 95.330 93.040 95.520 93.210 ;
        RECT 95.690 93.040 95.880 93.210 ;
        RECT 96.050 93.040 96.080 93.210 ;
        RECT 96.690 93.210 97.640 93.240 ;
        RECT 93.600 91.580 93.930 92.360 ;
        RECT 95.130 92.280 96.080 93.040 ;
      LAYER li1 ;
        RECT 96.260 92.400 96.510 93.110 ;
      LAYER li1 ;
        RECT 96.690 93.040 96.720 93.210 ;
        RECT 96.890 93.040 97.080 93.210 ;
        RECT 97.250 93.040 97.440 93.210 ;
        RECT 97.610 93.040 97.640 93.210 ;
        RECT 98.250 93.210 99.200 93.240 ;
        RECT 96.690 92.580 97.640 93.040 ;
      LAYER li1 ;
        RECT 97.820 92.400 98.070 93.110 ;
        RECT 96.260 92.230 98.070 92.400 ;
      LAYER li1 ;
        RECT 98.250 93.040 98.280 93.210 ;
        RECT 98.450 93.040 98.640 93.210 ;
        RECT 98.810 93.040 99.000 93.210 ;
        RECT 99.170 93.040 99.200 93.210 ;
        RECT 100.010 93.210 101.620 93.240 ;
        RECT 98.250 92.360 99.200 93.040 ;
      LAYER li1 ;
        RECT 96.260 92.060 96.430 92.230 ;
      LAYER li1 ;
        RECT 99.380 92.180 99.710 93.110 ;
        RECT 100.010 93.040 100.060 93.210 ;
        RECT 100.230 93.040 100.500 93.210 ;
        RECT 100.670 93.040 100.940 93.210 ;
        RECT 101.110 93.040 101.350 93.210 ;
        RECT 101.520 93.040 101.620 93.210 ;
        RECT 100.010 92.760 101.620 93.040 ;
        RECT 94.140 90.920 94.470 91.910 ;
      LAYER li1 ;
        RECT 95.170 91.830 96.430 92.060 ;
      LAYER li1 ;
        RECT 98.470 92.050 99.710 92.180 ;
        RECT 96.610 92.010 99.710 92.050 ;
        RECT 96.610 91.880 98.640 92.010 ;
      LAYER li1 ;
        RECT 96.260 91.700 96.430 91.830 ;
        RECT 96.260 91.530 98.150 91.700 ;
      LAYER li1 ;
        RECT 93.370 90.050 94.820 90.920 ;
        RECT 93.370 89.880 93.620 90.050 ;
        RECT 93.790 89.880 93.980 90.050 ;
        RECT 94.150 89.880 94.420 90.050 ;
        RECT 94.590 89.880 94.820 90.050 ;
        RECT 93.370 89.850 94.820 89.880 ;
        RECT 95.130 90.100 96.080 91.430 ;
        RECT 95.130 89.930 95.160 90.100 ;
        RECT 95.330 89.930 95.520 90.100 ;
        RECT 95.690 89.930 95.880 90.100 ;
        RECT 96.050 89.930 96.080 90.100 ;
        RECT 95.130 89.850 96.080 89.930 ;
      LAYER li1 ;
        RECT 96.260 89.850 96.510 91.530 ;
      LAYER li1 ;
        RECT 96.690 90.100 97.640 91.350 ;
        RECT 96.690 89.930 96.720 90.100 ;
        RECT 96.890 89.930 97.080 90.100 ;
        RECT 97.250 89.930 97.440 90.100 ;
        RECT 97.610 89.930 97.640 90.100 ;
        RECT 96.690 89.850 97.640 89.930 ;
      LAYER li1 ;
        RECT 97.820 89.850 98.150 91.530 ;
        RECT 98.930 91.490 99.260 91.830 ;
      LAYER li1 ;
        RECT 98.330 90.100 99.280 91.310 ;
        RECT 98.330 89.930 98.360 90.100 ;
        RECT 98.530 89.930 98.720 90.100 ;
        RECT 98.890 89.930 99.080 90.100 ;
        RECT 99.250 89.930 99.280 90.100 ;
        RECT 98.330 89.850 99.280 89.930 ;
        RECT 99.460 89.850 99.710 92.010 ;
        RECT 100.320 92.360 101.620 92.760 ;
        RECT 101.850 93.210 102.800 93.240 ;
        RECT 101.850 93.040 101.880 93.210 ;
        RECT 102.050 93.040 102.240 93.210 ;
        RECT 102.410 93.040 102.600 93.210 ;
        RECT 102.770 93.040 102.800 93.210 ;
        RECT 103.410 93.210 104.360 93.240 ;
        RECT 100.320 91.580 100.650 92.360 ;
        RECT 101.850 92.280 102.800 93.040 ;
      LAYER li1 ;
        RECT 102.980 92.400 103.230 93.110 ;
      LAYER li1 ;
        RECT 103.410 93.040 103.440 93.210 ;
        RECT 103.610 93.040 103.800 93.210 ;
        RECT 103.970 93.040 104.160 93.210 ;
        RECT 104.330 93.040 104.360 93.210 ;
        RECT 104.970 93.210 105.920 93.240 ;
        RECT 103.410 92.580 104.360 93.040 ;
      LAYER li1 ;
        RECT 104.540 92.400 104.790 93.110 ;
        RECT 102.980 92.230 104.790 92.400 ;
      LAYER li1 ;
        RECT 104.970 93.040 105.000 93.210 ;
        RECT 105.170 93.040 105.360 93.210 ;
        RECT 105.530 93.040 105.720 93.210 ;
        RECT 105.890 93.040 105.920 93.210 ;
        RECT 106.730 93.210 108.340 93.240 ;
        RECT 109.120 93.210 110.010 93.240 ;
        RECT 112.010 93.210 113.620 93.240 ;
        RECT 104.970 92.360 105.920 93.040 ;
      LAYER li1 ;
        RECT 102.980 92.060 103.150 92.230 ;
      LAYER li1 ;
        RECT 106.100 92.180 106.430 93.110 ;
        RECT 106.730 93.040 106.780 93.210 ;
        RECT 106.950 93.040 107.220 93.210 ;
        RECT 107.390 93.040 107.660 93.210 ;
        RECT 107.830 93.040 108.070 93.210 ;
        RECT 108.240 93.040 108.340 93.210 ;
        RECT 106.730 92.760 108.340 93.040 ;
        RECT 100.860 90.920 101.190 91.910 ;
      LAYER li1 ;
        RECT 101.890 91.830 103.150 92.060 ;
      LAYER li1 ;
        RECT 105.190 92.050 106.430 92.180 ;
        RECT 103.330 92.010 106.430 92.050 ;
        RECT 103.330 91.880 105.360 92.010 ;
      LAYER li1 ;
        RECT 102.980 91.700 103.150 91.830 ;
        RECT 102.980 91.530 104.870 91.700 ;
      LAYER li1 ;
        RECT 100.090 90.050 101.540 90.920 ;
        RECT 100.090 89.880 100.340 90.050 ;
        RECT 100.510 89.880 100.700 90.050 ;
        RECT 100.870 89.880 101.140 90.050 ;
        RECT 101.310 89.880 101.540 90.050 ;
        RECT 100.090 89.850 101.540 89.880 ;
        RECT 101.850 90.100 102.800 91.430 ;
        RECT 101.850 89.930 101.880 90.100 ;
        RECT 102.050 89.930 102.240 90.100 ;
        RECT 102.410 89.930 102.600 90.100 ;
        RECT 102.770 89.930 102.800 90.100 ;
        RECT 101.850 89.850 102.800 89.930 ;
      LAYER li1 ;
        RECT 102.980 89.850 103.230 91.530 ;
      LAYER li1 ;
        RECT 103.410 90.100 104.360 91.350 ;
        RECT 103.410 89.930 103.440 90.100 ;
        RECT 103.610 89.930 103.800 90.100 ;
        RECT 103.970 89.930 104.160 90.100 ;
        RECT 104.330 89.930 104.360 90.100 ;
        RECT 103.410 89.850 104.360 89.930 ;
      LAYER li1 ;
        RECT 104.540 89.850 104.870 91.530 ;
        RECT 105.650 91.490 105.980 91.830 ;
      LAYER li1 ;
        RECT 105.050 90.100 106.000 91.310 ;
        RECT 105.050 89.930 105.080 90.100 ;
        RECT 105.250 89.930 105.440 90.100 ;
        RECT 105.610 89.930 105.800 90.100 ;
        RECT 105.970 89.930 106.000 90.100 ;
        RECT 105.050 89.850 106.000 89.930 ;
        RECT 106.180 89.850 106.430 92.010 ;
        RECT 107.040 92.360 108.340 92.760 ;
        RECT 108.610 92.500 108.940 93.110 ;
        RECT 109.290 93.040 109.480 93.210 ;
        RECT 109.650 93.040 109.840 93.210 ;
        RECT 109.120 92.680 110.010 93.040 ;
        RECT 110.190 92.500 110.520 93.110 ;
        RECT 107.040 91.580 107.370 92.360 ;
        RECT 108.610 92.330 110.520 92.500 ;
        RECT 108.610 92.280 108.940 92.330 ;
      LAYER li1 ;
        RECT 110.970 92.150 111.300 93.110 ;
      LAYER li1 ;
        RECT 112.010 93.040 112.060 93.210 ;
        RECT 112.230 93.040 112.500 93.210 ;
        RECT 112.670 93.040 112.940 93.210 ;
        RECT 113.110 93.040 113.350 93.210 ;
        RECT 113.520 93.040 113.620 93.210 ;
        RECT 112.010 92.760 113.620 93.040 ;
        RECT 107.580 90.920 107.910 91.910 ;
      LAYER li1 ;
        RECT 108.610 91.770 109.340 92.100 ;
        RECT 109.550 91.850 110.280 92.100 ;
        RECT 110.460 91.980 111.300 92.150 ;
      LAYER li1 ;
        RECT 112.320 92.360 113.620 92.760 ;
        RECT 113.850 93.210 114.440 93.240 ;
        RECT 113.850 93.040 113.880 93.210 ;
        RECT 114.050 93.040 114.240 93.210 ;
        RECT 114.410 93.040 114.440 93.210 ;
        RECT 115.370 93.210 116.980 93.240 ;
        RECT 117.670 93.210 118.920 93.240 ;
        RECT 119.690 93.210 121.300 93.240 ;
      LAYER li1 ;
        RECT 110.460 91.670 110.630 91.980 ;
        RECT 110.050 91.500 110.630 91.670 ;
      LAYER li1 ;
        RECT 106.810 90.050 108.260 90.920 ;
        RECT 106.810 89.880 107.060 90.050 ;
        RECT 107.230 89.880 107.420 90.050 ;
        RECT 107.590 89.880 107.860 90.050 ;
        RECT 108.030 89.880 108.260 90.050 ;
        RECT 106.810 89.850 108.260 89.880 ;
        RECT 108.570 90.100 109.520 91.430 ;
        RECT 108.570 89.930 108.600 90.100 ;
        RECT 108.770 89.930 108.960 90.100 ;
        RECT 109.130 89.930 109.320 90.100 ;
        RECT 109.490 89.930 109.520 90.100 ;
        RECT 108.570 89.850 109.520 89.930 ;
      LAYER li1 ;
        RECT 110.050 89.850 110.520 91.500 ;
        RECT 110.810 91.490 111.720 91.800 ;
      LAYER li1 ;
        RECT 112.320 91.580 112.650 92.360 ;
        RECT 113.850 92.280 114.440 93.040 ;
        RECT 110.700 90.100 111.650 91.310 ;
        RECT 112.860 90.920 113.190 91.910 ;
      LAYER li1 ;
        RECT 113.890 91.670 114.600 92.060 ;
        RECT 114.780 91.430 115.110 93.110 ;
      LAYER li1 ;
        RECT 115.370 93.040 115.420 93.210 ;
        RECT 115.590 93.040 115.860 93.210 ;
        RECT 116.030 93.040 116.300 93.210 ;
        RECT 116.470 93.040 116.710 93.210 ;
        RECT 116.880 93.040 116.980 93.210 ;
        RECT 115.370 92.760 116.980 93.040 ;
        RECT 115.680 92.360 116.980 92.760 ;
        RECT 115.680 91.580 116.010 92.360 ;
        RECT 110.700 89.930 110.730 90.100 ;
        RECT 110.900 89.930 111.090 90.100 ;
        RECT 111.260 89.930 111.450 90.100 ;
        RECT 111.620 89.930 111.650 90.100 ;
        RECT 110.700 89.850 111.650 89.930 ;
        RECT 112.090 90.050 113.540 90.920 ;
        RECT 112.090 89.880 112.340 90.050 ;
        RECT 112.510 89.880 112.700 90.050 ;
        RECT 112.870 89.880 113.140 90.050 ;
        RECT 113.310 89.880 113.540 90.050 ;
        RECT 112.090 89.850 113.540 89.880 ;
        RECT 113.850 90.100 114.440 91.430 ;
        RECT 113.850 89.930 113.880 90.100 ;
        RECT 114.050 89.930 114.240 90.100 ;
        RECT 114.410 89.930 114.440 90.100 ;
        RECT 113.850 89.850 114.440 89.930 ;
      LAYER li1 ;
        RECT 114.720 89.850 115.110 91.430 ;
      LAYER li1 ;
        RECT 116.220 90.920 116.550 91.910 ;
      LAYER li1 ;
        RECT 117.240 91.430 117.490 93.110 ;
      LAYER li1 ;
        RECT 117.840 93.040 118.030 93.210 ;
        RECT 118.200 93.040 118.390 93.210 ;
        RECT 118.560 93.040 118.750 93.210 ;
        RECT 117.670 92.670 118.920 93.040 ;
        RECT 119.100 92.490 119.350 93.110 ;
        RECT 119.690 93.040 119.740 93.210 ;
        RECT 119.910 93.040 120.180 93.210 ;
        RECT 120.350 93.040 120.620 93.210 ;
        RECT 120.790 93.040 121.030 93.210 ;
        RECT 121.200 93.040 121.300 93.210 ;
        RECT 119.690 92.760 121.300 93.040 ;
        RECT 117.800 92.320 119.350 92.490 ;
        RECT 117.800 91.860 118.130 92.320 ;
        RECT 115.450 90.050 116.900 90.920 ;
        RECT 115.450 89.880 115.700 90.050 ;
        RECT 115.870 89.880 116.060 90.050 ;
        RECT 116.230 89.880 116.500 90.050 ;
        RECT 116.670 89.880 116.900 90.050 ;
        RECT 115.450 89.850 116.900 89.880 ;
      LAYER li1 ;
        RECT 117.240 89.850 117.670 91.430 ;
      LAYER li1 ;
        RECT 117.850 90.100 118.410 91.430 ;
      LAYER li1 ;
        RECT 118.590 90.350 118.920 92.140 ;
      LAYER li1 ;
        RECT 119.100 90.600 119.350 92.320 ;
        RECT 120.000 92.360 121.300 92.760 ;
        RECT 121.530 93.210 122.480 93.240 ;
        RECT 121.530 93.040 121.560 93.210 ;
        RECT 121.730 93.040 121.920 93.210 ;
        RECT 122.090 93.040 122.280 93.210 ;
        RECT 122.450 93.040 122.480 93.210 ;
        RECT 123.090 93.210 124.040 93.240 ;
        RECT 120.000 91.580 120.330 92.360 ;
        RECT 121.530 92.280 122.480 93.040 ;
      LAYER li1 ;
        RECT 122.660 92.400 122.910 93.110 ;
      LAYER li1 ;
        RECT 123.090 93.040 123.120 93.210 ;
        RECT 123.290 93.040 123.480 93.210 ;
        RECT 123.650 93.040 123.840 93.210 ;
        RECT 124.010 93.040 124.040 93.210 ;
        RECT 124.650 93.210 125.600 93.240 ;
        RECT 123.090 92.580 124.040 93.040 ;
      LAYER li1 ;
        RECT 124.220 92.400 124.470 93.110 ;
        RECT 122.660 92.230 124.470 92.400 ;
      LAYER li1 ;
        RECT 124.650 93.040 124.680 93.210 ;
        RECT 124.850 93.040 125.040 93.210 ;
        RECT 125.210 93.040 125.400 93.210 ;
        RECT 125.570 93.040 125.600 93.210 ;
        RECT 126.820 93.220 129.550 93.250 ;
        RECT 124.650 92.360 125.600 93.040 ;
      LAYER li1 ;
        RECT 122.660 92.060 122.830 92.230 ;
      LAYER li1 ;
        RECT 125.780 92.180 126.110 93.110 ;
        RECT 126.820 93.050 126.990 93.220 ;
        RECT 127.160 93.050 127.430 93.220 ;
        RECT 127.600 93.050 127.840 93.220 ;
        RECT 128.010 93.050 128.270 93.220 ;
        RECT 128.440 93.050 128.710 93.220 ;
        RECT 128.880 93.050 129.120 93.220 ;
        RECT 129.290 93.050 129.550 93.220 ;
        RECT 126.820 92.250 129.550 93.050 ;
        RECT 130.660 93.220 133.390 93.250 ;
        RECT 130.660 93.050 130.830 93.220 ;
        RECT 131.000 93.050 131.270 93.220 ;
        RECT 131.440 93.050 131.680 93.220 ;
        RECT 131.850 93.050 132.110 93.220 ;
        RECT 132.280 93.050 132.550 93.220 ;
        RECT 132.720 93.050 132.960 93.220 ;
        RECT 133.130 93.050 133.390 93.220 ;
        RECT 130.660 92.250 133.390 93.050 ;
        RECT 134.500 93.220 137.230 93.250 ;
        RECT 134.500 93.050 134.670 93.220 ;
        RECT 134.840 93.050 135.110 93.220 ;
        RECT 135.280 93.050 135.520 93.220 ;
        RECT 135.690 93.050 135.950 93.220 ;
        RECT 136.120 93.050 136.390 93.220 ;
        RECT 136.560 93.050 136.800 93.220 ;
        RECT 136.970 93.050 137.230 93.220 ;
        RECT 134.500 92.250 137.230 93.050 ;
        RECT 138.340 93.220 141.070 93.250 ;
        RECT 138.340 93.050 138.510 93.220 ;
        RECT 138.680 93.050 138.950 93.220 ;
        RECT 139.120 93.050 139.360 93.220 ;
        RECT 139.530 93.050 139.790 93.220 ;
        RECT 139.960 93.050 140.230 93.220 ;
        RECT 140.400 93.050 140.640 93.220 ;
        RECT 140.810 93.050 141.070 93.220 ;
        RECT 138.340 92.250 141.070 93.050 ;
        RECT 120.540 90.920 120.870 91.910 ;
      LAYER li1 ;
        RECT 121.570 91.830 122.830 92.060 ;
      LAYER li1 ;
        RECT 124.870 92.050 126.110 92.180 ;
        RECT 123.010 92.010 126.110 92.050 ;
        RECT 123.010 91.880 125.040 92.010 ;
      LAYER li1 ;
        RECT 122.660 91.700 122.830 91.830 ;
        RECT 122.660 91.530 124.550 91.700 ;
      LAYER li1 ;
        RECT 117.850 89.930 117.860 90.100 ;
        RECT 118.030 89.930 118.220 90.100 ;
        RECT 118.390 89.930 118.410 90.100 ;
        RECT 117.850 89.850 118.410 89.930 ;
        RECT 119.770 90.050 121.220 90.920 ;
        RECT 119.770 89.880 120.020 90.050 ;
        RECT 120.190 89.880 120.380 90.050 ;
        RECT 120.550 89.880 120.820 90.050 ;
        RECT 120.990 89.880 121.220 90.050 ;
        RECT 119.770 89.850 121.220 89.880 ;
        RECT 121.530 90.100 122.480 91.430 ;
        RECT 121.530 89.930 121.560 90.100 ;
        RECT 121.730 89.930 121.920 90.100 ;
        RECT 122.090 89.930 122.280 90.100 ;
        RECT 122.450 89.930 122.480 90.100 ;
        RECT 121.530 89.850 122.480 89.930 ;
      LAYER li1 ;
        RECT 122.660 89.850 122.910 91.530 ;
      LAYER li1 ;
        RECT 123.090 90.100 124.040 91.350 ;
        RECT 123.090 89.930 123.120 90.100 ;
        RECT 123.290 89.930 123.480 90.100 ;
        RECT 123.650 89.930 123.840 90.100 ;
        RECT 124.010 89.930 124.040 90.100 ;
        RECT 123.090 89.850 124.040 89.930 ;
      LAYER li1 ;
        RECT 124.220 89.850 124.550 91.530 ;
        RECT 125.330 91.490 125.660 91.830 ;
      LAYER li1 ;
        RECT 124.730 90.100 125.680 91.310 ;
        RECT 124.730 89.930 124.760 90.100 ;
        RECT 124.930 89.930 125.120 90.100 ;
        RECT 125.290 89.930 125.480 90.100 ;
        RECT 125.650 89.930 125.680 90.100 ;
        RECT 124.730 89.850 125.680 89.930 ;
        RECT 125.860 89.850 126.110 92.010 ;
        RECT 126.980 91.580 127.310 92.250 ;
        RECT 127.710 90.930 128.040 91.910 ;
        RECT 128.260 91.580 128.590 92.250 ;
        RECT 128.990 90.930 129.320 91.910 ;
        RECT 130.820 91.580 131.150 92.250 ;
        RECT 131.550 90.930 131.880 91.910 ;
        RECT 132.100 91.580 132.430 92.250 ;
        RECT 132.830 90.930 133.160 91.910 ;
        RECT 134.660 91.580 134.990 92.250 ;
        RECT 135.390 90.930 135.720 91.910 ;
        RECT 135.940 91.580 136.270 92.250 ;
        RECT 136.670 90.930 137.000 91.910 ;
        RECT 138.500 91.580 138.830 92.250 ;
        RECT 139.230 90.930 139.560 91.910 ;
        RECT 139.780 91.580 140.110 92.250 ;
        RECT 140.510 90.930 140.840 91.910 ;
        RECT 126.740 90.050 129.480 90.930 ;
        RECT 126.740 89.880 126.950 90.050 ;
        RECT 127.120 89.880 127.390 90.050 ;
        RECT 127.560 89.880 127.800 90.050 ;
        RECT 127.970 89.880 128.230 90.050 ;
        RECT 128.400 89.880 128.670 90.050 ;
        RECT 128.840 89.880 129.080 90.050 ;
        RECT 129.250 89.880 129.480 90.050 ;
        RECT 126.740 89.860 129.480 89.880 ;
        RECT 130.580 90.050 133.320 90.930 ;
        RECT 130.580 89.880 130.790 90.050 ;
        RECT 130.960 89.880 131.230 90.050 ;
        RECT 131.400 89.880 131.640 90.050 ;
        RECT 131.810 89.880 132.070 90.050 ;
        RECT 132.240 89.880 132.510 90.050 ;
        RECT 132.680 89.880 132.920 90.050 ;
        RECT 133.090 89.880 133.320 90.050 ;
        RECT 130.580 89.860 133.320 89.880 ;
        RECT 134.420 90.050 137.160 90.930 ;
        RECT 134.420 89.880 134.630 90.050 ;
        RECT 134.800 89.880 135.070 90.050 ;
        RECT 135.240 89.880 135.480 90.050 ;
        RECT 135.650 89.880 135.910 90.050 ;
        RECT 136.080 89.880 136.350 90.050 ;
        RECT 136.520 89.880 136.760 90.050 ;
        RECT 136.930 89.880 137.160 90.050 ;
        RECT 134.420 89.860 137.160 89.880 ;
        RECT 138.260 90.050 141.000 90.930 ;
        RECT 138.260 89.880 138.470 90.050 ;
        RECT 138.640 89.880 138.910 90.050 ;
        RECT 139.080 89.880 139.320 90.050 ;
        RECT 139.490 89.880 139.750 90.050 ;
        RECT 139.920 89.880 140.190 90.050 ;
        RECT 140.360 89.880 140.600 90.050 ;
        RECT 140.770 89.880 141.000 90.050 ;
        RECT 138.260 89.860 141.000 89.880 ;
        RECT 5.760 89.450 5.920 89.630 ;
        RECT 6.090 89.450 6.400 89.630 ;
        RECT 6.570 89.450 6.880 89.630 ;
        RECT 7.050 89.450 7.360 89.630 ;
        RECT 7.530 89.450 7.840 89.630 ;
        RECT 8.010 89.450 8.320 89.630 ;
        RECT 8.490 89.450 8.800 89.630 ;
        RECT 8.970 89.450 9.280 89.630 ;
        RECT 9.450 89.450 9.760 89.630 ;
        RECT 9.930 89.450 10.240 89.630 ;
        RECT 10.410 89.450 10.720 89.630 ;
        RECT 10.890 89.450 11.200 89.630 ;
        RECT 11.370 89.450 11.680 89.630 ;
        RECT 11.850 89.450 12.160 89.630 ;
        RECT 12.330 89.620 12.640 89.630 ;
        RECT 12.810 89.620 13.120 89.630 ;
        RECT 12.330 89.450 12.480 89.620 ;
        RECT 12.960 89.450 13.120 89.620 ;
        RECT 13.290 89.450 13.600 89.630 ;
        RECT 13.770 89.450 14.080 89.630 ;
        RECT 14.250 89.450 14.560 89.630 ;
        RECT 14.730 89.450 15.040 89.630 ;
        RECT 15.210 89.450 15.520 89.630 ;
        RECT 15.690 89.450 16.000 89.630 ;
        RECT 16.170 89.450 16.480 89.630 ;
        RECT 16.650 89.450 16.960 89.630 ;
        RECT 17.130 89.450 17.440 89.630 ;
        RECT 17.610 89.450 17.920 89.630 ;
        RECT 18.090 89.450 18.400 89.630 ;
        RECT 18.570 89.450 18.880 89.630 ;
        RECT 19.050 89.450 19.360 89.630 ;
        RECT 19.530 89.450 19.840 89.630 ;
        RECT 20.010 89.460 20.160 89.630 ;
        RECT 20.640 89.460 20.800 89.630 ;
        RECT 20.010 89.450 20.320 89.460 ;
        RECT 20.490 89.450 20.800 89.460 ;
        RECT 20.970 89.450 21.280 89.630 ;
        RECT 21.450 89.450 21.760 89.630 ;
        RECT 21.930 89.450 22.240 89.630 ;
        RECT 22.410 89.450 22.720 89.630 ;
        RECT 22.890 89.450 23.200 89.630 ;
        RECT 23.370 89.450 23.680 89.630 ;
        RECT 23.850 89.450 24.160 89.630 ;
        RECT 24.330 89.450 24.640 89.630 ;
        RECT 24.810 89.450 25.120 89.630 ;
        RECT 25.290 89.450 25.600 89.630 ;
        RECT 25.770 89.450 26.080 89.630 ;
        RECT 26.250 89.450 26.560 89.630 ;
        RECT 26.730 89.450 27.040 89.630 ;
        RECT 27.210 89.450 27.520 89.630 ;
        RECT 27.690 89.450 28.000 89.630 ;
        RECT 28.170 89.450 28.480 89.630 ;
        RECT 28.650 89.450 28.960 89.630 ;
        RECT 29.130 89.450 29.440 89.630 ;
        RECT 29.610 89.450 29.920 89.630 ;
        RECT 30.090 89.450 30.400 89.630 ;
        RECT 30.570 89.450 30.880 89.630 ;
        RECT 31.050 89.450 31.360 89.630 ;
        RECT 31.530 89.450 31.840 89.630 ;
        RECT 32.010 89.450 32.320 89.630 ;
        RECT 32.490 89.450 32.800 89.630 ;
        RECT 32.970 89.450 33.280 89.630 ;
        RECT 33.450 89.450 33.760 89.630 ;
        RECT 33.930 89.450 34.240 89.630 ;
        RECT 34.410 89.450 34.720 89.630 ;
        RECT 34.890 89.450 35.200 89.630 ;
        RECT 35.370 89.450 35.680 89.630 ;
        RECT 35.850 89.450 36.160 89.630 ;
        RECT 36.330 89.450 36.640 89.630 ;
        RECT 36.810 89.450 37.120 89.630 ;
        RECT 37.290 89.450 37.600 89.630 ;
        RECT 37.770 89.450 38.080 89.630 ;
        RECT 38.250 89.450 38.560 89.630 ;
        RECT 38.730 89.450 39.040 89.630 ;
        RECT 39.210 89.450 39.520 89.630 ;
        RECT 39.690 89.450 40.000 89.630 ;
        RECT 40.170 89.450 40.480 89.630 ;
        RECT 40.650 89.450 40.960 89.630 ;
        RECT 41.130 89.450 41.440 89.630 ;
        RECT 41.610 89.450 41.920 89.630 ;
        RECT 42.090 89.450 42.400 89.630 ;
        RECT 42.570 89.450 42.880 89.630 ;
        RECT 43.050 89.450 43.360 89.630 ;
        RECT 43.530 89.450 43.840 89.630 ;
        RECT 44.010 89.450 44.320 89.630 ;
        RECT 44.490 89.450 44.800 89.630 ;
        RECT 44.970 89.450 45.280 89.630 ;
        RECT 45.450 89.450 45.760 89.630 ;
        RECT 45.930 89.450 46.240 89.630 ;
        RECT 46.410 89.450 46.720 89.630 ;
        RECT 46.890 89.450 47.200 89.630 ;
        RECT 47.370 89.450 47.680 89.630 ;
        RECT 47.850 89.450 48.160 89.630 ;
        RECT 48.330 89.450 48.640 89.630 ;
        RECT 48.810 89.450 49.120 89.630 ;
        RECT 49.290 89.450 49.600 89.630 ;
        RECT 49.770 89.450 50.080 89.630 ;
        RECT 50.250 89.450 50.560 89.630 ;
        RECT 50.730 89.450 51.040 89.630 ;
        RECT 51.210 89.450 51.520 89.630 ;
        RECT 51.690 89.450 52.000 89.630 ;
        RECT 52.170 89.450 52.480 89.630 ;
        RECT 52.650 89.450 52.960 89.630 ;
        RECT 53.130 89.450 53.440 89.630 ;
        RECT 53.610 89.450 53.920 89.630 ;
        RECT 54.090 89.450 54.400 89.630 ;
        RECT 54.570 89.450 54.880 89.630 ;
        RECT 55.050 89.450 55.360 89.630 ;
        RECT 55.530 89.450 55.840 89.630 ;
        RECT 56.010 89.620 56.320 89.630 ;
        RECT 56.490 89.620 56.800 89.630 ;
        RECT 56.010 89.450 56.160 89.620 ;
        RECT 56.640 89.450 56.800 89.620 ;
        RECT 56.970 89.450 57.280 89.630 ;
        RECT 57.450 89.450 57.760 89.630 ;
        RECT 57.930 89.450 58.240 89.630 ;
        RECT 58.410 89.450 58.720 89.630 ;
        RECT 58.890 89.450 59.200 89.630 ;
        RECT 59.370 89.450 59.680 89.630 ;
        RECT 59.850 89.450 60.160 89.630 ;
        RECT 60.330 89.450 60.640 89.630 ;
        RECT 60.810 89.450 61.120 89.630 ;
        RECT 61.290 89.450 61.600 89.630 ;
        RECT 61.770 89.450 62.080 89.630 ;
        RECT 62.250 89.450 62.560 89.630 ;
        RECT 62.730 89.450 63.040 89.630 ;
        RECT 63.210 89.450 63.520 89.630 ;
        RECT 63.690 89.450 64.000 89.630 ;
        RECT 64.170 89.450 64.480 89.630 ;
        RECT 64.650 89.450 64.960 89.630 ;
        RECT 65.130 89.450 65.440 89.630 ;
        RECT 65.610 89.450 65.920 89.630 ;
        RECT 66.090 89.450 66.400 89.630 ;
        RECT 66.570 89.450 66.880 89.630 ;
        RECT 67.050 89.450 67.360 89.630 ;
        RECT 67.530 89.450 67.840 89.630 ;
        RECT 68.010 89.460 68.160 89.630 ;
        RECT 68.640 89.460 68.800 89.630 ;
        RECT 68.010 89.450 68.320 89.460 ;
        RECT 68.490 89.450 68.800 89.460 ;
        RECT 68.970 89.450 69.280 89.630 ;
        RECT 69.450 89.450 69.760 89.630 ;
        RECT 69.930 89.450 70.240 89.630 ;
        RECT 70.410 89.450 70.720 89.630 ;
        RECT 70.890 89.450 71.200 89.630 ;
        RECT 71.370 89.450 71.680 89.630 ;
        RECT 71.850 89.450 72.160 89.630 ;
        RECT 72.330 89.450 72.640 89.630 ;
        RECT 72.810 89.450 73.120 89.630 ;
        RECT 73.290 89.450 73.600 89.630 ;
        RECT 73.770 89.450 74.080 89.630 ;
        RECT 74.250 89.450 74.560 89.630 ;
        RECT 74.730 89.450 75.040 89.630 ;
        RECT 75.210 89.450 75.520 89.630 ;
        RECT 75.690 89.450 76.000 89.630 ;
        RECT 76.170 89.450 76.480 89.630 ;
        RECT 76.650 89.450 76.960 89.630 ;
        RECT 77.130 89.450 77.440 89.630 ;
        RECT 77.610 89.450 77.920 89.630 ;
        RECT 78.090 89.450 78.400 89.630 ;
        RECT 78.570 89.450 78.880 89.630 ;
        RECT 79.050 89.450 79.360 89.630 ;
        RECT 79.530 89.450 79.840 89.630 ;
        RECT 80.010 89.450 80.320 89.630 ;
        RECT 80.490 89.450 80.800 89.630 ;
        RECT 80.970 89.450 81.280 89.630 ;
        RECT 81.450 89.450 81.760 89.630 ;
        RECT 81.930 89.450 82.240 89.630 ;
        RECT 82.410 89.450 82.720 89.630 ;
        RECT 82.890 89.450 83.200 89.630 ;
        RECT 83.370 89.450 83.680 89.630 ;
        RECT 83.850 89.450 84.160 89.630 ;
        RECT 84.330 89.450 84.640 89.630 ;
        RECT 84.810 89.450 85.120 89.630 ;
        RECT 85.290 89.450 85.600 89.630 ;
        RECT 85.770 89.450 86.080 89.630 ;
        RECT 86.250 89.450 86.560 89.630 ;
        RECT 86.730 89.450 87.040 89.630 ;
        RECT 87.210 89.450 87.520 89.630 ;
        RECT 87.690 89.450 88.000 89.630 ;
        RECT 88.170 89.450 88.480 89.630 ;
        RECT 88.650 89.450 88.960 89.630 ;
        RECT 89.130 89.450 89.440 89.630 ;
        RECT 89.610 89.450 89.920 89.630 ;
        RECT 90.090 89.450 90.400 89.630 ;
        RECT 90.570 89.450 90.880 89.630 ;
        RECT 91.050 89.450 91.360 89.630 ;
        RECT 91.530 89.450 91.840 89.630 ;
        RECT 92.010 89.450 92.320 89.630 ;
        RECT 92.490 89.450 92.800 89.630 ;
        RECT 92.970 89.450 93.280 89.630 ;
        RECT 93.450 89.450 93.760 89.630 ;
        RECT 93.930 89.450 94.240 89.630 ;
        RECT 94.410 89.450 94.720 89.630 ;
        RECT 94.890 89.450 95.200 89.630 ;
        RECT 95.370 89.450 95.680 89.630 ;
        RECT 95.850 89.450 96.160 89.630 ;
        RECT 96.330 89.450 96.640 89.630 ;
        RECT 96.810 89.450 97.120 89.630 ;
        RECT 97.290 89.450 97.600 89.630 ;
        RECT 97.770 89.450 98.080 89.630 ;
        RECT 98.250 89.450 98.560 89.630 ;
        RECT 98.730 89.450 99.040 89.630 ;
        RECT 99.210 89.450 99.520 89.630 ;
        RECT 99.690 89.450 100.000 89.630 ;
        RECT 100.170 89.450 100.480 89.630 ;
        RECT 100.650 89.450 100.960 89.630 ;
        RECT 101.130 89.460 101.280 89.630 ;
        RECT 101.760 89.460 101.920 89.630 ;
        RECT 101.130 89.450 101.440 89.460 ;
        RECT 101.610 89.450 101.920 89.460 ;
        RECT 102.090 89.450 102.400 89.630 ;
        RECT 102.570 89.450 102.880 89.630 ;
        RECT 103.050 89.450 103.360 89.630 ;
        RECT 103.530 89.450 103.840 89.630 ;
        RECT 104.010 89.450 104.320 89.630 ;
        RECT 104.490 89.450 104.800 89.630 ;
        RECT 104.970 89.450 105.280 89.630 ;
        RECT 105.450 89.450 105.760 89.630 ;
        RECT 105.930 89.450 106.240 89.630 ;
        RECT 106.410 89.450 106.720 89.630 ;
        RECT 106.890 89.450 107.200 89.630 ;
        RECT 107.370 89.450 107.680 89.630 ;
        RECT 107.850 89.450 108.160 89.630 ;
        RECT 108.330 89.450 108.640 89.630 ;
        RECT 108.810 89.450 109.120 89.630 ;
        RECT 109.290 89.450 109.600 89.630 ;
        RECT 109.770 89.450 110.080 89.630 ;
        RECT 110.250 89.450 110.560 89.630 ;
        RECT 110.730 89.450 111.040 89.630 ;
        RECT 111.210 89.450 111.520 89.630 ;
        RECT 111.690 89.450 112.000 89.630 ;
        RECT 112.170 89.450 112.480 89.630 ;
        RECT 112.650 89.450 112.960 89.630 ;
        RECT 113.130 89.450 113.440 89.630 ;
        RECT 113.610 89.450 113.920 89.630 ;
        RECT 114.090 89.450 114.400 89.630 ;
        RECT 114.570 89.450 114.880 89.630 ;
        RECT 115.050 89.450 115.360 89.630 ;
        RECT 115.530 89.450 115.840 89.630 ;
        RECT 116.010 89.450 116.320 89.630 ;
        RECT 116.490 89.450 116.800 89.630 ;
        RECT 116.970 89.450 117.280 89.630 ;
        RECT 117.450 89.620 117.600 89.630 ;
        RECT 118.080 89.620 118.240 89.630 ;
        RECT 117.450 89.450 117.760 89.620 ;
        RECT 117.930 89.450 118.240 89.620 ;
        RECT 118.410 89.450 118.720 89.630 ;
        RECT 118.890 89.450 119.200 89.630 ;
        RECT 119.370 89.450 119.680 89.630 ;
        RECT 119.850 89.450 120.160 89.630 ;
        RECT 120.330 89.450 120.640 89.630 ;
        RECT 120.810 89.450 121.120 89.630 ;
        RECT 121.290 89.450 121.600 89.630 ;
        RECT 121.770 89.450 122.080 89.630 ;
        RECT 122.250 89.450 122.560 89.630 ;
        RECT 122.730 89.450 123.040 89.630 ;
        RECT 123.210 89.450 123.520 89.630 ;
        RECT 123.690 89.450 124.000 89.630 ;
        RECT 124.170 89.450 124.480 89.630 ;
        RECT 124.650 89.450 124.960 89.630 ;
        RECT 125.130 89.450 125.440 89.630 ;
        RECT 125.610 89.450 125.920 89.630 ;
        RECT 126.090 89.450 126.400 89.630 ;
        RECT 126.570 89.450 126.880 89.630 ;
        RECT 127.050 89.450 127.360 89.630 ;
        RECT 127.530 89.450 127.840 89.630 ;
        RECT 128.010 89.450 128.320 89.630 ;
        RECT 128.490 89.450 128.800 89.630 ;
        RECT 128.970 89.450 129.280 89.630 ;
        RECT 129.450 89.450 129.760 89.630 ;
        RECT 129.930 89.450 130.240 89.630 ;
        RECT 130.410 89.450 130.720 89.630 ;
        RECT 130.890 89.450 131.200 89.630 ;
        RECT 131.370 89.450 131.680 89.630 ;
        RECT 131.850 89.450 132.160 89.630 ;
        RECT 132.330 89.450 132.640 89.630 ;
        RECT 132.810 89.450 133.120 89.630 ;
        RECT 133.290 89.450 133.600 89.630 ;
        RECT 133.770 89.460 133.920 89.630 ;
        RECT 134.400 89.460 134.560 89.630 ;
        RECT 133.770 89.450 134.080 89.460 ;
        RECT 134.250 89.450 134.560 89.460 ;
        RECT 134.730 89.450 135.040 89.630 ;
        RECT 135.210 89.450 135.520 89.630 ;
        RECT 135.690 89.450 136.000 89.630 ;
        RECT 136.170 89.450 136.480 89.630 ;
        RECT 136.650 89.450 136.960 89.630 ;
        RECT 137.130 89.450 137.440 89.630 ;
        RECT 137.610 89.450 137.920 89.630 ;
        RECT 138.090 89.450 138.400 89.630 ;
        RECT 138.570 89.450 138.880 89.630 ;
        RECT 139.050 89.450 139.360 89.630 ;
        RECT 139.530 89.450 139.840 89.630 ;
        RECT 140.010 89.450 140.320 89.630 ;
        RECT 140.490 89.450 140.800 89.630 ;
        RECT 140.970 89.450 141.280 89.630 ;
        RECT 141.450 89.450 141.600 89.630 ;
        RECT 6.260 89.200 9.000 89.220 ;
        RECT 6.260 89.030 6.470 89.200 ;
        RECT 6.640 89.030 6.910 89.200 ;
        RECT 7.080 89.030 7.320 89.200 ;
        RECT 7.490 89.030 7.750 89.200 ;
        RECT 7.920 89.030 8.190 89.200 ;
        RECT 8.360 89.030 8.600 89.200 ;
        RECT 8.770 89.030 9.000 89.200 ;
        RECT 6.260 88.150 9.000 89.030 ;
        RECT 10.100 89.200 12.840 89.220 ;
        RECT 10.100 89.030 10.310 89.200 ;
        RECT 10.480 89.030 10.750 89.200 ;
        RECT 10.920 89.030 11.160 89.200 ;
        RECT 11.330 89.030 11.590 89.200 ;
        RECT 11.760 89.030 12.030 89.200 ;
        RECT 12.200 89.030 12.440 89.200 ;
        RECT 12.610 89.030 12.840 89.200 ;
        RECT 10.100 88.150 12.840 89.030 ;
        RECT 13.940 89.200 16.680 89.220 ;
        RECT 13.940 89.030 14.150 89.200 ;
        RECT 14.320 89.030 14.590 89.200 ;
        RECT 14.760 89.030 15.000 89.200 ;
        RECT 15.170 89.030 15.430 89.200 ;
        RECT 15.600 89.030 15.870 89.200 ;
        RECT 16.040 89.030 16.280 89.200 ;
        RECT 16.450 89.030 16.680 89.200 ;
        RECT 13.940 88.150 16.680 89.030 ;
        RECT 17.530 89.200 18.980 89.230 ;
        RECT 17.530 89.030 17.780 89.200 ;
        RECT 17.950 89.030 18.140 89.200 ;
        RECT 18.310 89.030 18.580 89.200 ;
        RECT 18.750 89.030 18.980 89.200 ;
        RECT 17.530 88.160 18.980 89.030 ;
        RECT 20.730 89.150 21.320 89.230 ;
        RECT 20.730 88.980 20.760 89.150 ;
        RECT 20.930 88.980 21.120 89.150 ;
        RECT 21.290 88.980 21.320 89.150 ;
        RECT 6.500 86.830 6.830 87.500 ;
        RECT 7.230 87.170 7.560 88.150 ;
        RECT 7.780 86.830 8.110 87.500 ;
        RECT 8.510 87.170 8.840 88.150 ;
        RECT 10.340 86.830 10.670 87.500 ;
        RECT 11.070 87.170 11.400 88.150 ;
        RECT 11.620 86.830 11.950 87.500 ;
        RECT 12.350 87.170 12.680 88.150 ;
        RECT 14.180 86.830 14.510 87.500 ;
        RECT 14.910 87.170 15.240 88.150 ;
        RECT 15.460 86.830 15.790 87.500 ;
        RECT 16.190 87.170 16.520 88.150 ;
        RECT 6.340 85.830 9.070 86.830 ;
        RECT 10.180 85.830 12.910 86.830 ;
        RECT 14.020 85.830 16.750 86.830 ;
        RECT 17.760 86.720 18.090 87.500 ;
        RECT 18.300 87.170 18.630 88.160 ;
        RECT 20.730 87.650 21.320 88.980 ;
      LAYER li1 ;
        RECT 21.600 87.650 21.990 89.230 ;
      LAYER li1 ;
        RECT 22.330 89.200 23.780 89.230 ;
        RECT 22.330 89.030 22.580 89.200 ;
        RECT 22.750 89.030 22.940 89.200 ;
        RECT 23.110 89.030 23.380 89.200 ;
        RECT 23.550 89.030 23.780 89.200 ;
        RECT 22.330 88.160 23.780 89.030 ;
        RECT 24.090 89.150 24.680 89.230 ;
        RECT 24.090 88.980 24.120 89.150 ;
        RECT 24.290 88.980 24.480 89.150 ;
        RECT 24.650 88.980 24.680 89.150 ;
      LAYER li1 ;
        RECT 20.770 87.020 21.480 87.410 ;
      LAYER li1 ;
        RECT 17.760 86.320 19.060 86.720 ;
        RECT 17.450 85.840 19.060 86.320 ;
        RECT 20.730 85.840 21.320 86.800 ;
      LAYER li1 ;
        RECT 21.660 85.970 21.990 87.650 ;
      LAYER li1 ;
        RECT 22.560 86.720 22.890 87.500 ;
        RECT 23.100 87.170 23.430 88.160 ;
        RECT 24.090 87.650 24.680 88.980 ;
      LAYER li1 ;
        RECT 24.960 87.650 25.350 89.230 ;
      LAYER li1 ;
        RECT 25.690 89.200 27.140 89.230 ;
        RECT 25.690 89.030 25.940 89.200 ;
        RECT 26.110 89.030 26.300 89.200 ;
        RECT 26.470 89.030 26.740 89.200 ;
        RECT 26.910 89.030 27.140 89.200 ;
        RECT 25.690 88.160 27.140 89.030 ;
      LAYER li1 ;
        RECT 24.130 87.020 24.840 87.410 ;
      LAYER li1 ;
        RECT 22.560 86.320 23.860 86.720 ;
        RECT 22.250 85.840 23.860 86.320 ;
        RECT 24.090 85.840 24.680 86.800 ;
      LAYER li1 ;
        RECT 25.020 85.970 25.350 87.650 ;
      LAYER li1 ;
        RECT 25.920 86.720 26.250 87.500 ;
        RECT 26.460 87.170 26.790 88.160 ;
      LAYER li1 ;
        RECT 27.480 87.650 27.910 89.230 ;
      LAYER li1 ;
        RECT 28.090 89.150 28.650 89.230 ;
        RECT 28.090 88.980 28.100 89.150 ;
        RECT 28.270 88.980 28.460 89.150 ;
        RECT 28.630 88.980 28.650 89.150 ;
        RECT 28.090 87.650 28.650 88.980 ;
        RECT 30.010 89.200 31.460 89.230 ;
        RECT 30.010 89.030 30.260 89.200 ;
        RECT 30.430 89.030 30.620 89.200 ;
        RECT 30.790 89.030 31.060 89.200 ;
        RECT 31.230 89.030 31.460 89.200 ;
        RECT 25.920 86.320 27.220 86.720 ;
        RECT 25.610 85.840 27.220 86.320 ;
      LAYER li1 ;
        RECT 27.480 85.970 27.730 87.650 ;
      LAYER li1 ;
        RECT 28.040 86.760 28.370 87.220 ;
      LAYER li1 ;
        RECT 28.830 86.940 29.160 88.730 ;
      LAYER li1 ;
        RECT 29.340 86.760 29.590 88.480 ;
        RECT 30.010 88.160 31.460 89.030 ;
        RECT 31.770 89.150 32.720 89.230 ;
        RECT 31.770 88.980 31.800 89.150 ;
        RECT 31.970 88.980 32.160 89.150 ;
        RECT 32.330 88.980 32.520 89.150 ;
        RECT 32.690 88.980 32.720 89.150 ;
        RECT 28.040 86.590 29.590 86.760 ;
        RECT 27.910 85.840 29.160 86.410 ;
        RECT 29.340 85.970 29.590 86.590 ;
        RECT 30.240 86.720 30.570 87.500 ;
        RECT 30.780 87.170 31.110 88.160 ;
        RECT 31.770 87.650 32.720 88.980 ;
      LAYER li1 ;
        RECT 32.900 87.550 33.150 89.230 ;
      LAYER li1 ;
        RECT 33.330 89.150 34.280 89.230 ;
        RECT 33.330 88.980 33.360 89.150 ;
        RECT 33.530 88.980 33.720 89.150 ;
        RECT 33.890 88.980 34.080 89.150 ;
        RECT 34.250 88.980 34.280 89.150 ;
        RECT 33.330 87.730 34.280 88.980 ;
      LAYER li1 ;
        RECT 34.460 87.550 34.790 89.230 ;
      LAYER li1 ;
        RECT 34.970 89.150 35.920 89.230 ;
        RECT 34.970 88.980 35.000 89.150 ;
        RECT 35.170 88.980 35.360 89.150 ;
        RECT 35.530 88.980 35.720 89.150 ;
        RECT 35.890 88.980 35.920 89.150 ;
        RECT 34.970 87.770 35.920 88.980 ;
      LAYER li1 ;
        RECT 32.900 87.380 34.790 87.550 ;
        RECT 32.900 87.250 33.070 87.380 ;
        RECT 35.570 87.250 35.900 87.590 ;
        RECT 31.810 87.020 33.070 87.250 ;
      LAYER li1 ;
        RECT 33.250 87.070 35.280 87.200 ;
        RECT 36.100 87.070 36.350 89.230 ;
        RECT 36.730 89.200 38.180 89.230 ;
        RECT 36.730 89.030 36.980 89.200 ;
        RECT 37.150 89.030 37.340 89.200 ;
        RECT 37.510 89.030 37.780 89.200 ;
        RECT 37.950 89.030 38.180 89.200 ;
        RECT 36.730 88.160 38.180 89.030 ;
        RECT 38.490 89.150 39.440 89.230 ;
        RECT 38.490 88.980 38.520 89.150 ;
        RECT 38.690 88.980 38.880 89.150 ;
        RECT 39.050 88.980 39.240 89.150 ;
        RECT 39.410 88.980 39.440 89.150 ;
        RECT 33.250 87.030 36.350 87.070 ;
      LAYER li1 ;
        RECT 32.900 86.850 33.070 87.020 ;
      LAYER li1 ;
        RECT 35.110 86.900 36.350 87.030 ;
        RECT 30.240 86.320 31.540 86.720 ;
        RECT 29.930 85.840 31.540 86.320 ;
        RECT 31.770 85.840 32.720 86.800 ;
      LAYER li1 ;
        RECT 32.900 86.680 34.710 86.850 ;
        RECT 32.900 85.970 33.150 86.680 ;
      LAYER li1 ;
        RECT 33.330 85.840 34.280 86.500 ;
      LAYER li1 ;
        RECT 34.460 85.970 34.710 86.680 ;
      LAYER li1 ;
        RECT 34.890 85.840 35.840 86.720 ;
        RECT 36.020 85.970 36.350 86.900 ;
        RECT 36.960 86.720 37.290 87.500 ;
        RECT 37.500 87.170 37.830 88.160 ;
        RECT 38.490 87.650 39.440 88.980 ;
      LAYER li1 ;
        RECT 39.620 87.550 39.870 89.230 ;
      LAYER li1 ;
        RECT 40.050 89.150 41.000 89.230 ;
        RECT 40.050 88.980 40.080 89.150 ;
        RECT 40.250 88.980 40.440 89.150 ;
        RECT 40.610 88.980 40.800 89.150 ;
        RECT 40.970 88.980 41.000 89.150 ;
        RECT 40.050 87.730 41.000 88.980 ;
      LAYER li1 ;
        RECT 41.180 87.550 41.510 89.230 ;
      LAYER li1 ;
        RECT 41.690 89.150 42.640 89.230 ;
        RECT 41.690 88.980 41.720 89.150 ;
        RECT 41.890 88.980 42.080 89.150 ;
        RECT 42.250 88.980 42.440 89.150 ;
        RECT 42.610 88.980 42.640 89.150 ;
        RECT 41.690 87.770 42.640 88.980 ;
      LAYER li1 ;
        RECT 39.620 87.380 41.510 87.550 ;
        RECT 39.620 87.250 39.790 87.380 ;
        RECT 42.290 87.250 42.620 87.590 ;
        RECT 38.530 87.020 39.790 87.250 ;
      LAYER li1 ;
        RECT 39.970 87.070 42.000 87.200 ;
        RECT 42.820 87.070 43.070 89.230 ;
        RECT 43.450 89.200 44.900 89.230 ;
        RECT 43.450 89.030 43.700 89.200 ;
        RECT 43.870 89.030 44.060 89.200 ;
        RECT 44.230 89.030 44.500 89.200 ;
        RECT 44.670 89.030 44.900 89.200 ;
        RECT 43.450 88.160 44.900 89.030 ;
        RECT 45.210 89.150 46.160 89.230 ;
        RECT 45.210 88.980 45.240 89.150 ;
        RECT 45.410 88.980 45.600 89.150 ;
        RECT 45.770 88.980 45.960 89.150 ;
        RECT 46.130 88.980 46.160 89.150 ;
        RECT 39.970 87.030 43.070 87.070 ;
      LAYER li1 ;
        RECT 39.620 86.850 39.790 87.020 ;
      LAYER li1 ;
        RECT 41.830 86.900 43.070 87.030 ;
        RECT 36.960 86.320 38.260 86.720 ;
        RECT 36.650 85.840 38.260 86.320 ;
        RECT 38.490 85.840 39.440 86.800 ;
      LAYER li1 ;
        RECT 39.620 86.680 41.430 86.850 ;
        RECT 39.620 85.970 39.870 86.680 ;
      LAYER li1 ;
        RECT 40.050 85.840 41.000 86.500 ;
      LAYER li1 ;
        RECT 41.180 85.970 41.430 86.680 ;
      LAYER li1 ;
        RECT 41.610 85.840 42.560 86.720 ;
        RECT 42.740 85.970 43.070 86.900 ;
        RECT 43.680 86.720 44.010 87.500 ;
        RECT 44.220 87.170 44.550 88.160 ;
        RECT 45.210 87.650 46.160 88.980 ;
      LAYER li1 ;
        RECT 46.340 87.550 46.590 89.230 ;
      LAYER li1 ;
        RECT 46.770 89.150 47.720 89.230 ;
        RECT 46.770 88.980 46.800 89.150 ;
        RECT 46.970 88.980 47.160 89.150 ;
        RECT 47.330 88.980 47.520 89.150 ;
        RECT 47.690 88.980 47.720 89.150 ;
        RECT 46.770 87.730 47.720 88.980 ;
      LAYER li1 ;
        RECT 47.900 87.550 48.230 89.230 ;
      LAYER li1 ;
        RECT 48.410 89.150 49.360 89.230 ;
        RECT 48.410 88.980 48.440 89.150 ;
        RECT 48.610 88.980 48.800 89.150 ;
        RECT 48.970 88.980 49.160 89.150 ;
        RECT 49.330 88.980 49.360 89.150 ;
        RECT 48.410 87.770 49.360 88.980 ;
      LAYER li1 ;
        RECT 46.340 87.380 48.230 87.550 ;
        RECT 46.340 87.250 46.510 87.380 ;
        RECT 49.010 87.250 49.340 87.590 ;
        RECT 45.250 87.020 46.510 87.250 ;
      LAYER li1 ;
        RECT 46.690 87.070 48.720 87.200 ;
        RECT 49.540 87.070 49.790 89.230 ;
        RECT 50.170 89.200 51.620 89.230 ;
        RECT 50.170 89.030 50.420 89.200 ;
        RECT 50.590 89.030 50.780 89.200 ;
        RECT 50.950 89.030 51.220 89.200 ;
        RECT 51.390 89.030 51.620 89.200 ;
        RECT 50.170 88.160 51.620 89.030 ;
        RECT 51.930 89.150 53.190 89.230 ;
        RECT 51.930 88.980 51.940 89.150 ;
        RECT 52.110 88.980 52.300 89.150 ;
        RECT 52.470 88.980 52.660 89.150 ;
        RECT 52.830 88.980 53.020 89.150 ;
        RECT 46.690 87.030 49.790 87.070 ;
      LAYER li1 ;
        RECT 46.340 86.850 46.510 87.020 ;
      LAYER li1 ;
        RECT 48.550 86.900 49.790 87.030 ;
        RECT 43.680 86.320 44.980 86.720 ;
        RECT 43.370 85.840 44.980 86.320 ;
        RECT 45.210 85.840 46.160 86.800 ;
      LAYER li1 ;
        RECT 46.340 86.680 48.150 86.850 ;
        RECT 46.340 85.970 46.590 86.680 ;
      LAYER li1 ;
        RECT 46.770 85.840 47.720 86.500 ;
      LAYER li1 ;
        RECT 47.900 85.970 48.150 86.680 ;
      LAYER li1 ;
        RECT 48.330 85.840 49.280 86.720 ;
        RECT 49.460 85.970 49.790 86.900 ;
        RECT 50.400 86.720 50.730 87.500 ;
        RECT 50.940 87.170 51.270 88.160 ;
        RECT 51.930 87.750 53.190 88.980 ;
      LAYER li1 ;
        RECT 53.720 88.730 53.890 89.230 ;
        RECT 53.370 87.650 53.890 88.730 ;
      LAYER li1 ;
        RECT 54.150 89.150 55.460 89.230 ;
        RECT 54.150 88.980 54.180 89.150 ;
        RECT 54.350 88.980 54.540 89.150 ;
        RECT 54.710 88.980 54.900 89.150 ;
        RECT 55.070 88.980 55.260 89.150 ;
        RECT 55.430 88.980 55.460 89.150 ;
        RECT 54.150 87.770 55.460 88.980 ;
        RECT 55.930 89.200 57.380 89.230 ;
        RECT 55.930 89.030 56.180 89.200 ;
        RECT 56.350 89.030 56.540 89.200 ;
        RECT 56.710 89.030 56.980 89.200 ;
        RECT 57.150 89.030 57.380 89.200 ;
        RECT 55.930 88.160 57.380 89.030 ;
      LAYER li1 ;
        RECT 53.370 87.570 53.640 87.650 ;
        RECT 52.580 87.400 53.640 87.570 ;
        RECT 51.970 87.010 52.390 87.340 ;
        RECT 52.580 86.830 52.750 87.400 ;
        RECT 54.090 87.280 54.600 87.590 ;
        RECT 54.850 87.280 55.560 87.590 ;
        RECT 52.930 87.010 53.440 87.220 ;
      LAYER li1 ;
        RECT 53.640 86.930 55.510 87.100 ;
        RECT 50.400 86.320 51.700 86.720 ;
        RECT 50.090 85.840 51.700 86.320 ;
        RECT 52.000 85.910 52.330 86.830 ;
      LAYER li1 ;
        RECT 52.580 86.090 53.110 86.830 ;
      LAYER li1 ;
        RECT 53.640 85.910 53.810 86.930 ;
        RECT 52.000 85.740 53.810 85.910 ;
        RECT 53.990 85.840 55.090 86.750 ;
        RECT 55.260 86.000 55.510 86.930 ;
        RECT 56.160 86.720 56.490 87.500 ;
        RECT 56.700 87.170 57.030 88.160 ;
      LAYER li1 ;
        RECT 57.730 87.450 58.200 89.230 ;
      LAYER li1 ;
        RECT 58.380 89.150 59.630 89.230 ;
        RECT 58.550 88.980 58.740 89.150 ;
        RECT 58.910 88.980 59.100 89.150 ;
        RECT 59.270 88.980 59.460 89.150 ;
        RECT 58.380 87.770 59.630 88.980 ;
        RECT 56.160 86.320 57.460 86.720 ;
        RECT 55.850 85.840 57.460 86.320 ;
      LAYER li1 ;
        RECT 57.730 86.000 57.980 87.450 ;
        RECT 58.690 87.280 59.600 87.590 ;
      LAYER li1 ;
        RECT 58.150 87.100 58.440 87.270 ;
        RECT 59.810 87.100 59.980 89.230 ;
        RECT 60.570 89.150 61.830 89.230 ;
        RECT 60.740 88.980 60.930 89.150 ;
        RECT 61.100 88.980 61.290 89.150 ;
        RECT 61.460 88.980 61.650 89.150 ;
        RECT 61.820 88.980 61.830 89.150 ;
      LAYER li1 ;
        RECT 60.160 87.220 60.390 88.730 ;
      LAYER li1 ;
        RECT 60.570 87.650 61.830 88.980 ;
        RECT 62.170 89.200 63.620 89.230 ;
        RECT 62.170 89.030 62.420 89.200 ;
        RECT 62.590 89.030 62.780 89.200 ;
        RECT 62.950 89.030 63.220 89.200 ;
        RECT 63.390 89.030 63.620 89.200 ;
        RECT 62.170 88.160 63.620 89.030 ;
        RECT 58.150 86.930 59.980 87.100 ;
      LAYER li1 ;
        RECT 60.150 87.050 60.390 87.220 ;
        RECT 60.160 87.020 60.390 87.050 ;
        RECT 60.610 86.980 61.800 87.310 ;
      LAYER li1 ;
        RECT 58.150 85.840 58.920 86.750 ;
        RECT 59.100 85.970 59.430 86.930 ;
        RECT 61.460 86.750 61.790 86.800 ;
        RECT 59.880 86.580 61.790 86.750 ;
        RECT 59.880 85.970 60.210 86.580 ;
        RECT 60.390 85.840 61.280 86.400 ;
        RECT 61.460 85.970 61.790 86.580 ;
        RECT 62.400 86.720 62.730 87.500 ;
        RECT 62.940 87.170 63.270 88.160 ;
      LAYER li1 ;
        RECT 63.960 87.650 64.390 89.230 ;
      LAYER li1 ;
        RECT 64.570 89.150 65.130 89.230 ;
        RECT 64.570 88.980 64.580 89.150 ;
        RECT 64.750 88.980 64.940 89.150 ;
        RECT 65.110 88.980 65.130 89.150 ;
        RECT 64.570 87.650 65.130 88.980 ;
        RECT 66.490 89.200 67.940 89.230 ;
        RECT 66.490 89.030 66.740 89.200 ;
        RECT 66.910 89.030 67.100 89.200 ;
        RECT 67.270 89.030 67.540 89.200 ;
        RECT 67.710 89.030 67.940 89.200 ;
        RECT 62.400 86.320 63.700 86.720 ;
        RECT 62.090 85.840 63.700 86.320 ;
      LAYER li1 ;
        RECT 63.960 85.970 64.210 87.650 ;
      LAYER li1 ;
        RECT 64.520 86.760 64.850 87.220 ;
      LAYER li1 ;
        RECT 65.310 86.940 65.640 88.730 ;
      LAYER li1 ;
        RECT 65.820 86.760 66.070 88.480 ;
        RECT 66.490 88.160 67.940 89.030 ;
        RECT 68.730 89.150 69.320 89.230 ;
        RECT 68.730 88.980 68.760 89.150 ;
        RECT 68.930 88.980 69.120 89.150 ;
        RECT 69.290 88.980 69.320 89.150 ;
        RECT 64.520 86.590 66.070 86.760 ;
        RECT 64.390 85.840 65.640 86.410 ;
        RECT 65.820 85.970 66.070 86.590 ;
        RECT 66.720 86.720 67.050 87.500 ;
        RECT 67.260 87.170 67.590 88.160 ;
        RECT 68.730 87.650 69.320 88.980 ;
      LAYER li1 ;
        RECT 69.600 87.650 69.990 89.230 ;
      LAYER li1 ;
        RECT 70.330 89.200 71.780 89.230 ;
        RECT 70.330 89.030 70.580 89.200 ;
        RECT 70.750 89.030 70.940 89.200 ;
        RECT 71.110 89.030 71.380 89.200 ;
        RECT 71.550 89.030 71.780 89.200 ;
        RECT 70.330 88.160 71.780 89.030 ;
        RECT 72.090 89.150 73.020 89.230 ;
        RECT 72.090 88.980 72.110 89.150 ;
        RECT 72.280 88.980 72.470 89.150 ;
        RECT 72.640 88.980 72.830 89.150 ;
        RECT 73.000 88.980 73.020 89.150 ;
      LAYER li1 ;
        RECT 68.770 87.020 69.480 87.410 ;
      LAYER li1 ;
        RECT 66.720 86.320 68.020 86.720 ;
        RECT 66.410 85.840 68.020 86.320 ;
        RECT 68.730 85.840 69.320 86.800 ;
      LAYER li1 ;
        RECT 69.660 85.970 69.990 87.650 ;
      LAYER li1 ;
        RECT 70.560 86.720 70.890 87.500 ;
        RECT 71.100 87.170 71.430 88.160 ;
        RECT 72.090 87.650 73.020 88.980 ;
      LAYER li1 ;
        RECT 73.200 87.550 73.370 89.230 ;
      LAYER li1 ;
        RECT 73.550 89.150 74.800 89.230 ;
        RECT 73.720 88.980 73.910 89.150 ;
        RECT 74.080 88.980 74.270 89.150 ;
        RECT 74.440 88.980 74.630 89.150 ;
        RECT 73.550 87.730 74.800 88.980 ;
      LAYER li1 ;
        RECT 74.980 87.550 75.240 89.230 ;
      LAYER li1 ;
        RECT 75.610 89.200 77.060 89.230 ;
        RECT 75.610 89.030 75.860 89.200 ;
        RECT 76.030 89.030 76.220 89.200 ;
        RECT 76.390 89.030 76.660 89.200 ;
        RECT 76.830 89.030 77.060 89.200 ;
        RECT 75.610 88.160 77.060 89.030 ;
        RECT 77.370 89.150 78.320 89.230 ;
        RECT 77.370 88.980 77.400 89.150 ;
        RECT 77.570 88.980 77.760 89.150 ;
        RECT 77.930 88.980 78.120 89.150 ;
        RECT 78.290 88.980 78.320 89.150 ;
      LAYER li1 ;
        RECT 73.200 87.380 75.240 87.550 ;
        RECT 72.130 86.980 73.000 87.310 ;
      LAYER li1 ;
        RECT 70.560 86.320 71.860 86.720 ;
        RECT 70.250 85.840 71.860 86.320 ;
        RECT 72.090 85.840 73.710 86.800 ;
      LAYER li1 ;
        RECT 73.890 86.280 74.280 87.200 ;
        RECT 74.460 86.280 74.730 87.200 ;
        RECT 74.980 86.800 75.240 87.380 ;
        RECT 74.910 85.970 75.240 86.800 ;
      LAYER li1 ;
        RECT 75.840 86.720 76.170 87.500 ;
        RECT 76.380 87.170 76.710 88.160 ;
        RECT 77.370 87.650 78.320 88.980 ;
      LAYER li1 ;
        RECT 78.500 87.550 78.750 89.230 ;
      LAYER li1 ;
        RECT 78.930 89.150 79.880 89.230 ;
        RECT 78.930 88.980 78.960 89.150 ;
        RECT 79.130 88.980 79.320 89.150 ;
        RECT 79.490 88.980 79.680 89.150 ;
        RECT 79.850 88.980 79.880 89.150 ;
        RECT 78.930 87.730 79.880 88.980 ;
      LAYER li1 ;
        RECT 80.060 87.550 80.390 89.230 ;
      LAYER li1 ;
        RECT 80.570 89.150 81.520 89.230 ;
        RECT 80.570 88.980 80.600 89.150 ;
        RECT 80.770 88.980 80.960 89.150 ;
        RECT 81.130 88.980 81.320 89.150 ;
        RECT 81.490 88.980 81.520 89.150 ;
        RECT 80.570 87.770 81.520 88.980 ;
      LAYER li1 ;
        RECT 78.500 87.380 80.390 87.550 ;
        RECT 78.500 87.250 78.670 87.380 ;
        RECT 81.170 87.250 81.500 87.590 ;
        RECT 77.410 87.020 78.670 87.250 ;
      LAYER li1 ;
        RECT 78.850 87.070 80.880 87.200 ;
        RECT 81.700 87.070 81.950 89.230 ;
        RECT 82.330 89.200 83.780 89.230 ;
        RECT 82.330 89.030 82.580 89.200 ;
        RECT 82.750 89.030 82.940 89.200 ;
        RECT 83.110 89.030 83.380 89.200 ;
        RECT 83.550 89.030 83.780 89.200 ;
        RECT 82.330 88.160 83.780 89.030 ;
        RECT 84.090 89.150 85.040 89.230 ;
        RECT 84.090 88.980 84.120 89.150 ;
        RECT 84.290 88.980 84.480 89.150 ;
        RECT 84.650 88.980 84.840 89.150 ;
        RECT 85.010 88.980 85.040 89.150 ;
        RECT 78.850 87.030 81.950 87.070 ;
      LAYER li1 ;
        RECT 78.500 86.850 78.670 87.020 ;
      LAYER li1 ;
        RECT 80.710 86.900 81.950 87.030 ;
        RECT 75.840 86.320 77.140 86.720 ;
        RECT 75.530 85.840 77.140 86.320 ;
        RECT 77.370 85.840 78.320 86.800 ;
      LAYER li1 ;
        RECT 78.500 86.680 80.310 86.850 ;
        RECT 78.500 85.970 78.750 86.680 ;
      LAYER li1 ;
        RECT 78.930 85.840 79.880 86.500 ;
      LAYER li1 ;
        RECT 80.060 85.970 80.310 86.680 ;
      LAYER li1 ;
        RECT 80.490 85.840 81.440 86.720 ;
        RECT 81.620 85.970 81.950 86.900 ;
        RECT 82.560 86.720 82.890 87.500 ;
        RECT 83.100 87.170 83.430 88.160 ;
        RECT 84.090 87.650 85.040 88.980 ;
      LAYER li1 ;
        RECT 85.220 87.550 85.470 89.230 ;
      LAYER li1 ;
        RECT 85.650 89.150 86.600 89.230 ;
        RECT 85.650 88.980 85.680 89.150 ;
        RECT 85.850 88.980 86.040 89.150 ;
        RECT 86.210 88.980 86.400 89.150 ;
        RECT 86.570 88.980 86.600 89.150 ;
        RECT 85.650 87.730 86.600 88.980 ;
      LAYER li1 ;
        RECT 86.780 87.550 87.110 89.230 ;
      LAYER li1 ;
        RECT 87.290 89.150 88.240 89.230 ;
        RECT 87.290 88.980 87.320 89.150 ;
        RECT 87.490 88.980 87.680 89.150 ;
        RECT 87.850 88.980 88.040 89.150 ;
        RECT 88.210 88.980 88.240 89.150 ;
        RECT 87.290 87.770 88.240 88.980 ;
      LAYER li1 ;
        RECT 85.220 87.380 87.110 87.550 ;
        RECT 85.220 87.250 85.390 87.380 ;
        RECT 87.890 87.250 88.220 87.590 ;
        RECT 84.130 87.020 85.390 87.250 ;
      LAYER li1 ;
        RECT 85.570 87.070 87.600 87.200 ;
        RECT 88.420 87.070 88.670 89.230 ;
        RECT 89.300 89.200 92.040 89.220 ;
        RECT 89.300 89.030 89.510 89.200 ;
        RECT 89.680 89.030 89.950 89.200 ;
        RECT 90.120 89.030 90.360 89.200 ;
        RECT 90.530 89.030 90.790 89.200 ;
        RECT 90.960 89.030 91.230 89.200 ;
        RECT 91.400 89.030 91.640 89.200 ;
        RECT 91.810 89.030 92.040 89.200 ;
        RECT 89.300 88.150 92.040 89.030 ;
        RECT 93.690 89.150 94.640 89.230 ;
        RECT 93.690 88.980 93.720 89.150 ;
        RECT 93.890 88.980 94.080 89.150 ;
        RECT 94.250 88.980 94.440 89.150 ;
        RECT 94.610 88.980 94.640 89.150 ;
        RECT 85.570 87.030 88.670 87.070 ;
      LAYER li1 ;
        RECT 85.220 86.850 85.390 87.020 ;
      LAYER li1 ;
        RECT 87.430 86.900 88.670 87.030 ;
        RECT 82.560 86.320 83.860 86.720 ;
        RECT 82.250 85.840 83.860 86.320 ;
        RECT 84.090 85.840 85.040 86.800 ;
      LAYER li1 ;
        RECT 85.220 86.680 87.030 86.850 ;
        RECT 85.220 85.970 85.470 86.680 ;
      LAYER li1 ;
        RECT 85.650 85.840 86.600 86.500 ;
      LAYER li1 ;
        RECT 86.780 85.970 87.030 86.680 ;
      LAYER li1 ;
        RECT 87.210 85.840 88.160 86.720 ;
        RECT 88.340 85.970 88.670 86.900 ;
        RECT 89.540 86.830 89.870 87.500 ;
        RECT 90.270 87.170 90.600 88.150 ;
        RECT 90.820 86.830 91.150 87.500 ;
        RECT 91.550 87.170 91.880 88.150 ;
        RECT 93.690 87.650 94.640 88.980 ;
      LAYER li1 ;
        RECT 94.820 87.550 95.070 89.230 ;
      LAYER li1 ;
        RECT 95.250 89.150 96.200 89.230 ;
        RECT 95.250 88.980 95.280 89.150 ;
        RECT 95.450 88.980 95.640 89.150 ;
        RECT 95.810 88.980 96.000 89.150 ;
        RECT 96.170 88.980 96.200 89.150 ;
        RECT 95.250 87.730 96.200 88.980 ;
      LAYER li1 ;
        RECT 96.380 87.550 96.710 89.230 ;
      LAYER li1 ;
        RECT 96.890 89.150 97.840 89.230 ;
        RECT 96.890 88.980 96.920 89.150 ;
        RECT 97.090 88.980 97.280 89.150 ;
        RECT 97.450 88.980 97.640 89.150 ;
        RECT 97.810 88.980 97.840 89.150 ;
        RECT 96.890 87.770 97.840 88.980 ;
      LAYER li1 ;
        RECT 94.820 87.380 96.710 87.550 ;
        RECT 94.820 87.250 94.990 87.380 ;
        RECT 97.490 87.250 97.820 87.590 ;
        RECT 93.730 87.020 94.990 87.250 ;
      LAYER li1 ;
        RECT 95.170 87.070 97.200 87.200 ;
        RECT 98.020 87.070 98.270 89.230 ;
        RECT 98.650 89.200 100.100 89.230 ;
        RECT 98.650 89.030 98.900 89.200 ;
        RECT 99.070 89.030 99.260 89.200 ;
        RECT 99.430 89.030 99.700 89.200 ;
        RECT 99.870 89.030 100.100 89.200 ;
        RECT 98.650 88.160 100.100 89.030 ;
        RECT 95.170 87.030 98.270 87.070 ;
      LAYER li1 ;
        RECT 94.820 86.850 94.990 87.020 ;
      LAYER li1 ;
        RECT 97.030 86.900 98.270 87.030 ;
        RECT 89.380 85.830 92.110 86.830 ;
        RECT 93.690 85.840 94.640 86.800 ;
      LAYER li1 ;
        RECT 94.820 86.680 96.630 86.850 ;
        RECT 94.820 85.970 95.070 86.680 ;
      LAYER li1 ;
        RECT 95.250 85.840 96.200 86.500 ;
      LAYER li1 ;
        RECT 96.380 85.970 96.630 86.680 ;
      LAYER li1 ;
        RECT 96.810 85.840 97.760 86.720 ;
        RECT 97.940 85.970 98.270 86.900 ;
        RECT 98.880 86.720 99.210 87.500 ;
        RECT 99.420 87.170 99.750 88.160 ;
      LAYER li1 ;
        RECT 101.890 87.400 102.260 89.230 ;
      LAYER li1 ;
        RECT 102.440 89.150 103.020 89.230 ;
        RECT 107.290 89.200 108.740 89.230 ;
        RECT 102.440 88.980 102.460 89.150 ;
        RECT 102.630 88.980 102.820 89.150 ;
        RECT 102.990 88.980 103.020 89.150 ;
        RECT 102.440 87.650 103.020 88.980 ;
        RECT 105.170 89.150 106.480 89.180 ;
        RECT 105.170 88.980 105.200 89.150 ;
        RECT 105.370 88.980 105.560 89.150 ;
        RECT 105.730 88.980 105.920 89.150 ;
        RECT 106.090 88.980 106.280 89.150 ;
        RECT 106.450 88.980 106.480 89.150 ;
      LAYER li1 ;
        RECT 103.200 88.570 104.990 88.740 ;
      LAYER li1 ;
        RECT 98.880 86.320 100.180 86.720 ;
        RECT 98.570 85.840 100.180 86.320 ;
      LAYER li1 ;
        RECT 101.890 85.970 102.180 87.400 ;
      LAYER li1 ;
        RECT 102.380 87.000 102.710 87.220 ;
      LAYER li1 ;
        RECT 103.200 87.180 103.530 88.570 ;
      LAYER li1 ;
        RECT 104.310 88.060 104.640 88.390 ;
        RECT 103.710 87.890 104.640 88.060 ;
        RECT 103.710 87.000 103.880 87.890 ;
      LAYER li1 ;
        RECT 104.820 87.780 104.990 88.570 ;
      LAYER li1 ;
        RECT 105.170 87.970 106.480 88.980 ;
        RECT 107.290 89.030 107.540 89.200 ;
        RECT 107.710 89.030 107.900 89.200 ;
        RECT 108.070 89.030 108.340 89.200 ;
        RECT 108.510 89.030 108.740 89.200 ;
      LAYER li1 ;
        RECT 104.060 87.430 104.390 87.710 ;
        RECT 104.820 87.610 106.440 87.780 ;
        RECT 104.060 87.260 104.670 87.430 ;
      LAYER li1 ;
        RECT 102.380 86.830 104.320 87.000 ;
        RECT 102.360 85.840 103.970 86.650 ;
        RECT 104.150 86.390 104.320 86.830 ;
      LAYER li1 ;
        RECT 104.500 86.860 104.670 87.260 ;
        RECT 104.500 86.570 105.450 86.860 ;
      LAYER li1 ;
        RECT 105.630 86.750 105.880 87.250 ;
      LAYER li1 ;
        RECT 106.130 87.020 106.440 87.610 ;
      LAYER li1 ;
        RECT 106.660 86.750 106.910 88.390 ;
        RECT 107.290 88.160 108.740 89.030 ;
        RECT 109.050 89.150 110.720 89.230 ;
        RECT 109.050 88.980 109.080 89.150 ;
        RECT 109.250 88.980 109.440 89.150 ;
        RECT 109.610 88.980 109.800 89.150 ;
        RECT 109.970 88.980 110.160 89.150 ;
        RECT 110.330 88.980 110.520 89.150 ;
        RECT 110.690 88.980 110.720 89.150 ;
        RECT 105.630 86.580 106.910 86.750 ;
        RECT 104.150 85.970 104.640 86.390 ;
        RECT 104.820 85.840 106.480 86.390 ;
        RECT 106.660 85.970 106.910 86.580 ;
        RECT 107.520 86.720 107.850 87.500 ;
        RECT 108.060 87.170 108.390 88.160 ;
        RECT 109.050 87.770 110.720 88.980 ;
      LAYER li1 ;
        RECT 109.090 87.250 110.280 87.590 ;
        RECT 110.460 87.250 110.790 87.590 ;
        RECT 110.980 87.070 111.240 89.230 ;
      LAYER li1 ;
        RECT 111.610 89.200 113.060 89.230 ;
        RECT 111.610 89.030 111.860 89.200 ;
        RECT 112.030 89.030 112.220 89.200 ;
        RECT 112.390 89.030 112.660 89.200 ;
        RECT 112.830 89.030 113.060 89.200 ;
        RECT 111.610 88.160 113.060 89.030 ;
      LAYER li1 ;
        RECT 110.160 86.900 111.240 87.070 ;
      LAYER li1 ;
        RECT 107.520 86.320 108.820 86.720 ;
        RECT 107.210 85.840 108.820 86.320 ;
        RECT 109.050 85.840 109.980 86.800 ;
      LAYER li1 ;
        RECT 110.160 85.970 110.490 86.900 ;
      LAYER li1 ;
        RECT 111.840 86.720 112.170 87.500 ;
        RECT 112.380 87.170 112.710 88.160 ;
      LAYER li1 ;
        RECT 113.400 87.650 113.830 89.230 ;
      LAYER li1 ;
        RECT 114.010 89.150 114.570 89.230 ;
        RECT 114.010 88.980 114.020 89.150 ;
        RECT 114.190 88.980 114.380 89.150 ;
        RECT 114.550 88.980 114.570 89.150 ;
        RECT 114.010 87.650 114.570 88.980 ;
        RECT 115.930 89.200 117.380 89.230 ;
        RECT 115.930 89.030 116.180 89.200 ;
        RECT 116.350 89.030 116.540 89.200 ;
        RECT 116.710 89.030 116.980 89.200 ;
        RECT 117.150 89.030 117.380 89.200 ;
        RECT 110.680 85.840 111.270 86.720 ;
        RECT 111.840 86.320 113.140 86.720 ;
        RECT 111.530 85.840 113.140 86.320 ;
      LAYER li1 ;
        RECT 113.400 85.970 113.650 87.650 ;
      LAYER li1 ;
        RECT 113.960 86.760 114.290 87.220 ;
      LAYER li1 ;
        RECT 114.750 86.940 115.080 88.730 ;
      LAYER li1 ;
        RECT 115.260 86.760 115.510 88.480 ;
        RECT 115.930 88.160 117.380 89.030 ;
        RECT 113.960 86.590 115.510 86.760 ;
        RECT 113.830 85.840 115.080 86.410 ;
        RECT 115.260 85.970 115.510 86.590 ;
        RECT 116.160 86.720 116.490 87.500 ;
        RECT 116.700 87.170 117.030 88.160 ;
      LAYER li1 ;
        RECT 118.200 87.650 118.630 89.230 ;
      LAYER li1 ;
        RECT 118.810 89.150 119.370 89.230 ;
        RECT 118.810 88.980 118.820 89.150 ;
        RECT 118.990 88.980 119.180 89.150 ;
        RECT 119.350 88.980 119.370 89.150 ;
        RECT 118.810 87.650 119.370 88.980 ;
        RECT 120.980 89.200 123.720 89.220 ;
        RECT 120.980 89.030 121.190 89.200 ;
        RECT 121.360 89.030 121.630 89.200 ;
        RECT 121.800 89.030 122.040 89.200 ;
        RECT 122.210 89.030 122.470 89.200 ;
        RECT 122.640 89.030 122.910 89.200 ;
        RECT 123.080 89.030 123.320 89.200 ;
        RECT 123.490 89.030 123.720 89.200 ;
        RECT 116.160 86.320 117.460 86.720 ;
        RECT 115.850 85.840 117.460 86.320 ;
      LAYER li1 ;
        RECT 118.200 85.970 118.450 87.650 ;
      LAYER li1 ;
        RECT 118.760 86.760 119.090 87.220 ;
      LAYER li1 ;
        RECT 119.550 86.940 119.880 88.730 ;
      LAYER li1 ;
        RECT 120.060 86.760 120.310 88.480 ;
        RECT 120.980 88.150 123.720 89.030 ;
        RECT 124.820 89.200 127.560 89.220 ;
        RECT 124.820 89.030 125.030 89.200 ;
        RECT 125.200 89.030 125.470 89.200 ;
        RECT 125.640 89.030 125.880 89.200 ;
        RECT 126.050 89.030 126.310 89.200 ;
        RECT 126.480 89.030 126.750 89.200 ;
        RECT 126.920 89.030 127.160 89.200 ;
        RECT 127.330 89.030 127.560 89.200 ;
        RECT 124.820 88.150 127.560 89.030 ;
        RECT 128.660 89.200 131.400 89.220 ;
        RECT 128.660 89.030 128.870 89.200 ;
        RECT 129.040 89.030 129.310 89.200 ;
        RECT 129.480 89.030 129.720 89.200 ;
        RECT 129.890 89.030 130.150 89.200 ;
        RECT 130.320 89.030 130.590 89.200 ;
        RECT 130.760 89.030 131.000 89.200 ;
        RECT 131.170 89.030 131.400 89.200 ;
        RECT 128.660 88.150 131.400 89.030 ;
        RECT 132.250 89.200 133.700 89.230 ;
        RECT 132.250 89.030 132.500 89.200 ;
        RECT 132.670 89.030 132.860 89.200 ;
        RECT 133.030 89.030 133.300 89.200 ;
        RECT 133.470 89.030 133.700 89.200 ;
        RECT 132.250 88.160 133.700 89.030 ;
        RECT 134.620 89.150 135.270 89.260 ;
        RECT 134.620 88.980 134.680 89.150 ;
        RECT 134.850 88.980 135.040 89.150 ;
        RECT 135.210 88.980 135.270 89.150 ;
        RECT 134.620 88.920 135.270 88.980 ;
        RECT 134.620 88.650 135.020 88.920 ;
      LAYER li1 ;
        RECT 135.930 88.650 136.510 89.290 ;
      LAYER li1 ;
        RECT 137.300 89.200 140.040 89.220 ;
        RECT 137.300 89.030 137.510 89.200 ;
        RECT 137.680 89.030 137.950 89.200 ;
        RECT 138.120 89.030 138.360 89.200 ;
        RECT 138.530 89.030 138.790 89.200 ;
        RECT 138.960 89.030 139.230 89.200 ;
        RECT 139.400 89.030 139.640 89.200 ;
        RECT 139.810 89.030 140.040 89.200 ;
        RECT 121.220 86.830 121.550 87.500 ;
        RECT 121.950 87.170 122.280 88.150 ;
        RECT 122.500 86.830 122.830 87.500 ;
        RECT 123.230 87.170 123.560 88.150 ;
        RECT 125.060 86.830 125.390 87.500 ;
        RECT 125.790 87.170 126.120 88.150 ;
        RECT 126.340 86.830 126.670 87.500 ;
        RECT 127.070 87.170 127.400 88.150 ;
        RECT 128.900 86.830 129.230 87.500 ;
        RECT 129.630 87.170 129.960 88.150 ;
        RECT 130.180 86.830 130.510 87.500 ;
        RECT 130.910 87.170 131.240 88.150 ;
        RECT 118.760 86.590 120.310 86.760 ;
        RECT 118.630 85.840 119.880 86.410 ;
        RECT 120.060 85.970 120.310 86.590 ;
        RECT 121.060 85.830 123.790 86.830 ;
        RECT 124.900 85.830 127.630 86.830 ;
        RECT 128.740 85.830 131.470 86.830 ;
        RECT 132.480 86.720 132.810 87.500 ;
        RECT 133.020 87.170 133.350 88.160 ;
      LAYER li1 ;
        RECT 135.930 87.240 136.200 88.650 ;
      LAYER li1 ;
        RECT 137.300 88.150 140.040 89.030 ;
      LAYER li1 ;
        RECT 135.440 86.970 136.200 87.240 ;
      LAYER li1 ;
        RECT 132.480 86.320 133.780 86.720 ;
        RECT 132.170 85.840 133.780 86.320 ;
      LAYER li1 ;
        RECT 135.440 85.970 135.770 86.970 ;
      LAYER li1 ;
        RECT 137.540 86.830 137.870 87.500 ;
        RECT 138.270 87.170 138.600 88.150 ;
        RECT 138.820 86.830 139.150 87.500 ;
        RECT 139.550 87.170 139.880 88.150 ;
        RECT 136.180 86.100 136.590 86.540 ;
        RECT 135.940 85.760 136.590 86.100 ;
        RECT 137.380 85.830 140.110 86.830 ;
        RECT 5.760 85.380 5.920 85.560 ;
        RECT 6.090 85.380 6.400 85.560 ;
        RECT 6.570 85.380 6.880 85.560 ;
        RECT 7.050 85.380 7.360 85.560 ;
        RECT 7.530 85.380 7.840 85.560 ;
        RECT 8.010 85.380 8.320 85.560 ;
        RECT 8.490 85.380 8.800 85.560 ;
        RECT 8.970 85.380 9.280 85.560 ;
        RECT 9.450 85.380 9.760 85.560 ;
        RECT 9.930 85.380 10.240 85.560 ;
        RECT 10.410 85.380 10.720 85.560 ;
        RECT 10.890 85.380 11.200 85.560 ;
        RECT 11.370 85.380 11.680 85.560 ;
        RECT 11.850 85.380 12.160 85.560 ;
        RECT 12.330 85.380 12.640 85.560 ;
        RECT 12.810 85.380 13.120 85.560 ;
        RECT 13.290 85.380 13.600 85.560 ;
        RECT 13.770 85.380 14.080 85.560 ;
        RECT 14.250 85.380 14.560 85.560 ;
        RECT 14.730 85.380 15.040 85.560 ;
        RECT 15.210 85.380 15.520 85.560 ;
        RECT 15.690 85.380 16.000 85.560 ;
        RECT 16.170 85.380 16.480 85.560 ;
        RECT 16.650 85.380 16.960 85.560 ;
        RECT 17.130 85.380 17.440 85.560 ;
        RECT 17.610 85.380 17.920 85.560 ;
        RECT 18.090 85.380 18.400 85.560 ;
        RECT 18.570 85.380 18.880 85.560 ;
        RECT 19.050 85.380 19.360 85.560 ;
        RECT 19.530 85.380 19.840 85.560 ;
        RECT 20.010 85.380 20.160 85.560 ;
        RECT 20.640 85.380 20.800 85.560 ;
        RECT 20.970 85.380 21.280 85.560 ;
        RECT 21.450 85.380 21.760 85.560 ;
        RECT 21.930 85.380 22.240 85.560 ;
        RECT 22.410 85.380 22.720 85.560 ;
        RECT 22.890 85.380 23.200 85.560 ;
        RECT 23.370 85.380 23.680 85.560 ;
        RECT 23.850 85.380 24.160 85.560 ;
        RECT 24.330 85.380 24.640 85.560 ;
        RECT 24.810 85.380 25.120 85.560 ;
        RECT 25.290 85.380 25.600 85.560 ;
        RECT 25.770 85.380 26.080 85.560 ;
        RECT 26.250 85.380 26.560 85.560 ;
        RECT 26.730 85.380 27.040 85.560 ;
        RECT 27.210 85.380 27.520 85.560 ;
        RECT 27.690 85.380 28.000 85.560 ;
        RECT 28.170 85.380 28.480 85.560 ;
        RECT 28.650 85.380 28.960 85.560 ;
        RECT 29.130 85.380 29.440 85.560 ;
        RECT 29.610 85.380 29.920 85.560 ;
        RECT 30.090 85.380 30.400 85.560 ;
        RECT 30.570 85.380 30.880 85.560 ;
        RECT 31.050 85.380 31.360 85.560 ;
        RECT 31.530 85.380 31.840 85.560 ;
        RECT 32.010 85.380 32.320 85.560 ;
        RECT 32.490 85.380 32.800 85.560 ;
        RECT 32.970 85.380 33.280 85.560 ;
        RECT 33.450 85.380 33.760 85.560 ;
        RECT 33.930 85.380 34.240 85.560 ;
        RECT 34.410 85.380 34.720 85.560 ;
        RECT 34.890 85.380 35.200 85.560 ;
        RECT 35.370 85.380 35.680 85.560 ;
        RECT 35.850 85.380 36.160 85.560 ;
        RECT 36.330 85.380 36.640 85.560 ;
        RECT 36.810 85.380 37.120 85.560 ;
        RECT 37.290 85.380 37.600 85.560 ;
        RECT 37.770 85.380 38.080 85.560 ;
        RECT 38.250 85.380 38.560 85.560 ;
        RECT 38.730 85.380 39.040 85.560 ;
        RECT 39.210 85.380 39.520 85.560 ;
        RECT 39.690 85.380 40.000 85.560 ;
        RECT 40.170 85.380 40.480 85.560 ;
        RECT 40.650 85.380 40.960 85.560 ;
        RECT 41.130 85.380 41.440 85.560 ;
        RECT 41.610 85.380 41.920 85.560 ;
        RECT 42.090 85.380 42.400 85.560 ;
        RECT 42.570 85.380 42.880 85.560 ;
        RECT 43.050 85.380 43.360 85.560 ;
        RECT 43.530 85.380 43.840 85.560 ;
        RECT 44.010 85.380 44.320 85.560 ;
        RECT 44.490 85.380 44.800 85.560 ;
        RECT 44.970 85.380 45.280 85.560 ;
        RECT 45.450 85.380 45.760 85.560 ;
        RECT 45.930 85.380 46.240 85.560 ;
        RECT 46.410 85.380 46.720 85.560 ;
        RECT 46.890 85.380 47.200 85.560 ;
        RECT 47.370 85.380 47.680 85.560 ;
        RECT 47.850 85.380 48.160 85.560 ;
        RECT 48.330 85.380 48.640 85.560 ;
        RECT 48.810 85.380 49.120 85.560 ;
        RECT 49.290 85.380 49.600 85.560 ;
        RECT 49.770 85.380 50.080 85.560 ;
        RECT 50.250 85.380 50.560 85.560 ;
        RECT 50.730 85.380 51.040 85.560 ;
        RECT 51.210 85.380 51.520 85.560 ;
        RECT 51.690 85.380 52.000 85.560 ;
        RECT 52.170 85.380 52.480 85.560 ;
        RECT 52.650 85.380 52.960 85.560 ;
        RECT 53.130 85.380 53.440 85.560 ;
        RECT 53.610 85.380 53.920 85.560 ;
        RECT 54.090 85.380 54.400 85.560 ;
        RECT 54.570 85.380 54.880 85.560 ;
        RECT 55.050 85.380 55.360 85.560 ;
        RECT 55.530 85.380 55.840 85.560 ;
        RECT 56.010 85.380 56.320 85.560 ;
        RECT 56.490 85.380 56.800 85.560 ;
        RECT 56.970 85.380 57.280 85.560 ;
        RECT 57.450 85.380 57.760 85.560 ;
        RECT 57.930 85.380 58.240 85.560 ;
        RECT 58.410 85.380 58.720 85.560 ;
        RECT 58.890 85.380 59.200 85.560 ;
        RECT 59.370 85.380 59.680 85.560 ;
        RECT 59.850 85.380 60.160 85.560 ;
        RECT 60.330 85.380 60.640 85.560 ;
        RECT 60.810 85.380 61.120 85.560 ;
        RECT 61.290 85.380 61.600 85.560 ;
        RECT 61.770 85.380 62.080 85.560 ;
        RECT 62.250 85.380 62.560 85.560 ;
        RECT 62.730 85.380 63.040 85.560 ;
        RECT 63.210 85.380 63.520 85.560 ;
        RECT 63.690 85.380 64.000 85.560 ;
        RECT 64.170 85.380 64.480 85.560 ;
        RECT 64.650 85.380 64.960 85.560 ;
        RECT 65.130 85.380 65.440 85.560 ;
        RECT 65.610 85.380 65.920 85.560 ;
        RECT 66.090 85.380 66.400 85.560 ;
        RECT 66.570 85.380 66.880 85.560 ;
        RECT 67.050 85.380 67.360 85.560 ;
        RECT 67.530 85.380 67.840 85.560 ;
        RECT 68.010 85.380 68.160 85.560 ;
        RECT 68.640 85.380 68.800 85.560 ;
        RECT 68.970 85.380 69.280 85.560 ;
        RECT 69.450 85.380 69.760 85.560 ;
        RECT 69.930 85.380 70.240 85.560 ;
        RECT 70.410 85.380 70.720 85.560 ;
        RECT 70.890 85.380 71.200 85.560 ;
        RECT 71.370 85.380 71.680 85.560 ;
        RECT 71.850 85.380 72.160 85.560 ;
        RECT 72.330 85.380 72.640 85.560 ;
        RECT 72.810 85.380 73.120 85.560 ;
        RECT 73.290 85.380 73.600 85.560 ;
        RECT 73.770 85.380 74.080 85.560 ;
        RECT 74.250 85.380 74.560 85.560 ;
        RECT 74.730 85.380 75.040 85.560 ;
        RECT 75.210 85.380 75.520 85.560 ;
        RECT 75.690 85.380 76.000 85.560 ;
        RECT 76.170 85.380 76.480 85.560 ;
        RECT 76.650 85.380 76.960 85.560 ;
        RECT 77.130 85.380 77.440 85.560 ;
        RECT 77.610 85.380 77.920 85.560 ;
        RECT 78.090 85.380 78.400 85.560 ;
        RECT 78.570 85.380 78.880 85.560 ;
        RECT 79.050 85.380 79.360 85.560 ;
        RECT 79.530 85.380 79.840 85.560 ;
        RECT 80.010 85.380 80.320 85.560 ;
        RECT 80.490 85.380 80.800 85.560 ;
        RECT 80.970 85.380 81.280 85.560 ;
        RECT 81.450 85.380 81.760 85.560 ;
        RECT 81.930 85.380 82.240 85.560 ;
        RECT 82.410 85.380 82.720 85.560 ;
        RECT 82.890 85.380 83.200 85.560 ;
        RECT 83.370 85.380 83.680 85.560 ;
        RECT 83.850 85.380 84.160 85.560 ;
        RECT 84.330 85.380 84.640 85.560 ;
        RECT 84.810 85.380 85.120 85.560 ;
        RECT 85.290 85.380 85.600 85.560 ;
        RECT 85.770 85.380 86.080 85.560 ;
        RECT 86.250 85.380 86.560 85.560 ;
        RECT 86.730 85.380 87.040 85.560 ;
        RECT 87.210 85.380 87.520 85.560 ;
        RECT 87.690 85.380 88.000 85.560 ;
        RECT 88.170 85.380 88.480 85.560 ;
        RECT 88.650 85.380 88.960 85.560 ;
        RECT 89.130 85.380 89.440 85.560 ;
        RECT 89.610 85.380 89.920 85.560 ;
        RECT 90.090 85.380 90.400 85.560 ;
        RECT 90.570 85.380 90.880 85.560 ;
        RECT 91.050 85.380 91.360 85.560 ;
        RECT 91.530 85.380 91.840 85.560 ;
        RECT 92.010 85.380 92.320 85.560 ;
        RECT 92.490 85.380 92.800 85.560 ;
        RECT 92.970 85.380 93.280 85.560 ;
        RECT 93.450 85.380 93.760 85.560 ;
        RECT 93.930 85.380 94.240 85.560 ;
        RECT 94.410 85.380 94.720 85.560 ;
        RECT 94.890 85.380 95.200 85.560 ;
        RECT 95.370 85.380 95.680 85.560 ;
        RECT 95.850 85.380 96.160 85.560 ;
        RECT 96.330 85.380 96.640 85.560 ;
        RECT 96.810 85.380 97.120 85.560 ;
        RECT 97.290 85.380 97.600 85.560 ;
        RECT 97.770 85.380 98.080 85.560 ;
        RECT 98.250 85.380 98.560 85.560 ;
        RECT 98.730 85.380 99.040 85.560 ;
        RECT 99.210 85.380 99.520 85.560 ;
        RECT 99.690 85.380 100.000 85.560 ;
        RECT 100.170 85.380 100.480 85.560 ;
        RECT 100.650 85.380 100.960 85.560 ;
        RECT 101.130 85.380 101.280 85.560 ;
        RECT 101.760 85.380 101.920 85.560 ;
        RECT 102.090 85.380 102.400 85.560 ;
        RECT 102.570 85.380 102.880 85.560 ;
        RECT 103.050 85.380 103.360 85.560 ;
        RECT 103.530 85.380 103.840 85.560 ;
        RECT 104.010 85.380 104.320 85.560 ;
        RECT 104.490 85.380 104.800 85.560 ;
        RECT 104.970 85.380 105.280 85.560 ;
        RECT 105.450 85.380 105.760 85.560 ;
        RECT 105.930 85.380 106.240 85.560 ;
        RECT 106.410 85.380 106.720 85.560 ;
        RECT 106.890 85.380 107.200 85.560 ;
        RECT 107.370 85.380 107.680 85.560 ;
        RECT 107.850 85.380 108.160 85.560 ;
        RECT 108.330 85.380 108.640 85.560 ;
        RECT 108.810 85.380 109.120 85.560 ;
        RECT 109.290 85.380 109.600 85.560 ;
        RECT 109.770 85.380 110.080 85.560 ;
        RECT 110.250 85.380 110.560 85.560 ;
        RECT 110.730 85.380 111.040 85.560 ;
        RECT 111.210 85.380 111.520 85.560 ;
        RECT 111.690 85.380 112.000 85.560 ;
        RECT 112.170 85.380 112.480 85.560 ;
        RECT 112.650 85.380 112.960 85.560 ;
        RECT 113.130 85.380 113.440 85.560 ;
        RECT 113.610 85.380 113.920 85.560 ;
        RECT 114.090 85.380 114.400 85.560 ;
        RECT 114.570 85.380 114.880 85.560 ;
        RECT 115.050 85.380 115.360 85.560 ;
        RECT 115.530 85.380 115.840 85.560 ;
        RECT 116.010 85.380 116.320 85.560 ;
        RECT 116.490 85.380 116.800 85.560 ;
        RECT 116.970 85.380 117.280 85.560 ;
        RECT 117.450 85.380 117.600 85.560 ;
        RECT 118.080 85.380 118.240 85.560 ;
        RECT 118.410 85.380 118.720 85.560 ;
        RECT 118.890 85.380 119.200 85.560 ;
        RECT 119.370 85.380 119.680 85.560 ;
        RECT 119.850 85.380 120.160 85.560 ;
        RECT 120.330 85.380 120.640 85.560 ;
        RECT 120.810 85.380 121.120 85.560 ;
        RECT 121.290 85.380 121.600 85.560 ;
        RECT 121.770 85.380 122.080 85.560 ;
        RECT 122.250 85.380 122.560 85.560 ;
        RECT 122.730 85.380 123.040 85.560 ;
        RECT 123.210 85.380 123.520 85.560 ;
        RECT 123.690 85.380 124.000 85.560 ;
        RECT 124.170 85.380 124.480 85.560 ;
        RECT 124.650 85.380 124.960 85.560 ;
        RECT 125.130 85.380 125.440 85.560 ;
        RECT 125.610 85.380 125.920 85.560 ;
        RECT 126.090 85.380 126.400 85.560 ;
        RECT 126.570 85.380 126.880 85.560 ;
        RECT 127.050 85.380 127.360 85.560 ;
        RECT 127.530 85.380 127.840 85.560 ;
        RECT 128.010 85.380 128.320 85.560 ;
        RECT 128.490 85.380 128.800 85.560 ;
        RECT 128.970 85.380 129.280 85.560 ;
        RECT 129.450 85.380 129.760 85.560 ;
        RECT 129.930 85.380 130.240 85.560 ;
        RECT 130.410 85.380 130.720 85.560 ;
        RECT 130.890 85.380 131.200 85.560 ;
        RECT 131.370 85.380 131.680 85.560 ;
        RECT 131.850 85.380 132.160 85.560 ;
        RECT 132.330 85.380 132.640 85.560 ;
        RECT 132.810 85.380 133.120 85.560 ;
        RECT 133.290 85.380 133.600 85.560 ;
        RECT 133.770 85.380 133.920 85.560 ;
        RECT 134.400 85.380 134.560 85.560 ;
        RECT 134.730 85.380 135.040 85.560 ;
        RECT 135.210 85.380 135.520 85.560 ;
        RECT 135.690 85.380 136.000 85.560 ;
        RECT 136.170 85.380 136.480 85.560 ;
        RECT 136.650 85.380 136.960 85.560 ;
        RECT 137.130 85.380 137.440 85.560 ;
        RECT 137.610 85.380 137.920 85.560 ;
        RECT 138.090 85.380 138.400 85.560 ;
        RECT 138.570 85.380 138.880 85.560 ;
        RECT 139.050 85.380 139.360 85.560 ;
        RECT 139.530 85.380 139.840 85.560 ;
        RECT 140.010 85.380 140.320 85.560 ;
        RECT 140.490 85.380 140.800 85.560 ;
        RECT 140.970 85.380 141.280 85.560 ;
        RECT 141.450 85.380 141.600 85.560 ;
        RECT 5.930 85.070 7.540 85.100 ;
        RECT 5.930 84.900 5.980 85.070 ;
        RECT 6.150 84.900 6.420 85.070 ;
        RECT 6.590 84.900 6.860 85.070 ;
        RECT 7.030 84.900 7.270 85.070 ;
        RECT 7.440 84.900 7.540 85.070 ;
        RECT 8.240 85.070 9.190 85.100 ;
        RECT 5.930 84.620 7.540 84.900 ;
        RECT 6.240 84.220 7.540 84.620 ;
        RECT 6.240 83.440 6.570 84.220 ;
        RECT 6.780 82.780 7.110 83.770 ;
        RECT 7.790 83.110 8.060 84.970 ;
        RECT 8.240 84.900 8.270 85.070 ;
        RECT 8.440 84.900 8.630 85.070 ;
        RECT 8.800 84.900 8.990 85.070 ;
        RECT 9.160 84.900 9.190 85.070 ;
        RECT 9.880 85.070 10.470 85.100 ;
        RECT 8.240 84.470 9.190 84.900 ;
        RECT 9.370 84.470 9.700 84.970 ;
        RECT 8.920 83.110 9.250 83.610 ;
        RECT 7.790 82.940 9.250 83.110 ;
        RECT 6.010 81.910 7.460 82.780 ;
        RECT 7.790 82.010 8.120 82.940 ;
        RECT 6.010 81.740 6.260 81.910 ;
        RECT 6.430 81.740 6.620 81.910 ;
        RECT 6.790 81.740 7.060 81.910 ;
        RECT 7.230 81.740 7.460 81.910 ;
        RECT 8.310 81.960 8.900 82.740 ;
        RECT 8.310 81.790 8.340 81.960 ;
        RECT 8.510 81.790 8.700 81.960 ;
        RECT 8.870 81.790 8.900 81.960 ;
        RECT 8.310 81.760 8.900 81.790 ;
        RECT 9.080 81.830 9.250 82.940 ;
        RECT 9.430 83.550 9.700 84.470 ;
        RECT 9.880 84.900 9.910 85.070 ;
        RECT 10.080 84.900 10.270 85.070 ;
        RECT 10.440 84.900 10.470 85.070 ;
        RECT 14.840 85.070 15.790 85.100 ;
        RECT 9.880 84.220 10.470 84.900 ;
      LAYER li1 ;
        RECT 10.750 84.840 13.690 85.010 ;
        RECT 10.750 83.850 10.920 84.840 ;
      LAYER li1 ;
        RECT 9.430 83.320 9.960 83.550 ;
        RECT 9.430 82.010 9.680 83.320 ;
      LAYER li1 ;
        RECT 10.380 82.980 10.920 83.850 ;
        RECT 11.100 83.360 11.430 84.660 ;
      LAYER li1 ;
        RECT 11.610 84.140 11.880 84.640 ;
        RECT 12.330 84.390 12.660 84.640 ;
        RECT 12.330 84.220 13.340 84.390 ;
        RECT 11.610 83.150 11.780 84.140 ;
        RECT 12.660 83.550 12.990 84.040 ;
        RECT 11.560 82.980 11.780 83.150 ;
        RECT 11.960 83.320 12.990 83.550 ;
        RECT 13.170 83.990 13.340 84.220 ;
      LAYER li1 ;
        RECT 13.520 84.340 13.690 84.840 ;
      LAYER li1 ;
        RECT 14.840 84.900 14.870 85.070 ;
        RECT 15.040 84.900 15.230 85.070 ;
        RECT 15.400 84.900 15.590 85.070 ;
        RECT 15.760 84.900 15.790 85.070 ;
        RECT 14.840 84.520 15.790 84.900 ;
      LAYER li1 ;
        RECT 15.970 85.030 18.630 85.200 ;
        RECT 15.970 84.340 16.140 85.030 ;
        RECT 13.520 84.170 16.140 84.340 ;
      LAYER li1 ;
        RECT 13.170 83.820 15.790 83.990 ;
        RECT 11.560 82.800 11.730 82.980 ;
        RECT 11.960 82.800 12.130 83.320 ;
        RECT 13.170 83.140 13.340 83.820 ;
      LAYER li1 ;
        RECT 15.970 83.640 16.140 84.170 ;
      LAYER li1 ;
        RECT 9.920 82.630 11.730 82.800 ;
        RECT 9.920 82.010 10.170 82.630 ;
        RECT 10.350 82.280 11.380 82.450 ;
        RECT 10.350 81.830 10.520 82.280 ;
        RECT 6.010 81.710 7.460 81.740 ;
        RECT 9.080 81.660 10.520 81.830 ;
        RECT 10.700 81.960 11.030 82.100 ;
        RECT 10.700 81.790 10.730 81.960 ;
        RECT 10.900 81.790 11.030 81.960 ;
        RECT 10.700 81.760 11.030 81.790 ;
        RECT 11.210 81.830 11.380 82.280 ;
        RECT 11.560 82.010 11.730 82.630 ;
        RECT 11.910 82.470 12.130 82.800 ;
        RECT 12.310 82.970 13.340 83.140 ;
        RECT 13.520 83.290 13.850 83.640 ;
      LAYER li1 ;
        RECT 14.290 83.470 16.140 83.640 ;
      LAYER li1 ;
        RECT 16.320 84.140 16.650 84.850 ;
        RECT 17.110 84.680 18.280 84.850 ;
        RECT 17.110 84.140 17.440 84.680 ;
        RECT 16.320 83.290 16.580 84.140 ;
        RECT 17.650 83.880 17.930 84.380 ;
        RECT 13.520 83.120 16.580 83.290 ;
        RECT 12.310 82.270 12.480 82.970 ;
        RECT 13.170 82.940 13.340 82.970 ;
        RECT 12.660 82.590 12.990 82.790 ;
        RECT 13.170 82.770 14.940 82.940 ;
        RECT 12.660 82.470 14.430 82.590 ;
        RECT 12.780 82.420 14.430 82.470 ;
        RECT 12.260 82.010 12.590 82.270 ;
        RECT 12.780 81.830 12.950 82.420 ;
        RECT 11.210 81.660 12.950 81.830 ;
        RECT 13.130 81.960 14.080 82.240 ;
        RECT 13.130 81.790 13.160 81.960 ;
        RECT 13.330 81.790 13.520 81.960 ;
        RECT 13.690 81.790 13.880 81.960 ;
        RECT 14.050 81.790 14.080 81.960 ;
        RECT 13.130 81.760 14.080 81.790 ;
        RECT 14.260 81.830 14.430 82.420 ;
        RECT 14.610 82.010 14.940 82.770 ;
        RECT 16.250 82.540 16.580 83.120 ;
        RECT 16.760 83.710 17.930 83.880 ;
        RECT 16.760 82.360 16.930 83.710 ;
        RECT 17.310 83.030 17.640 83.530 ;
        RECT 18.110 83.280 18.280 84.680 ;
      LAYER li1 ;
        RECT 18.460 84.370 18.630 85.030 ;
      LAYER li1 ;
        RECT 18.810 85.070 19.760 85.100 ;
        RECT 18.810 84.900 18.840 85.070 ;
        RECT 19.010 84.900 19.200 85.070 ;
        RECT 19.370 84.900 19.560 85.070 ;
        RECT 19.730 84.900 19.760 85.070 ;
        RECT 21.420 85.070 22.370 85.100 ;
        RECT 18.810 84.550 19.760 84.900 ;
        RECT 20.300 84.470 20.630 84.970 ;
        RECT 21.420 84.900 21.450 85.070 ;
        RECT 21.620 84.900 21.810 85.070 ;
        RECT 21.980 84.900 22.170 85.070 ;
        RECT 22.340 84.900 22.370 85.070 ;
      LAYER li1 ;
        RECT 18.460 84.260 19.470 84.370 ;
        RECT 18.460 84.200 19.520 84.260 ;
        RECT 19.140 84.090 19.520 84.200 ;
      LAYER li1 ;
        RECT 18.490 83.630 18.820 84.020 ;
      LAYER li1 ;
        RECT 19.140 83.810 19.470 84.090 ;
      LAYER li1 ;
        RECT 20.300 83.630 20.530 84.470 ;
        RECT 20.910 83.970 21.240 84.470 ;
        RECT 21.420 83.970 22.370 84.900 ;
        RECT 23.210 85.070 24.820 85.100 ;
        RECT 25.510 85.070 26.760 85.100 ;
        RECT 27.530 85.070 29.140 85.100 ;
        RECT 23.210 84.900 23.260 85.070 ;
        RECT 23.430 84.900 23.700 85.070 ;
        RECT 23.870 84.900 24.140 85.070 ;
        RECT 24.310 84.900 24.550 85.070 ;
        RECT 24.720 84.900 24.820 85.070 ;
        RECT 18.490 83.460 20.530 83.630 ;
        RECT 17.820 83.110 20.180 83.280 ;
        RECT 17.820 82.790 17.990 83.110 ;
        RECT 20.360 82.930 20.530 83.460 ;
        RECT 15.120 82.190 16.930 82.360 ;
        RECT 17.110 82.620 17.990 82.790 ;
        RECT 15.120 81.830 15.290 82.190 ;
        RECT 14.260 81.660 15.290 81.830 ;
        RECT 15.470 81.960 16.420 82.010 ;
        RECT 15.470 81.790 15.500 81.960 ;
        RECT 15.670 81.790 15.860 81.960 ;
        RECT 16.030 81.790 16.220 81.960 ;
        RECT 16.390 81.790 16.420 81.960 ;
        RECT 15.470 81.710 16.420 81.790 ;
        RECT 17.110 81.710 17.360 82.620 ;
        RECT 18.170 81.960 19.120 82.790 ;
        RECT 19.520 82.760 20.530 82.930 ;
        RECT 21.030 83.790 21.240 83.970 ;
        RECT 21.030 83.460 22.400 83.790 ;
        RECT 19.520 82.290 19.770 82.760 ;
        RECT 19.950 81.960 20.850 82.580 ;
        RECT 21.030 82.460 21.280 83.460 ;
        RECT 18.170 81.790 18.200 81.960 ;
        RECT 18.370 81.790 18.560 81.960 ;
        RECT 18.730 81.790 18.920 81.960 ;
        RECT 19.090 81.790 19.120 81.960 ;
        RECT 20.120 81.790 20.310 81.960 ;
        RECT 20.480 81.790 20.670 81.960 ;
        RECT 20.840 81.790 20.850 81.960 ;
        RECT 18.170 81.760 19.120 81.790 ;
        RECT 19.950 81.760 20.850 81.790 ;
        RECT 21.460 81.960 22.400 83.270 ;
        RECT 21.460 81.790 21.480 81.960 ;
        RECT 21.650 81.790 21.840 81.960 ;
        RECT 22.010 81.790 22.200 81.960 ;
        RECT 22.370 81.790 22.400 81.960 ;
        RECT 21.460 81.730 22.400 81.790 ;
      LAYER li1 ;
        RECT 22.580 81.730 22.920 84.800 ;
      LAYER li1 ;
        RECT 23.210 84.620 24.820 84.900 ;
        RECT 23.520 84.220 24.820 84.620 ;
        RECT 23.520 83.440 23.850 84.220 ;
        RECT 24.060 82.780 24.390 83.770 ;
      LAYER li1 ;
        RECT 25.080 83.290 25.330 84.970 ;
      LAYER li1 ;
        RECT 25.680 84.900 25.870 85.070 ;
        RECT 26.040 84.900 26.230 85.070 ;
        RECT 26.400 84.900 26.590 85.070 ;
        RECT 25.510 84.530 26.760 84.900 ;
        RECT 26.940 84.350 27.190 84.970 ;
        RECT 27.530 84.900 27.580 85.070 ;
        RECT 27.750 84.900 28.020 85.070 ;
        RECT 28.190 84.900 28.460 85.070 ;
        RECT 28.630 84.900 28.870 85.070 ;
        RECT 29.040 84.900 29.140 85.070 ;
        RECT 27.530 84.620 29.140 84.900 ;
        RECT 25.640 84.180 27.190 84.350 ;
        RECT 25.640 83.720 25.970 84.180 ;
        RECT 23.290 81.910 24.740 82.780 ;
        RECT 23.290 81.740 23.540 81.910 ;
        RECT 23.710 81.740 23.900 81.910 ;
        RECT 24.070 81.740 24.340 81.910 ;
        RECT 24.510 81.740 24.740 81.910 ;
        RECT 23.290 81.710 24.740 81.740 ;
      LAYER li1 ;
        RECT 25.080 81.710 25.510 83.290 ;
      LAYER li1 ;
        RECT 25.690 81.960 26.250 83.290 ;
      LAYER li1 ;
        RECT 26.430 82.210 26.760 84.000 ;
      LAYER li1 ;
        RECT 26.940 82.460 27.190 84.180 ;
        RECT 27.840 84.220 29.140 84.620 ;
        RECT 29.440 85.030 31.250 85.200 ;
        RECT 27.840 83.440 28.170 84.220 ;
        RECT 29.440 84.110 29.770 85.030 ;
      LAYER li1 ;
        RECT 30.020 84.110 30.550 84.850 ;
      LAYER li1 ;
        RECT 28.380 82.780 28.710 83.770 ;
      LAYER li1 ;
        RECT 29.410 83.600 29.830 83.930 ;
        RECT 30.020 83.540 30.190 84.110 ;
      LAYER li1 ;
        RECT 31.080 84.010 31.250 85.030 ;
        RECT 31.430 85.070 32.530 85.100 ;
        RECT 31.430 84.900 31.480 85.070 ;
        RECT 31.650 84.900 31.840 85.070 ;
        RECT 32.010 84.900 32.200 85.070 ;
        RECT 32.370 84.900 32.530 85.070 ;
        RECT 33.290 85.070 34.900 85.100 ;
        RECT 35.590 85.070 36.840 85.100 ;
        RECT 37.610 85.070 39.220 85.100 ;
        RECT 31.430 84.190 32.530 84.900 ;
        RECT 32.700 84.010 32.950 84.940 ;
        RECT 33.290 84.900 33.340 85.070 ;
        RECT 33.510 84.900 33.780 85.070 ;
        RECT 33.950 84.900 34.220 85.070 ;
        RECT 34.390 84.900 34.630 85.070 ;
        RECT 34.800 84.900 34.900 85.070 ;
        RECT 33.290 84.620 34.900 84.900 ;
      LAYER li1 ;
        RECT 30.370 83.720 30.880 83.930 ;
      LAYER li1 ;
        RECT 31.080 83.840 32.950 84.010 ;
        RECT 33.600 84.220 34.900 84.620 ;
      LAYER li1 ;
        RECT 30.020 83.370 31.080 83.540 ;
        RECT 30.810 83.290 31.080 83.370 ;
        RECT 31.530 83.350 32.040 83.660 ;
        RECT 32.290 83.350 33.000 83.660 ;
      LAYER li1 ;
        RECT 33.600 83.440 33.930 84.220 ;
        RECT 25.690 81.790 25.700 81.960 ;
        RECT 25.870 81.790 26.060 81.960 ;
        RECT 26.230 81.790 26.250 81.960 ;
        RECT 25.690 81.710 26.250 81.790 ;
        RECT 27.610 81.910 29.060 82.780 ;
        RECT 27.610 81.740 27.860 81.910 ;
        RECT 28.030 81.740 28.220 81.910 ;
        RECT 28.390 81.740 28.660 81.910 ;
        RECT 28.830 81.740 29.060 81.910 ;
        RECT 27.610 81.710 29.060 81.740 ;
        RECT 29.370 81.960 30.630 83.190 ;
      LAYER li1 ;
        RECT 30.810 82.210 31.330 83.290 ;
      LAYER li1 ;
        RECT 29.370 81.790 29.380 81.960 ;
        RECT 29.550 81.790 29.740 81.960 ;
        RECT 29.910 81.790 30.100 81.960 ;
        RECT 30.270 81.790 30.460 81.960 ;
        RECT 29.370 81.710 30.630 81.790 ;
      LAYER li1 ;
        RECT 31.160 81.710 31.330 82.210 ;
      LAYER li1 ;
        RECT 31.590 81.960 32.900 83.170 ;
        RECT 34.140 82.780 34.470 83.770 ;
      LAYER li1 ;
        RECT 35.160 83.290 35.410 84.970 ;
      LAYER li1 ;
        RECT 35.760 84.900 35.950 85.070 ;
        RECT 36.120 84.900 36.310 85.070 ;
        RECT 36.480 84.900 36.670 85.070 ;
        RECT 35.590 84.530 36.840 84.900 ;
        RECT 37.020 84.350 37.270 84.970 ;
        RECT 37.610 84.900 37.660 85.070 ;
        RECT 37.830 84.900 38.100 85.070 ;
        RECT 38.270 84.900 38.540 85.070 ;
        RECT 38.710 84.900 38.950 85.070 ;
        RECT 39.120 84.900 39.220 85.070 ;
        RECT 37.610 84.620 39.220 84.900 ;
        RECT 35.720 84.180 37.270 84.350 ;
        RECT 35.720 83.720 36.050 84.180 ;
        RECT 31.590 81.790 31.620 81.960 ;
        RECT 31.790 81.790 31.980 81.960 ;
        RECT 32.150 81.790 32.340 81.960 ;
        RECT 32.510 81.790 32.700 81.960 ;
        RECT 32.870 81.790 32.900 81.960 ;
        RECT 31.590 81.710 32.900 81.790 ;
        RECT 33.370 81.910 34.820 82.780 ;
        RECT 33.370 81.740 33.620 81.910 ;
        RECT 33.790 81.740 33.980 81.910 ;
        RECT 34.150 81.740 34.420 81.910 ;
        RECT 34.590 81.740 34.820 81.910 ;
        RECT 33.370 81.710 34.820 81.740 ;
      LAYER li1 ;
        RECT 35.160 81.710 35.590 83.290 ;
      LAYER li1 ;
        RECT 35.770 81.960 36.330 83.290 ;
      LAYER li1 ;
        RECT 36.510 82.210 36.840 84.000 ;
      LAYER li1 ;
        RECT 37.020 82.460 37.270 84.180 ;
        RECT 37.920 84.220 39.220 84.620 ;
        RECT 39.450 85.070 40.400 85.100 ;
        RECT 39.450 84.900 39.480 85.070 ;
        RECT 39.650 84.900 39.840 85.070 ;
        RECT 40.010 84.900 40.200 85.070 ;
        RECT 40.370 84.900 40.400 85.070 ;
        RECT 41.010 85.070 41.960 85.100 ;
        RECT 37.920 83.440 38.250 84.220 ;
        RECT 39.450 84.140 40.400 84.900 ;
      LAYER li1 ;
        RECT 40.580 84.260 40.830 84.970 ;
      LAYER li1 ;
        RECT 41.010 84.900 41.040 85.070 ;
        RECT 41.210 84.900 41.400 85.070 ;
        RECT 41.570 84.900 41.760 85.070 ;
        RECT 41.930 84.900 41.960 85.070 ;
        RECT 42.570 85.070 43.520 85.100 ;
        RECT 41.010 84.440 41.960 84.900 ;
      LAYER li1 ;
        RECT 42.140 84.260 42.390 84.970 ;
        RECT 40.580 84.090 42.390 84.260 ;
      LAYER li1 ;
        RECT 42.570 84.900 42.600 85.070 ;
        RECT 42.770 84.900 42.960 85.070 ;
        RECT 43.130 84.900 43.320 85.070 ;
        RECT 43.490 84.900 43.520 85.070 ;
        RECT 44.740 85.080 47.470 85.110 ;
        RECT 42.570 84.220 43.520 84.900 ;
      LAYER li1 ;
        RECT 40.580 83.920 40.750 84.090 ;
      LAYER li1 ;
        RECT 43.700 84.040 44.030 84.970 ;
        RECT 44.740 84.910 44.910 85.080 ;
        RECT 45.080 84.910 45.350 85.080 ;
        RECT 45.520 84.910 45.760 85.080 ;
        RECT 45.930 84.910 46.190 85.080 ;
        RECT 46.360 84.910 46.630 85.080 ;
        RECT 46.800 84.910 47.040 85.080 ;
        RECT 47.210 84.910 47.470 85.080 ;
        RECT 44.740 84.110 47.470 84.910 ;
        RECT 49.050 85.070 50.000 85.100 ;
        RECT 49.050 84.900 49.080 85.070 ;
        RECT 49.250 84.900 49.440 85.070 ;
        RECT 49.610 84.900 49.800 85.070 ;
        RECT 49.970 84.900 50.000 85.070 ;
        RECT 50.610 85.070 51.560 85.100 ;
        RECT 49.050 84.140 50.000 84.900 ;
      LAYER li1 ;
        RECT 50.180 84.260 50.430 84.970 ;
      LAYER li1 ;
        RECT 50.610 84.900 50.640 85.070 ;
        RECT 50.810 84.900 51.000 85.070 ;
        RECT 51.170 84.900 51.360 85.070 ;
        RECT 51.530 84.900 51.560 85.070 ;
        RECT 52.170 85.070 53.120 85.100 ;
        RECT 50.610 84.440 51.560 84.900 ;
      LAYER li1 ;
        RECT 51.740 84.260 51.990 84.970 ;
      LAYER li1 ;
        RECT 38.460 82.780 38.790 83.770 ;
      LAYER li1 ;
        RECT 39.490 83.690 40.750 83.920 ;
      LAYER li1 ;
        RECT 42.790 83.910 44.030 84.040 ;
        RECT 40.930 83.870 44.030 83.910 ;
        RECT 40.930 83.740 42.960 83.870 ;
      LAYER li1 ;
        RECT 40.580 83.560 40.750 83.690 ;
        RECT 40.580 83.390 42.470 83.560 ;
      LAYER li1 ;
        RECT 35.770 81.790 35.780 81.960 ;
        RECT 35.950 81.790 36.140 81.960 ;
        RECT 36.310 81.790 36.330 81.960 ;
        RECT 35.770 81.710 36.330 81.790 ;
        RECT 37.690 81.910 39.140 82.780 ;
        RECT 37.690 81.740 37.940 81.910 ;
        RECT 38.110 81.740 38.300 81.910 ;
        RECT 38.470 81.740 38.740 81.910 ;
        RECT 38.910 81.740 39.140 81.910 ;
        RECT 37.690 81.710 39.140 81.740 ;
        RECT 39.450 81.960 40.400 83.290 ;
        RECT 39.450 81.790 39.480 81.960 ;
        RECT 39.650 81.790 39.840 81.960 ;
        RECT 40.010 81.790 40.200 81.960 ;
        RECT 40.370 81.790 40.400 81.960 ;
        RECT 39.450 81.710 40.400 81.790 ;
      LAYER li1 ;
        RECT 40.580 81.710 40.830 83.390 ;
      LAYER li1 ;
        RECT 41.010 81.960 41.960 83.210 ;
        RECT 41.010 81.790 41.040 81.960 ;
        RECT 41.210 81.790 41.400 81.960 ;
        RECT 41.570 81.790 41.760 81.960 ;
        RECT 41.930 81.790 41.960 81.960 ;
        RECT 41.010 81.710 41.960 81.790 ;
      LAYER li1 ;
        RECT 42.140 81.710 42.470 83.390 ;
        RECT 43.250 83.350 43.580 83.690 ;
      LAYER li1 ;
        RECT 42.650 81.960 43.600 83.170 ;
        RECT 42.650 81.790 42.680 81.960 ;
        RECT 42.850 81.790 43.040 81.960 ;
        RECT 43.210 81.790 43.400 81.960 ;
        RECT 43.570 81.790 43.600 81.960 ;
        RECT 42.650 81.710 43.600 81.790 ;
        RECT 43.780 81.710 44.030 83.870 ;
        RECT 44.900 83.440 45.230 84.110 ;
        RECT 45.630 82.790 45.960 83.770 ;
        RECT 46.180 83.440 46.510 84.110 ;
      LAYER li1 ;
        RECT 50.180 84.090 51.990 84.260 ;
      LAYER li1 ;
        RECT 52.170 84.900 52.200 85.070 ;
        RECT 52.370 84.900 52.560 85.070 ;
        RECT 52.730 84.900 52.920 85.070 ;
        RECT 53.090 84.900 53.120 85.070 ;
        RECT 53.930 85.070 55.540 85.100 ;
        RECT 52.170 84.220 53.120 84.900 ;
      LAYER li1 ;
        RECT 50.180 83.920 50.350 84.090 ;
      LAYER li1 ;
        RECT 53.300 84.040 53.630 84.970 ;
        RECT 53.930 84.900 53.980 85.070 ;
        RECT 54.150 84.900 54.420 85.070 ;
        RECT 54.590 84.900 54.860 85.070 ;
        RECT 55.030 84.900 55.270 85.070 ;
        RECT 55.440 84.900 55.540 85.070 ;
        RECT 53.930 84.620 55.540 84.900 ;
        RECT 46.910 82.790 47.240 83.770 ;
      LAYER li1 ;
        RECT 49.090 83.690 50.350 83.920 ;
      LAYER li1 ;
        RECT 52.390 83.910 53.630 84.040 ;
        RECT 50.530 83.870 53.630 83.910 ;
        RECT 50.530 83.740 52.560 83.870 ;
      LAYER li1 ;
        RECT 50.180 83.560 50.350 83.690 ;
        RECT 50.180 83.390 52.070 83.560 ;
      LAYER li1 ;
        RECT 44.660 81.910 47.400 82.790 ;
        RECT 44.660 81.740 44.870 81.910 ;
        RECT 45.040 81.740 45.310 81.910 ;
        RECT 45.480 81.740 45.720 81.910 ;
        RECT 45.890 81.740 46.150 81.910 ;
        RECT 46.320 81.740 46.590 81.910 ;
        RECT 46.760 81.740 47.000 81.910 ;
        RECT 47.170 81.740 47.400 81.910 ;
        RECT 44.660 81.720 47.400 81.740 ;
        RECT 49.050 81.960 50.000 83.290 ;
        RECT 49.050 81.790 49.080 81.960 ;
        RECT 49.250 81.790 49.440 81.960 ;
        RECT 49.610 81.790 49.800 81.960 ;
        RECT 49.970 81.790 50.000 81.960 ;
        RECT 49.050 81.710 50.000 81.790 ;
      LAYER li1 ;
        RECT 50.180 81.710 50.430 83.390 ;
      LAYER li1 ;
        RECT 50.610 81.960 51.560 83.210 ;
        RECT 50.610 81.790 50.640 81.960 ;
        RECT 50.810 81.790 51.000 81.960 ;
        RECT 51.170 81.790 51.360 81.960 ;
        RECT 51.530 81.790 51.560 81.960 ;
        RECT 50.610 81.710 51.560 81.790 ;
      LAYER li1 ;
        RECT 51.740 81.710 52.070 83.390 ;
        RECT 52.850 83.350 53.180 83.690 ;
      LAYER li1 ;
        RECT 52.250 81.960 53.200 83.170 ;
        RECT 52.250 81.790 52.280 81.960 ;
        RECT 52.450 81.790 52.640 81.960 ;
        RECT 52.810 81.790 53.000 81.960 ;
        RECT 53.170 81.790 53.200 81.960 ;
        RECT 52.250 81.710 53.200 81.790 ;
        RECT 53.380 81.710 53.630 83.870 ;
        RECT 54.240 84.220 55.540 84.620 ;
        RECT 55.770 85.070 56.720 85.100 ;
        RECT 55.770 84.900 55.800 85.070 ;
        RECT 55.970 84.900 56.160 85.070 ;
        RECT 56.330 84.900 56.520 85.070 ;
        RECT 56.690 84.900 56.720 85.070 ;
        RECT 57.330 85.070 58.280 85.100 ;
        RECT 54.240 83.440 54.570 84.220 ;
        RECT 55.770 84.140 56.720 84.900 ;
      LAYER li1 ;
        RECT 56.900 84.260 57.150 84.970 ;
      LAYER li1 ;
        RECT 57.330 84.900 57.360 85.070 ;
        RECT 57.530 84.900 57.720 85.070 ;
        RECT 57.890 84.900 58.080 85.070 ;
        RECT 58.250 84.900 58.280 85.070 ;
        RECT 58.890 85.070 59.840 85.100 ;
        RECT 57.330 84.440 58.280 84.900 ;
      LAYER li1 ;
        RECT 58.460 84.260 58.710 84.970 ;
        RECT 56.900 84.090 58.710 84.260 ;
      LAYER li1 ;
        RECT 58.890 84.900 58.920 85.070 ;
        RECT 59.090 84.900 59.280 85.070 ;
        RECT 59.450 84.900 59.640 85.070 ;
        RECT 59.810 84.900 59.840 85.070 ;
        RECT 61.060 85.080 63.790 85.110 ;
        RECT 58.890 84.220 59.840 84.900 ;
      LAYER li1 ;
        RECT 56.900 83.920 57.070 84.090 ;
      LAYER li1 ;
        RECT 60.020 84.040 60.350 84.970 ;
        RECT 61.060 84.910 61.230 85.080 ;
        RECT 61.400 84.910 61.670 85.080 ;
        RECT 61.840 84.910 62.080 85.080 ;
        RECT 62.250 84.910 62.510 85.080 ;
        RECT 62.680 84.910 62.950 85.080 ;
        RECT 63.120 84.910 63.360 85.080 ;
        RECT 63.530 84.910 63.790 85.080 ;
        RECT 65.350 85.070 66.600 85.100 ;
        RECT 67.780 85.080 70.510 85.110 ;
        RECT 61.060 84.110 63.790 84.910 ;
        RECT 54.780 82.780 55.110 83.770 ;
      LAYER li1 ;
        RECT 55.810 83.690 57.070 83.920 ;
      LAYER li1 ;
        RECT 59.110 83.910 60.350 84.040 ;
        RECT 57.250 83.870 60.350 83.910 ;
        RECT 57.250 83.740 59.280 83.870 ;
      LAYER li1 ;
        RECT 56.900 83.560 57.070 83.690 ;
        RECT 56.900 83.390 58.790 83.560 ;
      LAYER li1 ;
        RECT 54.010 81.910 55.460 82.780 ;
        RECT 54.010 81.740 54.260 81.910 ;
        RECT 54.430 81.740 54.620 81.910 ;
        RECT 54.790 81.740 55.060 81.910 ;
        RECT 55.230 81.740 55.460 81.910 ;
        RECT 54.010 81.710 55.460 81.740 ;
        RECT 55.770 81.960 56.720 83.290 ;
        RECT 55.770 81.790 55.800 81.960 ;
        RECT 55.970 81.790 56.160 81.960 ;
        RECT 56.330 81.790 56.520 81.960 ;
        RECT 56.690 81.790 56.720 81.960 ;
        RECT 55.770 81.710 56.720 81.790 ;
      LAYER li1 ;
        RECT 56.900 81.710 57.150 83.390 ;
      LAYER li1 ;
        RECT 57.330 81.960 58.280 83.210 ;
        RECT 57.330 81.790 57.360 81.960 ;
        RECT 57.530 81.790 57.720 81.960 ;
        RECT 57.890 81.790 58.080 81.960 ;
        RECT 58.250 81.790 58.280 81.960 ;
        RECT 57.330 81.710 58.280 81.790 ;
      LAYER li1 ;
        RECT 58.460 81.710 58.790 83.390 ;
        RECT 59.570 83.350 59.900 83.690 ;
      LAYER li1 ;
        RECT 58.970 81.960 59.920 83.170 ;
        RECT 58.970 81.790 59.000 81.960 ;
        RECT 59.170 81.790 59.360 81.960 ;
        RECT 59.530 81.790 59.720 81.960 ;
        RECT 59.890 81.790 59.920 81.960 ;
        RECT 58.970 81.710 59.920 81.790 ;
        RECT 60.100 81.710 60.350 83.870 ;
        RECT 61.220 83.440 61.550 84.110 ;
        RECT 61.950 82.790 62.280 83.770 ;
        RECT 62.500 83.440 62.830 84.110 ;
        RECT 63.230 82.790 63.560 83.770 ;
      LAYER li1 ;
        RECT 64.920 83.290 65.170 84.970 ;
      LAYER li1 ;
        RECT 65.520 84.900 65.710 85.070 ;
        RECT 65.880 84.900 66.070 85.070 ;
        RECT 66.240 84.900 66.430 85.070 ;
        RECT 65.350 84.530 66.600 84.900 ;
        RECT 66.780 84.350 67.030 84.970 ;
        RECT 65.480 84.180 67.030 84.350 ;
        RECT 65.480 83.720 65.810 84.180 ;
        RECT 60.980 81.910 63.720 82.790 ;
        RECT 60.980 81.740 61.190 81.910 ;
        RECT 61.360 81.740 61.630 81.910 ;
        RECT 61.800 81.740 62.040 81.910 ;
        RECT 62.210 81.740 62.470 81.910 ;
        RECT 62.640 81.740 62.910 81.910 ;
        RECT 63.080 81.740 63.320 81.910 ;
        RECT 63.490 81.740 63.720 81.910 ;
        RECT 60.980 81.720 63.720 81.740 ;
      LAYER li1 ;
        RECT 64.920 81.710 65.350 83.290 ;
      LAYER li1 ;
        RECT 65.530 81.960 66.090 83.290 ;
      LAYER li1 ;
        RECT 66.270 82.210 66.600 84.000 ;
      LAYER li1 ;
        RECT 66.780 82.460 67.030 84.180 ;
        RECT 67.780 84.910 67.950 85.080 ;
        RECT 68.120 84.910 68.390 85.080 ;
        RECT 68.560 84.910 68.800 85.080 ;
        RECT 68.970 84.910 69.230 85.080 ;
        RECT 69.400 84.910 69.670 85.080 ;
        RECT 69.840 84.910 70.080 85.080 ;
        RECT 70.250 84.910 70.510 85.080 ;
        RECT 67.780 84.110 70.510 84.910 ;
        RECT 72.090 85.070 73.400 85.100 ;
        RECT 72.090 84.900 72.120 85.070 ;
        RECT 72.290 84.900 72.480 85.070 ;
        RECT 72.650 84.900 72.840 85.070 ;
        RECT 73.010 84.900 73.200 85.070 ;
        RECT 73.370 84.900 73.400 85.070 ;
        RECT 74.570 85.070 76.180 85.100 ;
        RECT 72.090 84.120 73.400 84.900 ;
      LAYER li1 ;
        RECT 73.850 84.290 74.180 84.950 ;
      LAYER li1 ;
        RECT 74.570 84.900 74.620 85.070 ;
        RECT 74.790 84.900 75.060 85.070 ;
        RECT 75.230 84.900 75.500 85.070 ;
        RECT 75.670 84.900 75.910 85.070 ;
        RECT 76.080 84.900 76.180 85.070 ;
        RECT 76.850 85.070 77.710 85.100 ;
        RECT 74.570 84.620 76.180 84.900 ;
      LAYER li1 ;
        RECT 73.580 84.120 74.180 84.290 ;
      LAYER li1 ;
        RECT 74.880 84.220 76.180 84.620 ;
        RECT 67.940 83.440 68.270 84.110 ;
        RECT 68.670 82.790 69.000 83.770 ;
        RECT 69.220 83.440 69.550 84.110 ;
      LAYER li1 ;
        RECT 73.580 83.940 73.800 84.120 ;
      LAYER li1 ;
        RECT 69.950 82.790 70.280 83.770 ;
      LAYER li1 ;
        RECT 72.130 83.530 73.020 83.920 ;
        RECT 73.220 83.770 73.800 83.940 ;
      LAYER li1 ;
        RECT 65.530 81.790 65.540 81.960 ;
        RECT 65.710 81.790 65.900 81.960 ;
        RECT 66.070 81.790 66.090 81.960 ;
        RECT 65.530 81.710 66.090 81.790 ;
        RECT 67.700 81.910 70.440 82.790 ;
        RECT 67.700 81.740 67.910 81.910 ;
        RECT 68.080 81.740 68.350 81.910 ;
        RECT 68.520 81.740 68.760 81.910 ;
        RECT 68.930 81.740 69.190 81.910 ;
        RECT 69.360 81.740 69.630 81.910 ;
        RECT 69.800 81.740 70.040 81.910 ;
        RECT 70.210 81.740 70.440 81.910 ;
        RECT 67.700 81.720 70.440 81.740 ;
        RECT 72.090 81.960 73.040 83.290 ;
        RECT 72.090 81.790 72.120 81.960 ;
        RECT 72.290 81.790 72.480 81.960 ;
        RECT 72.650 81.790 72.840 81.960 ;
        RECT 73.010 81.790 73.040 81.960 ;
        RECT 72.090 81.710 73.040 81.790 ;
      LAYER li1 ;
        RECT 73.220 81.710 73.470 83.770 ;
        RECT 73.980 83.610 74.280 83.940 ;
      LAYER li1 ;
        RECT 74.880 83.440 75.210 84.220 ;
        RECT 76.470 83.910 76.680 84.970 ;
        RECT 76.850 84.900 76.900 85.070 ;
        RECT 77.070 84.900 77.490 85.070 ;
        RECT 77.660 84.900 77.710 85.070 ;
        RECT 78.940 85.070 79.610 85.100 ;
        RECT 76.850 84.560 77.710 84.900 ;
        RECT 77.890 84.560 78.290 84.970 ;
        RECT 78.940 84.900 79.010 85.070 ;
        RECT 79.180 84.900 79.370 85.070 ;
        RECT 79.540 84.900 79.610 85.070 ;
        RECT 80.330 85.070 81.940 85.100 ;
      LAYER li1 ;
        RECT 76.850 84.080 77.640 84.390 ;
      LAYER li1 ;
        RECT 77.890 83.910 78.060 84.560 ;
      LAYER li1 ;
        RECT 78.240 84.080 78.770 84.390 ;
      LAYER li1 ;
        RECT 78.940 84.140 79.610 84.900 ;
        RECT 73.660 81.960 74.250 83.290 ;
        RECT 75.420 82.780 75.750 83.770 ;
        RECT 76.470 83.740 79.580 83.910 ;
        RECT 73.660 81.790 73.690 81.960 ;
        RECT 73.860 81.790 74.050 81.960 ;
        RECT 74.220 81.790 74.250 81.960 ;
        RECT 73.660 81.710 74.250 81.790 ;
        RECT 74.650 81.910 76.100 82.780 ;
        RECT 76.470 82.690 76.720 83.740 ;
      LAYER li1 ;
        RECT 76.930 82.210 77.860 83.560 ;
      LAYER li1 ;
        RECT 79.250 83.530 79.580 83.740 ;
        RECT 78.030 82.040 79.600 83.290 ;
        RECT 74.650 81.740 74.900 81.910 ;
        RECT 75.070 81.740 75.260 81.910 ;
        RECT 75.430 81.740 75.700 81.910 ;
        RECT 75.870 81.740 76.100 81.910 ;
        RECT 74.650 81.710 76.100 81.740 ;
        RECT 77.940 81.960 79.600 82.040 ;
        RECT 77.940 81.790 77.990 81.960 ;
        RECT 78.160 81.790 78.350 81.960 ;
        RECT 78.520 81.790 78.710 81.960 ;
        RECT 78.880 81.790 79.070 81.960 ;
        RECT 79.240 81.790 79.430 81.960 ;
        RECT 77.940 81.710 79.600 81.790 ;
      LAYER li1 ;
        RECT 79.780 81.710 80.040 84.970 ;
      LAYER li1 ;
        RECT 80.330 84.900 80.380 85.070 ;
        RECT 80.550 84.900 80.820 85.070 ;
        RECT 80.990 84.900 81.260 85.070 ;
        RECT 81.430 84.900 81.670 85.070 ;
        RECT 81.840 84.900 81.940 85.070 ;
        RECT 80.330 84.620 81.940 84.900 ;
        RECT 80.640 84.220 81.940 84.620 ;
        RECT 82.170 85.070 82.760 85.100 ;
        RECT 84.220 85.070 85.830 85.100 ;
        RECT 86.090 85.070 87.700 85.100 ;
        RECT 82.170 84.900 82.200 85.070 ;
        RECT 82.370 84.900 82.560 85.070 ;
        RECT 82.730 84.900 82.760 85.070 ;
        RECT 80.640 83.440 80.970 84.220 ;
        RECT 82.170 84.140 82.760 84.900 ;
      LAYER li1 ;
        RECT 83.790 84.660 84.040 84.970 ;
      LAYER li1 ;
        RECT 84.390 84.900 84.580 85.070 ;
        RECT 84.750 84.900 84.940 85.070 ;
        RECT 85.110 84.900 85.300 85.070 ;
        RECT 85.470 84.900 85.660 85.070 ;
        RECT 86.090 84.900 86.140 85.070 ;
        RECT 86.310 84.900 86.580 85.070 ;
        RECT 86.750 84.900 87.020 85.070 ;
        RECT 87.190 84.900 87.430 85.070 ;
        RECT 87.600 84.900 87.700 85.070 ;
      LAYER li1 ;
        RECT 83.170 84.490 84.040 84.660 ;
      LAYER li1 ;
        RECT 81.180 82.780 81.510 83.770 ;
      LAYER li1 ;
        RECT 82.210 83.630 82.920 83.960 ;
        RECT 83.170 83.290 83.370 84.490 ;
        RECT 83.790 84.140 84.040 84.490 ;
      LAYER li1 ;
        RECT 84.220 84.140 85.830 84.900 ;
        RECT 86.090 84.620 87.700 84.900 ;
        RECT 86.400 84.220 87.700 84.620 ;
        RECT 87.930 85.070 88.880 85.100 ;
        RECT 87.930 84.900 87.960 85.070 ;
        RECT 88.130 84.900 88.320 85.070 ;
        RECT 88.490 84.900 88.680 85.070 ;
        RECT 88.850 84.900 88.880 85.070 ;
        RECT 89.490 85.070 90.440 85.100 ;
      LAYER li1 ;
        RECT 84.130 83.720 84.840 83.960 ;
        RECT 85.020 83.720 85.800 83.960 ;
      LAYER li1 ;
        RECT 80.410 81.910 81.860 82.780 ;
        RECT 80.410 81.740 80.660 81.910 ;
        RECT 80.830 81.740 81.020 81.910 ;
        RECT 81.190 81.740 81.460 81.910 ;
        RECT 81.630 81.740 81.860 81.910 ;
        RECT 80.410 81.710 81.860 81.740 ;
        RECT 82.230 81.830 82.560 83.290 ;
      LAYER li1 ;
        RECT 83.010 82.010 83.370 83.290 ;
      LAYER li1 ;
        RECT 83.790 83.370 85.680 83.540 ;
        RECT 86.400 83.440 86.730 84.220 ;
        RECT 87.930 84.140 88.880 84.900 ;
      LAYER li1 ;
        RECT 89.060 84.260 89.310 84.970 ;
      LAYER li1 ;
        RECT 89.490 84.900 89.520 85.070 ;
        RECT 89.690 84.900 89.880 85.070 ;
        RECT 90.050 84.900 90.240 85.070 ;
        RECT 90.410 84.900 90.440 85.070 ;
        RECT 91.050 85.070 92.000 85.100 ;
        RECT 89.490 84.440 90.440 84.900 ;
      LAYER li1 ;
        RECT 90.620 84.260 90.870 84.970 ;
        RECT 89.060 84.090 90.870 84.260 ;
      LAYER li1 ;
        RECT 91.050 84.900 91.080 85.070 ;
        RECT 91.250 84.900 91.440 85.070 ;
        RECT 91.610 84.900 91.800 85.070 ;
        RECT 91.970 84.900 92.000 85.070 ;
        RECT 92.810 85.070 94.420 85.100 ;
        RECT 91.050 84.220 92.000 84.900 ;
      LAYER li1 ;
        RECT 89.060 83.920 89.230 84.090 ;
      LAYER li1 ;
        RECT 92.180 84.040 92.510 84.970 ;
        RECT 92.810 84.900 92.860 85.070 ;
        RECT 93.030 84.900 93.300 85.070 ;
        RECT 93.470 84.900 93.740 85.070 ;
        RECT 93.910 84.900 94.150 85.070 ;
        RECT 94.320 84.900 94.420 85.070 ;
        RECT 92.810 84.620 94.420 84.900 ;
        RECT 83.790 81.830 84.040 83.370 ;
        RECT 82.230 81.660 84.040 81.830 ;
        RECT 84.220 81.960 85.170 83.190 ;
        RECT 84.220 81.790 84.250 81.960 ;
        RECT 84.420 81.790 84.610 81.960 ;
        RECT 84.780 81.790 84.970 81.960 ;
        RECT 85.140 81.790 85.170 81.960 ;
        RECT 84.220 81.710 85.170 81.790 ;
        RECT 85.350 81.710 85.680 83.370 ;
        RECT 86.940 82.780 87.270 83.770 ;
      LAYER li1 ;
        RECT 87.970 83.690 89.230 83.920 ;
      LAYER li1 ;
        RECT 91.270 83.910 92.510 84.040 ;
        RECT 89.410 83.870 92.510 83.910 ;
        RECT 89.410 83.740 91.440 83.870 ;
      LAYER li1 ;
        RECT 89.060 83.560 89.230 83.690 ;
        RECT 89.060 83.390 90.950 83.560 ;
      LAYER li1 ;
        RECT 86.170 81.910 87.620 82.780 ;
        RECT 86.170 81.740 86.420 81.910 ;
        RECT 86.590 81.740 86.780 81.910 ;
        RECT 86.950 81.740 87.220 81.910 ;
        RECT 87.390 81.740 87.620 81.910 ;
        RECT 86.170 81.710 87.620 81.740 ;
        RECT 87.930 81.960 88.880 83.290 ;
        RECT 87.930 81.790 87.960 81.960 ;
        RECT 88.130 81.790 88.320 81.960 ;
        RECT 88.490 81.790 88.680 81.960 ;
        RECT 88.850 81.790 88.880 81.960 ;
        RECT 87.930 81.710 88.880 81.790 ;
      LAYER li1 ;
        RECT 89.060 81.710 89.310 83.390 ;
      LAYER li1 ;
        RECT 89.490 81.960 90.440 83.210 ;
        RECT 89.490 81.790 89.520 81.960 ;
        RECT 89.690 81.790 89.880 81.960 ;
        RECT 90.050 81.790 90.240 81.960 ;
        RECT 90.410 81.790 90.440 81.960 ;
        RECT 89.490 81.710 90.440 81.790 ;
      LAYER li1 ;
        RECT 90.620 81.710 90.950 83.390 ;
        RECT 91.730 83.350 92.060 83.690 ;
      LAYER li1 ;
        RECT 91.130 81.960 92.080 83.170 ;
        RECT 91.130 81.790 91.160 81.960 ;
        RECT 91.330 81.790 91.520 81.960 ;
        RECT 91.690 81.790 91.880 81.960 ;
        RECT 92.050 81.790 92.080 81.960 ;
        RECT 91.130 81.710 92.080 81.790 ;
        RECT 92.260 81.710 92.510 83.870 ;
        RECT 93.120 84.220 94.420 84.620 ;
        RECT 94.650 85.070 95.600 85.100 ;
        RECT 94.650 84.900 94.680 85.070 ;
        RECT 94.850 84.900 95.040 85.070 ;
        RECT 95.210 84.900 95.400 85.070 ;
        RECT 95.570 84.900 95.600 85.070 ;
        RECT 96.210 85.070 97.160 85.100 ;
        RECT 93.120 83.440 93.450 84.220 ;
        RECT 94.650 84.140 95.600 84.900 ;
      LAYER li1 ;
        RECT 95.780 84.260 96.030 84.970 ;
      LAYER li1 ;
        RECT 96.210 84.900 96.240 85.070 ;
        RECT 96.410 84.900 96.600 85.070 ;
        RECT 96.770 84.900 96.960 85.070 ;
        RECT 97.130 84.900 97.160 85.070 ;
        RECT 97.770 85.070 98.720 85.100 ;
        RECT 96.210 84.440 97.160 84.900 ;
      LAYER li1 ;
        RECT 97.340 84.260 97.590 84.970 ;
        RECT 95.780 84.090 97.590 84.260 ;
      LAYER li1 ;
        RECT 97.770 84.900 97.800 85.070 ;
        RECT 97.970 84.900 98.160 85.070 ;
        RECT 98.330 84.900 98.520 85.070 ;
        RECT 98.690 84.900 98.720 85.070 ;
        RECT 99.530 85.070 101.140 85.100 ;
        RECT 97.770 84.220 98.720 84.900 ;
      LAYER li1 ;
        RECT 95.780 83.920 95.950 84.090 ;
      LAYER li1 ;
        RECT 98.900 84.040 99.230 84.970 ;
        RECT 99.530 84.900 99.580 85.070 ;
        RECT 99.750 84.900 100.020 85.070 ;
        RECT 100.190 84.900 100.460 85.070 ;
        RECT 100.630 84.900 100.870 85.070 ;
        RECT 101.040 84.900 101.140 85.070 ;
        RECT 99.530 84.620 101.140 84.900 ;
        RECT 93.660 82.780 93.990 83.770 ;
      LAYER li1 ;
        RECT 94.690 83.690 95.950 83.920 ;
      LAYER li1 ;
        RECT 97.990 83.910 99.230 84.040 ;
        RECT 96.130 83.870 99.230 83.910 ;
        RECT 96.130 83.740 98.160 83.870 ;
      LAYER li1 ;
        RECT 95.780 83.560 95.950 83.690 ;
        RECT 95.780 83.390 97.670 83.560 ;
      LAYER li1 ;
        RECT 92.890 81.910 94.340 82.780 ;
        RECT 92.890 81.740 93.140 81.910 ;
        RECT 93.310 81.740 93.500 81.910 ;
        RECT 93.670 81.740 93.940 81.910 ;
        RECT 94.110 81.740 94.340 81.910 ;
        RECT 92.890 81.710 94.340 81.740 ;
        RECT 94.650 81.960 95.600 83.290 ;
        RECT 94.650 81.790 94.680 81.960 ;
        RECT 94.850 81.790 95.040 81.960 ;
        RECT 95.210 81.790 95.400 81.960 ;
        RECT 95.570 81.790 95.600 81.960 ;
        RECT 94.650 81.710 95.600 81.790 ;
      LAYER li1 ;
        RECT 95.780 81.710 96.030 83.390 ;
      LAYER li1 ;
        RECT 96.210 81.960 97.160 83.210 ;
        RECT 96.210 81.790 96.240 81.960 ;
        RECT 96.410 81.790 96.600 81.960 ;
        RECT 96.770 81.790 96.960 81.960 ;
        RECT 97.130 81.790 97.160 81.960 ;
        RECT 96.210 81.710 97.160 81.790 ;
      LAYER li1 ;
        RECT 97.340 81.710 97.670 83.390 ;
        RECT 98.450 83.350 98.780 83.690 ;
      LAYER li1 ;
        RECT 97.850 81.960 98.800 83.170 ;
        RECT 97.850 81.790 97.880 81.960 ;
        RECT 98.050 81.790 98.240 81.960 ;
        RECT 98.410 81.790 98.600 81.960 ;
        RECT 98.770 81.790 98.800 81.960 ;
        RECT 97.850 81.710 98.800 81.790 ;
        RECT 98.980 81.710 99.230 83.870 ;
        RECT 99.840 84.220 101.140 84.620 ;
        RECT 101.370 85.070 101.960 85.100 ;
        RECT 101.370 84.900 101.400 85.070 ;
        RECT 101.570 84.900 101.760 85.070 ;
        RECT 101.930 84.900 101.960 85.070 ;
        RECT 102.890 85.070 104.500 85.100 ;
        RECT 99.840 83.440 100.170 84.220 ;
        RECT 101.370 84.140 101.960 84.900 ;
        RECT 100.380 82.780 100.710 83.770 ;
      LAYER li1 ;
        RECT 101.410 83.530 102.120 83.920 ;
        RECT 102.300 83.290 102.630 84.970 ;
      LAYER li1 ;
        RECT 102.890 84.900 102.940 85.070 ;
        RECT 103.110 84.900 103.380 85.070 ;
        RECT 103.550 84.900 103.820 85.070 ;
        RECT 103.990 84.900 104.230 85.070 ;
        RECT 104.400 84.900 104.500 85.070 ;
        RECT 105.680 85.070 106.630 85.100 ;
        RECT 102.890 84.620 104.500 84.900 ;
        RECT 103.200 84.220 104.500 84.620 ;
        RECT 103.200 83.440 103.530 84.220 ;
        RECT 99.610 81.910 101.060 82.780 ;
        RECT 99.610 81.740 99.860 81.910 ;
        RECT 100.030 81.740 100.220 81.910 ;
        RECT 100.390 81.740 100.660 81.910 ;
        RECT 100.830 81.740 101.060 81.910 ;
        RECT 99.610 81.710 101.060 81.740 ;
        RECT 101.370 81.960 101.960 83.290 ;
        RECT 101.370 81.790 101.400 81.960 ;
        RECT 101.570 81.790 101.760 81.960 ;
        RECT 101.930 81.790 101.960 81.960 ;
        RECT 101.370 81.710 101.960 81.790 ;
      LAYER li1 ;
        RECT 102.240 81.710 102.630 83.290 ;
      LAYER li1 ;
        RECT 103.740 82.780 104.070 83.770 ;
        RECT 105.230 83.110 105.500 84.970 ;
        RECT 105.680 84.900 105.710 85.070 ;
        RECT 105.880 84.900 106.070 85.070 ;
        RECT 106.240 84.900 106.430 85.070 ;
        RECT 106.600 84.900 106.630 85.070 ;
        RECT 107.320 85.070 107.910 85.100 ;
        RECT 105.680 84.470 106.630 84.900 ;
        RECT 106.810 84.470 107.140 84.970 ;
        RECT 106.360 83.110 106.690 83.610 ;
        RECT 105.230 82.940 106.690 83.110 ;
        RECT 102.970 81.910 104.420 82.780 ;
        RECT 105.230 82.010 105.560 82.940 ;
        RECT 102.970 81.740 103.220 81.910 ;
        RECT 103.390 81.740 103.580 81.910 ;
        RECT 103.750 81.740 104.020 81.910 ;
        RECT 104.190 81.740 104.420 81.910 ;
        RECT 105.750 81.960 106.340 82.740 ;
        RECT 105.750 81.790 105.780 81.960 ;
        RECT 105.950 81.790 106.140 81.960 ;
        RECT 106.310 81.790 106.340 81.960 ;
        RECT 105.750 81.760 106.340 81.790 ;
        RECT 106.520 81.830 106.690 82.940 ;
        RECT 106.870 83.550 107.140 84.470 ;
        RECT 107.320 84.900 107.350 85.070 ;
        RECT 107.520 84.900 107.710 85.070 ;
        RECT 107.880 84.900 107.910 85.070 ;
        RECT 112.280 85.070 113.230 85.100 ;
        RECT 107.320 84.220 107.910 84.900 ;
      LAYER li1 ;
        RECT 108.190 84.840 111.130 85.010 ;
        RECT 108.190 83.850 108.360 84.840 ;
      LAYER li1 ;
        RECT 106.870 83.320 107.400 83.550 ;
        RECT 106.870 82.010 107.120 83.320 ;
      LAYER li1 ;
        RECT 107.820 82.980 108.360 83.850 ;
        RECT 108.540 83.360 108.870 84.660 ;
      LAYER li1 ;
        RECT 109.050 84.140 109.320 84.640 ;
        RECT 109.770 84.390 110.100 84.640 ;
        RECT 109.770 84.220 110.780 84.390 ;
        RECT 109.050 83.150 109.220 84.140 ;
        RECT 110.100 83.550 110.430 84.040 ;
        RECT 109.000 82.980 109.220 83.150 ;
        RECT 109.400 83.320 110.430 83.550 ;
        RECT 110.610 83.990 110.780 84.220 ;
      LAYER li1 ;
        RECT 110.960 84.340 111.130 84.840 ;
      LAYER li1 ;
        RECT 112.280 84.900 112.310 85.070 ;
        RECT 112.480 84.900 112.670 85.070 ;
        RECT 112.840 84.900 113.030 85.070 ;
        RECT 113.200 84.900 113.230 85.070 ;
        RECT 112.280 84.520 113.230 84.900 ;
      LAYER li1 ;
        RECT 113.410 85.030 116.070 85.200 ;
        RECT 113.410 84.340 113.580 85.030 ;
        RECT 110.960 84.170 113.580 84.340 ;
      LAYER li1 ;
        RECT 110.610 83.820 113.230 83.990 ;
        RECT 109.000 82.800 109.170 82.980 ;
        RECT 109.400 82.800 109.570 83.320 ;
        RECT 110.610 83.140 110.780 83.820 ;
      LAYER li1 ;
        RECT 113.410 83.640 113.580 84.170 ;
      LAYER li1 ;
        RECT 107.360 82.630 109.170 82.800 ;
        RECT 107.360 82.010 107.610 82.630 ;
        RECT 107.790 82.280 108.820 82.450 ;
        RECT 107.790 81.830 107.960 82.280 ;
        RECT 102.970 81.710 104.420 81.740 ;
        RECT 106.520 81.660 107.960 81.830 ;
        RECT 108.140 81.960 108.470 82.100 ;
        RECT 108.140 81.790 108.170 81.960 ;
        RECT 108.340 81.790 108.470 81.960 ;
        RECT 108.140 81.760 108.470 81.790 ;
        RECT 108.650 81.830 108.820 82.280 ;
        RECT 109.000 82.010 109.170 82.630 ;
        RECT 109.350 82.470 109.570 82.800 ;
        RECT 109.750 82.970 110.780 83.140 ;
        RECT 110.960 83.290 111.290 83.640 ;
      LAYER li1 ;
        RECT 111.730 83.470 113.580 83.640 ;
      LAYER li1 ;
        RECT 113.760 84.140 114.090 84.850 ;
        RECT 114.550 84.680 115.720 84.850 ;
        RECT 114.550 84.140 114.880 84.680 ;
        RECT 113.760 83.290 114.020 84.140 ;
        RECT 115.090 83.880 115.370 84.380 ;
        RECT 110.960 83.120 114.020 83.290 ;
        RECT 109.750 82.270 109.920 82.970 ;
        RECT 110.610 82.940 110.780 82.970 ;
        RECT 110.100 82.590 110.430 82.790 ;
        RECT 110.610 82.770 112.380 82.940 ;
        RECT 110.100 82.470 111.870 82.590 ;
        RECT 110.220 82.420 111.870 82.470 ;
        RECT 109.700 82.010 110.030 82.270 ;
        RECT 110.220 81.830 110.390 82.420 ;
        RECT 108.650 81.660 110.390 81.830 ;
        RECT 110.570 81.960 111.520 82.240 ;
        RECT 110.570 81.790 110.600 81.960 ;
        RECT 110.770 81.790 110.960 81.960 ;
        RECT 111.130 81.790 111.320 81.960 ;
        RECT 111.490 81.790 111.520 81.960 ;
        RECT 110.570 81.760 111.520 81.790 ;
        RECT 111.700 81.830 111.870 82.420 ;
        RECT 112.050 82.010 112.380 82.770 ;
        RECT 113.690 82.540 114.020 83.120 ;
        RECT 114.200 83.710 115.370 83.880 ;
        RECT 114.200 82.360 114.370 83.710 ;
        RECT 114.750 83.030 115.080 83.530 ;
        RECT 115.550 83.280 115.720 84.680 ;
      LAYER li1 ;
        RECT 115.900 84.370 116.070 85.030 ;
      LAYER li1 ;
        RECT 116.250 85.070 117.200 85.100 ;
        RECT 116.250 84.900 116.280 85.070 ;
        RECT 116.450 84.900 116.640 85.070 ;
        RECT 116.810 84.900 117.000 85.070 ;
        RECT 117.170 84.900 117.200 85.070 ;
        RECT 118.860 85.070 119.810 85.100 ;
        RECT 116.250 84.550 117.200 84.900 ;
        RECT 117.740 84.470 118.070 84.970 ;
        RECT 118.860 84.900 118.890 85.070 ;
        RECT 119.060 84.900 119.250 85.070 ;
        RECT 119.420 84.900 119.610 85.070 ;
        RECT 119.780 84.900 119.810 85.070 ;
      LAYER li1 ;
        RECT 115.900 84.260 116.910 84.370 ;
        RECT 115.900 84.200 116.960 84.260 ;
        RECT 116.580 84.090 116.960 84.200 ;
      LAYER li1 ;
        RECT 115.930 83.630 116.260 84.020 ;
      LAYER li1 ;
        RECT 116.580 83.810 116.910 84.090 ;
      LAYER li1 ;
        RECT 117.740 83.630 117.970 84.470 ;
        RECT 118.350 83.970 118.680 84.470 ;
        RECT 118.860 83.970 119.810 84.900 ;
        RECT 121.060 85.080 123.790 85.110 ;
        RECT 121.060 84.910 121.230 85.080 ;
        RECT 121.400 84.910 121.670 85.080 ;
        RECT 121.840 84.910 122.080 85.080 ;
        RECT 122.250 84.910 122.510 85.080 ;
        RECT 122.680 84.910 122.950 85.080 ;
        RECT 123.120 84.910 123.360 85.080 ;
        RECT 123.530 84.910 123.790 85.080 ;
        RECT 121.060 84.110 123.790 84.910 ;
        RECT 124.900 85.080 127.630 85.110 ;
        RECT 124.900 84.910 125.070 85.080 ;
        RECT 125.240 84.910 125.510 85.080 ;
        RECT 125.680 84.910 125.920 85.080 ;
        RECT 126.090 84.910 126.350 85.080 ;
        RECT 126.520 84.910 126.790 85.080 ;
        RECT 126.960 84.910 127.200 85.080 ;
        RECT 127.370 84.910 127.630 85.080 ;
        RECT 124.900 84.110 127.630 84.910 ;
        RECT 128.740 85.080 131.470 85.110 ;
        RECT 128.740 84.910 128.910 85.080 ;
        RECT 129.080 84.910 129.350 85.080 ;
        RECT 129.520 84.910 129.760 85.080 ;
        RECT 129.930 84.910 130.190 85.080 ;
        RECT 130.360 84.910 130.630 85.080 ;
        RECT 130.800 84.910 131.040 85.080 ;
        RECT 131.210 84.910 131.470 85.080 ;
        RECT 128.740 84.110 131.470 84.910 ;
        RECT 132.580 85.080 135.310 85.110 ;
        RECT 132.580 84.910 132.750 85.080 ;
        RECT 132.920 84.910 133.190 85.080 ;
        RECT 133.360 84.910 133.600 85.080 ;
        RECT 133.770 84.910 134.030 85.080 ;
        RECT 134.200 84.910 134.470 85.080 ;
        RECT 134.640 84.910 134.880 85.080 ;
        RECT 135.050 84.910 135.310 85.080 ;
        RECT 132.580 84.110 135.310 84.910 ;
        RECT 136.420 85.080 139.150 85.110 ;
        RECT 136.420 84.910 136.590 85.080 ;
        RECT 136.760 84.910 137.030 85.080 ;
        RECT 137.200 84.910 137.440 85.080 ;
        RECT 137.610 84.910 137.870 85.080 ;
        RECT 138.040 84.910 138.310 85.080 ;
        RECT 138.480 84.910 138.720 85.080 ;
        RECT 138.890 84.910 139.150 85.080 ;
        RECT 136.420 84.110 139.150 84.910 ;
        RECT 139.850 85.070 141.460 85.100 ;
        RECT 139.850 84.900 139.900 85.070 ;
        RECT 140.070 84.900 140.340 85.070 ;
        RECT 140.510 84.900 140.780 85.070 ;
        RECT 140.950 84.900 141.190 85.070 ;
        RECT 141.360 84.900 141.460 85.070 ;
        RECT 139.850 84.620 141.460 84.900 ;
        RECT 140.160 84.220 141.460 84.620 ;
        RECT 115.930 83.460 117.970 83.630 ;
        RECT 115.260 83.110 117.620 83.280 ;
        RECT 115.260 82.790 115.430 83.110 ;
        RECT 117.800 82.930 117.970 83.460 ;
        RECT 112.560 82.190 114.370 82.360 ;
        RECT 114.550 82.620 115.430 82.790 ;
        RECT 112.560 81.830 112.730 82.190 ;
        RECT 111.700 81.660 112.730 81.830 ;
        RECT 112.910 81.960 113.860 82.010 ;
        RECT 112.910 81.790 112.940 81.960 ;
        RECT 113.110 81.790 113.300 81.960 ;
        RECT 113.470 81.790 113.660 81.960 ;
        RECT 113.830 81.790 113.860 81.960 ;
        RECT 112.910 81.710 113.860 81.790 ;
        RECT 114.550 81.710 114.800 82.620 ;
        RECT 115.610 81.960 116.560 82.790 ;
        RECT 116.960 82.760 117.970 82.930 ;
        RECT 118.470 83.790 118.680 83.970 ;
        RECT 118.470 83.460 119.840 83.790 ;
        RECT 116.960 82.290 117.210 82.760 ;
        RECT 117.390 81.960 118.290 82.580 ;
        RECT 118.470 82.460 118.720 83.460 ;
        RECT 121.220 83.440 121.550 84.110 ;
        RECT 115.610 81.790 115.640 81.960 ;
        RECT 115.810 81.790 116.000 81.960 ;
        RECT 116.170 81.790 116.360 81.960 ;
        RECT 116.530 81.790 116.560 81.960 ;
        RECT 117.560 81.790 117.750 81.960 ;
        RECT 117.920 81.790 118.110 81.960 ;
        RECT 118.280 81.790 118.290 81.960 ;
        RECT 115.610 81.760 116.560 81.790 ;
        RECT 117.390 81.760 118.290 81.790 ;
        RECT 118.900 81.960 119.840 83.270 ;
        RECT 121.950 82.790 122.280 83.770 ;
        RECT 122.500 83.440 122.830 84.110 ;
        RECT 123.230 82.790 123.560 83.770 ;
        RECT 125.060 83.440 125.390 84.110 ;
        RECT 125.790 82.790 126.120 83.770 ;
        RECT 126.340 83.440 126.670 84.110 ;
        RECT 127.070 82.790 127.400 83.770 ;
        RECT 128.900 83.440 129.230 84.110 ;
        RECT 129.630 82.790 129.960 83.770 ;
        RECT 130.180 83.440 130.510 84.110 ;
        RECT 130.910 82.790 131.240 83.770 ;
        RECT 132.740 83.440 133.070 84.110 ;
        RECT 133.470 82.790 133.800 83.770 ;
        RECT 134.020 83.440 134.350 84.110 ;
        RECT 134.750 82.790 135.080 83.770 ;
        RECT 136.580 83.440 136.910 84.110 ;
        RECT 137.310 82.790 137.640 83.770 ;
        RECT 137.860 83.440 138.190 84.110 ;
        RECT 138.590 82.790 138.920 83.770 ;
        RECT 140.160 83.440 140.490 84.220 ;
        RECT 118.900 81.790 118.920 81.960 ;
        RECT 119.090 81.790 119.280 81.960 ;
        RECT 119.450 81.790 119.640 81.960 ;
        RECT 119.810 81.790 119.840 81.960 ;
        RECT 118.900 81.730 119.840 81.790 ;
        RECT 120.980 81.910 123.720 82.790 ;
        RECT 120.980 81.740 121.190 81.910 ;
        RECT 121.360 81.740 121.630 81.910 ;
        RECT 121.800 81.740 122.040 81.910 ;
        RECT 122.210 81.740 122.470 81.910 ;
        RECT 122.640 81.740 122.910 81.910 ;
        RECT 123.080 81.740 123.320 81.910 ;
        RECT 123.490 81.740 123.720 81.910 ;
        RECT 120.980 81.720 123.720 81.740 ;
        RECT 124.820 81.910 127.560 82.790 ;
        RECT 124.820 81.740 125.030 81.910 ;
        RECT 125.200 81.740 125.470 81.910 ;
        RECT 125.640 81.740 125.880 81.910 ;
        RECT 126.050 81.740 126.310 81.910 ;
        RECT 126.480 81.740 126.750 81.910 ;
        RECT 126.920 81.740 127.160 81.910 ;
        RECT 127.330 81.740 127.560 81.910 ;
        RECT 124.820 81.720 127.560 81.740 ;
        RECT 128.660 81.910 131.400 82.790 ;
        RECT 128.660 81.740 128.870 81.910 ;
        RECT 129.040 81.740 129.310 81.910 ;
        RECT 129.480 81.740 129.720 81.910 ;
        RECT 129.890 81.740 130.150 81.910 ;
        RECT 130.320 81.740 130.590 81.910 ;
        RECT 130.760 81.740 131.000 81.910 ;
        RECT 131.170 81.740 131.400 81.910 ;
        RECT 128.660 81.720 131.400 81.740 ;
        RECT 132.500 81.910 135.240 82.790 ;
        RECT 132.500 81.740 132.710 81.910 ;
        RECT 132.880 81.740 133.150 81.910 ;
        RECT 133.320 81.740 133.560 81.910 ;
        RECT 133.730 81.740 133.990 81.910 ;
        RECT 134.160 81.740 134.430 81.910 ;
        RECT 134.600 81.740 134.840 81.910 ;
        RECT 135.010 81.740 135.240 81.910 ;
        RECT 132.500 81.720 135.240 81.740 ;
        RECT 136.340 81.910 139.080 82.790 ;
        RECT 140.700 82.780 141.030 83.770 ;
        RECT 136.340 81.740 136.550 81.910 ;
        RECT 136.720 81.740 136.990 81.910 ;
        RECT 137.160 81.740 137.400 81.910 ;
        RECT 137.570 81.740 137.830 81.910 ;
        RECT 138.000 81.740 138.270 81.910 ;
        RECT 138.440 81.740 138.680 81.910 ;
        RECT 138.850 81.740 139.080 81.910 ;
        RECT 136.340 81.720 139.080 81.740 ;
        RECT 139.930 81.910 141.380 82.780 ;
        RECT 139.930 81.740 140.180 81.910 ;
        RECT 140.350 81.740 140.540 81.910 ;
        RECT 140.710 81.740 140.980 81.910 ;
        RECT 141.150 81.740 141.380 81.910 ;
        RECT 139.930 81.710 141.380 81.740 ;
        RECT 5.760 81.310 5.920 81.490 ;
        RECT 6.090 81.310 6.400 81.490 ;
        RECT 6.570 81.310 6.880 81.490 ;
        RECT 7.050 81.310 7.360 81.490 ;
        RECT 7.530 81.310 7.840 81.490 ;
        RECT 8.010 81.310 8.320 81.490 ;
        RECT 8.490 81.310 8.800 81.490 ;
        RECT 8.970 81.310 9.280 81.490 ;
        RECT 9.450 81.310 9.760 81.490 ;
        RECT 9.930 81.310 10.240 81.490 ;
        RECT 10.410 81.310 10.720 81.490 ;
        RECT 10.890 81.310 11.200 81.490 ;
        RECT 11.370 81.310 11.680 81.490 ;
        RECT 11.850 81.310 12.160 81.490 ;
        RECT 12.330 81.310 12.640 81.490 ;
        RECT 12.810 81.310 13.120 81.490 ;
        RECT 13.290 81.310 13.600 81.490 ;
        RECT 13.770 81.310 14.080 81.490 ;
        RECT 14.250 81.480 14.400 81.490 ;
        RECT 14.880 81.480 15.040 81.490 ;
        RECT 14.250 81.310 14.560 81.480 ;
        RECT 14.730 81.310 15.040 81.480 ;
        RECT 15.210 81.310 15.520 81.490 ;
        RECT 15.690 81.310 16.000 81.490 ;
        RECT 16.170 81.310 16.480 81.490 ;
        RECT 16.650 81.310 16.960 81.490 ;
        RECT 17.130 81.310 17.440 81.490 ;
        RECT 17.610 81.310 17.920 81.490 ;
        RECT 18.090 81.310 18.400 81.490 ;
        RECT 18.570 81.310 18.880 81.490 ;
        RECT 19.050 81.310 19.360 81.490 ;
        RECT 19.530 81.310 19.840 81.490 ;
        RECT 20.010 81.310 20.320 81.490 ;
        RECT 20.490 81.310 20.800 81.490 ;
        RECT 20.970 81.310 21.280 81.490 ;
        RECT 21.450 81.310 21.760 81.490 ;
        RECT 21.930 81.310 22.240 81.490 ;
        RECT 22.410 81.310 22.720 81.490 ;
        RECT 22.890 81.310 23.200 81.490 ;
        RECT 23.370 81.310 23.680 81.490 ;
        RECT 23.850 81.310 24.160 81.490 ;
        RECT 24.330 81.310 24.640 81.490 ;
        RECT 24.810 81.310 25.120 81.490 ;
        RECT 25.290 81.310 25.600 81.490 ;
        RECT 25.770 81.310 26.080 81.490 ;
        RECT 26.250 81.310 26.560 81.490 ;
        RECT 26.730 81.310 27.040 81.490 ;
        RECT 27.210 81.310 27.520 81.490 ;
        RECT 27.690 81.310 28.000 81.490 ;
        RECT 28.170 81.310 28.480 81.490 ;
        RECT 28.650 81.310 28.960 81.490 ;
        RECT 29.130 81.310 29.440 81.490 ;
        RECT 29.610 81.310 29.920 81.490 ;
        RECT 30.090 81.310 30.400 81.490 ;
        RECT 30.570 81.310 30.880 81.490 ;
        RECT 31.050 81.310 31.360 81.490 ;
        RECT 31.530 81.310 31.840 81.490 ;
        RECT 32.010 81.310 32.320 81.490 ;
        RECT 32.490 81.310 32.800 81.490 ;
        RECT 32.970 81.310 33.280 81.490 ;
        RECT 33.450 81.310 33.760 81.490 ;
        RECT 33.930 81.310 34.240 81.490 ;
        RECT 34.410 81.310 34.720 81.490 ;
        RECT 34.890 81.310 35.200 81.490 ;
        RECT 35.370 81.310 35.680 81.490 ;
        RECT 35.850 81.310 36.160 81.490 ;
        RECT 36.330 81.310 36.640 81.490 ;
        RECT 36.810 81.310 37.120 81.490 ;
        RECT 37.290 81.310 37.600 81.490 ;
        RECT 37.770 81.310 38.080 81.490 ;
        RECT 38.250 81.310 38.560 81.490 ;
        RECT 38.730 81.310 39.040 81.490 ;
        RECT 39.210 81.310 39.520 81.490 ;
        RECT 39.690 81.310 40.000 81.490 ;
        RECT 40.170 81.310 40.480 81.490 ;
        RECT 40.650 81.310 40.960 81.490 ;
        RECT 41.130 81.310 41.440 81.490 ;
        RECT 41.610 81.310 41.920 81.490 ;
        RECT 42.090 81.310 42.400 81.490 ;
        RECT 42.570 81.310 42.880 81.490 ;
        RECT 43.050 81.310 43.360 81.490 ;
        RECT 43.530 81.310 43.840 81.490 ;
        RECT 44.010 81.310 44.320 81.490 ;
        RECT 44.490 81.310 44.800 81.490 ;
        RECT 44.970 81.310 45.280 81.490 ;
        RECT 45.450 81.310 45.760 81.490 ;
        RECT 45.930 81.310 46.240 81.490 ;
        RECT 46.410 81.310 46.720 81.490 ;
        RECT 46.890 81.310 47.200 81.490 ;
        RECT 47.370 81.310 47.680 81.490 ;
        RECT 47.850 81.310 48.160 81.490 ;
        RECT 48.330 81.310 48.640 81.490 ;
        RECT 48.810 81.310 49.120 81.490 ;
        RECT 49.290 81.310 49.600 81.490 ;
        RECT 49.770 81.310 50.080 81.490 ;
        RECT 50.250 81.310 50.560 81.490 ;
        RECT 50.730 81.310 51.040 81.490 ;
        RECT 51.210 81.310 51.520 81.490 ;
        RECT 51.690 81.310 52.000 81.490 ;
        RECT 52.170 81.310 52.480 81.490 ;
        RECT 52.650 81.310 52.960 81.490 ;
        RECT 53.130 81.310 53.440 81.490 ;
        RECT 53.610 81.310 53.920 81.490 ;
        RECT 54.090 81.310 54.400 81.490 ;
        RECT 54.570 81.310 54.880 81.490 ;
        RECT 55.050 81.310 55.360 81.490 ;
        RECT 55.530 81.310 55.840 81.490 ;
        RECT 56.010 81.310 56.320 81.490 ;
        RECT 56.490 81.310 56.800 81.490 ;
        RECT 56.970 81.310 57.280 81.490 ;
        RECT 57.450 81.310 57.760 81.490 ;
        RECT 57.930 81.310 58.240 81.490 ;
        RECT 58.410 81.310 58.720 81.490 ;
        RECT 58.890 81.310 59.200 81.490 ;
        RECT 59.370 81.310 59.680 81.490 ;
        RECT 59.850 81.310 60.160 81.490 ;
        RECT 60.330 81.310 60.640 81.490 ;
        RECT 60.810 81.310 61.120 81.490 ;
        RECT 61.290 81.310 61.600 81.490 ;
        RECT 61.770 81.310 62.080 81.490 ;
        RECT 62.250 81.310 62.560 81.490 ;
        RECT 62.730 81.310 63.040 81.490 ;
        RECT 63.210 81.310 63.520 81.490 ;
        RECT 63.690 81.310 64.000 81.490 ;
        RECT 64.170 81.480 64.480 81.490 ;
        RECT 64.650 81.480 64.960 81.490 ;
        RECT 64.170 81.310 64.320 81.480 ;
        RECT 64.800 81.310 64.960 81.480 ;
        RECT 65.130 81.310 65.440 81.490 ;
        RECT 65.610 81.310 65.920 81.490 ;
        RECT 66.090 81.310 66.400 81.490 ;
        RECT 66.570 81.310 66.880 81.490 ;
        RECT 67.050 81.310 67.360 81.490 ;
        RECT 67.530 81.310 67.840 81.490 ;
        RECT 68.010 81.310 68.320 81.490 ;
        RECT 68.490 81.310 68.800 81.490 ;
        RECT 68.970 81.310 69.280 81.490 ;
        RECT 69.450 81.310 69.760 81.490 ;
        RECT 69.930 81.310 70.240 81.490 ;
        RECT 70.410 81.310 70.720 81.490 ;
        RECT 70.890 81.480 71.040 81.490 ;
        RECT 71.520 81.480 71.680 81.490 ;
        RECT 70.890 81.310 71.200 81.480 ;
        RECT 71.370 81.310 71.680 81.480 ;
        RECT 71.850 81.310 72.160 81.490 ;
        RECT 72.330 81.310 72.640 81.490 ;
        RECT 72.810 81.310 73.120 81.490 ;
        RECT 73.290 81.310 73.600 81.490 ;
        RECT 73.770 81.310 74.080 81.490 ;
        RECT 74.250 81.310 74.560 81.490 ;
        RECT 74.730 81.310 75.040 81.490 ;
        RECT 75.210 81.310 75.520 81.490 ;
        RECT 75.690 81.310 76.000 81.490 ;
        RECT 76.170 81.310 76.480 81.490 ;
        RECT 76.650 81.310 76.960 81.490 ;
        RECT 77.130 81.310 77.440 81.490 ;
        RECT 77.610 81.310 77.920 81.490 ;
        RECT 78.090 81.310 78.400 81.490 ;
        RECT 78.570 81.310 78.880 81.490 ;
        RECT 79.050 81.310 79.360 81.490 ;
        RECT 79.530 81.310 79.840 81.490 ;
        RECT 80.010 81.310 80.320 81.490 ;
        RECT 80.490 81.480 80.640 81.490 ;
        RECT 81.120 81.480 81.280 81.490 ;
        RECT 80.490 81.310 80.800 81.480 ;
        RECT 80.970 81.310 81.280 81.480 ;
        RECT 81.450 81.310 81.760 81.490 ;
        RECT 81.930 81.310 82.240 81.490 ;
        RECT 82.410 81.310 82.720 81.490 ;
        RECT 82.890 81.310 83.200 81.490 ;
        RECT 83.370 81.310 83.680 81.490 ;
        RECT 83.850 81.310 84.160 81.490 ;
        RECT 84.330 81.310 84.640 81.490 ;
        RECT 84.810 81.310 85.120 81.490 ;
        RECT 85.290 81.310 85.600 81.490 ;
        RECT 85.770 81.310 86.080 81.490 ;
        RECT 86.250 81.310 86.560 81.490 ;
        RECT 86.730 81.310 87.040 81.490 ;
        RECT 87.210 81.310 87.520 81.490 ;
        RECT 87.690 81.310 88.000 81.490 ;
        RECT 88.170 81.310 88.480 81.490 ;
        RECT 88.650 81.310 88.960 81.490 ;
        RECT 89.130 81.310 89.440 81.490 ;
        RECT 89.610 81.310 89.920 81.490 ;
        RECT 90.090 81.310 90.400 81.490 ;
        RECT 90.570 81.310 90.880 81.490 ;
        RECT 91.050 81.310 91.360 81.490 ;
        RECT 91.530 81.310 91.840 81.490 ;
        RECT 92.010 81.310 92.320 81.490 ;
        RECT 92.490 81.310 92.800 81.490 ;
        RECT 92.970 81.310 93.280 81.490 ;
        RECT 93.450 81.310 93.760 81.490 ;
        RECT 93.930 81.310 94.240 81.490 ;
        RECT 94.410 81.310 94.720 81.490 ;
        RECT 94.890 81.310 95.200 81.490 ;
        RECT 95.370 81.310 95.680 81.490 ;
        RECT 95.850 81.310 96.160 81.490 ;
        RECT 96.330 81.310 96.640 81.490 ;
        RECT 96.810 81.310 97.120 81.490 ;
        RECT 97.290 81.310 97.600 81.490 ;
        RECT 97.770 81.310 98.080 81.490 ;
        RECT 98.250 81.310 98.560 81.490 ;
        RECT 98.730 81.310 99.040 81.490 ;
        RECT 99.210 81.310 99.520 81.490 ;
        RECT 99.690 81.310 100.000 81.490 ;
        RECT 100.170 81.310 100.480 81.490 ;
        RECT 100.650 81.310 100.960 81.490 ;
        RECT 101.130 81.310 101.440 81.490 ;
        RECT 101.610 81.310 101.920 81.490 ;
        RECT 102.090 81.310 102.400 81.490 ;
        RECT 102.570 81.310 102.880 81.490 ;
        RECT 103.050 81.310 103.360 81.490 ;
        RECT 103.530 81.310 103.840 81.490 ;
        RECT 104.010 81.310 104.320 81.490 ;
        RECT 104.490 81.480 104.800 81.490 ;
        RECT 104.970 81.480 105.280 81.490 ;
        RECT 104.490 81.310 104.640 81.480 ;
        RECT 105.120 81.310 105.280 81.480 ;
        RECT 105.450 81.310 105.760 81.490 ;
        RECT 105.930 81.310 106.240 81.490 ;
        RECT 106.410 81.310 106.720 81.490 ;
        RECT 106.890 81.310 107.200 81.490 ;
        RECT 107.370 81.310 107.680 81.490 ;
        RECT 107.850 81.310 108.160 81.490 ;
        RECT 108.330 81.310 108.640 81.490 ;
        RECT 108.810 81.310 109.120 81.490 ;
        RECT 109.290 81.310 109.600 81.490 ;
        RECT 109.770 81.310 110.080 81.490 ;
        RECT 110.250 81.310 110.560 81.490 ;
        RECT 110.730 81.310 111.040 81.490 ;
        RECT 111.210 81.310 111.520 81.490 ;
        RECT 111.690 81.310 112.000 81.490 ;
        RECT 112.170 81.310 112.480 81.490 ;
        RECT 112.650 81.310 112.960 81.490 ;
        RECT 113.130 81.310 113.440 81.490 ;
        RECT 113.610 81.310 113.920 81.490 ;
        RECT 114.090 81.310 114.400 81.490 ;
        RECT 114.570 81.310 114.880 81.490 ;
        RECT 115.050 81.310 115.360 81.490 ;
        RECT 115.530 81.310 115.840 81.490 ;
        RECT 116.010 81.310 116.320 81.490 ;
        RECT 116.490 81.310 116.800 81.490 ;
        RECT 116.970 81.310 117.280 81.490 ;
        RECT 117.450 81.310 117.760 81.490 ;
        RECT 117.930 81.310 118.240 81.490 ;
        RECT 118.410 81.310 118.720 81.490 ;
        RECT 118.890 81.310 119.200 81.490 ;
        RECT 119.370 81.310 119.680 81.490 ;
        RECT 119.850 81.310 120.160 81.490 ;
        RECT 120.330 81.310 120.640 81.490 ;
        RECT 120.810 81.310 121.120 81.490 ;
        RECT 121.290 81.310 121.600 81.490 ;
        RECT 121.770 81.310 122.080 81.490 ;
        RECT 122.250 81.310 122.560 81.490 ;
        RECT 122.730 81.310 123.040 81.490 ;
        RECT 123.210 81.310 123.520 81.490 ;
        RECT 123.690 81.310 124.000 81.490 ;
        RECT 124.170 81.310 124.480 81.490 ;
        RECT 124.650 81.310 124.960 81.490 ;
        RECT 125.130 81.310 125.440 81.490 ;
        RECT 125.610 81.310 125.920 81.490 ;
        RECT 126.090 81.310 126.400 81.490 ;
        RECT 126.570 81.310 126.880 81.490 ;
        RECT 127.050 81.310 127.360 81.490 ;
        RECT 127.530 81.310 127.840 81.490 ;
        RECT 128.010 81.310 128.320 81.490 ;
        RECT 128.490 81.310 128.800 81.490 ;
        RECT 128.970 81.310 129.280 81.490 ;
        RECT 129.450 81.310 129.760 81.490 ;
        RECT 129.930 81.310 130.240 81.490 ;
        RECT 130.410 81.310 130.720 81.490 ;
        RECT 130.890 81.310 131.200 81.490 ;
        RECT 131.370 81.310 131.680 81.490 ;
        RECT 131.850 81.310 132.160 81.490 ;
        RECT 132.330 81.310 132.640 81.490 ;
        RECT 132.810 81.310 133.120 81.490 ;
        RECT 133.290 81.310 133.600 81.490 ;
        RECT 133.770 81.310 134.080 81.490 ;
        RECT 134.250 81.310 134.560 81.490 ;
        RECT 134.730 81.310 135.040 81.490 ;
        RECT 135.210 81.310 135.520 81.490 ;
        RECT 135.690 81.310 136.000 81.490 ;
        RECT 136.170 81.310 136.480 81.490 ;
        RECT 136.650 81.310 136.960 81.490 ;
        RECT 137.130 81.310 137.440 81.490 ;
        RECT 137.610 81.310 137.920 81.490 ;
        RECT 138.090 81.310 138.400 81.490 ;
        RECT 138.570 81.310 138.880 81.490 ;
        RECT 139.050 81.310 139.360 81.490 ;
        RECT 139.530 81.310 139.840 81.490 ;
        RECT 140.010 81.310 140.320 81.490 ;
        RECT 140.490 81.310 140.800 81.490 ;
        RECT 140.970 81.310 141.280 81.490 ;
        RECT 141.450 81.480 141.760 81.490 ;
        RECT 141.930 81.480 142.080 81.490 ;
        RECT 141.450 81.310 141.600 81.480 ;
        RECT 6.260 81.060 9.000 81.080 ;
        RECT 6.260 80.890 6.470 81.060 ;
        RECT 6.640 80.890 6.910 81.060 ;
        RECT 7.080 80.890 7.320 81.060 ;
        RECT 7.490 80.890 7.750 81.060 ;
        RECT 7.920 80.890 8.190 81.060 ;
        RECT 8.360 80.890 8.600 81.060 ;
        RECT 8.770 80.890 9.000 81.060 ;
        RECT 6.260 80.010 9.000 80.890 ;
        RECT 10.100 81.060 12.840 81.080 ;
        RECT 10.100 80.890 10.310 81.060 ;
        RECT 10.480 80.890 10.750 81.060 ;
        RECT 10.920 80.890 11.160 81.060 ;
        RECT 11.330 80.890 11.590 81.060 ;
        RECT 11.760 80.890 12.030 81.060 ;
        RECT 12.200 80.890 12.440 81.060 ;
        RECT 12.610 80.890 12.840 81.060 ;
        RECT 10.100 80.010 12.840 80.890 ;
        RECT 6.500 78.690 6.830 79.360 ;
        RECT 7.230 79.030 7.560 80.010 ;
        RECT 7.780 78.690 8.110 79.360 ;
        RECT 8.510 79.030 8.840 80.010 ;
        RECT 10.340 78.690 10.670 79.360 ;
        RECT 11.070 79.030 11.400 80.010 ;
        RECT 11.620 78.690 11.950 79.360 ;
        RECT 12.350 79.030 12.680 80.010 ;
      LAYER li1 ;
        RECT 15.000 79.510 15.430 81.090 ;
      LAYER li1 ;
        RECT 15.610 81.010 16.170 81.090 ;
        RECT 15.610 80.840 15.620 81.010 ;
        RECT 15.790 80.840 15.980 81.010 ;
        RECT 16.150 80.840 16.170 81.010 ;
        RECT 15.610 79.510 16.170 80.840 ;
        RECT 17.780 81.060 20.520 81.080 ;
        RECT 17.780 80.890 17.990 81.060 ;
        RECT 18.160 80.890 18.430 81.060 ;
        RECT 18.600 80.890 18.840 81.060 ;
        RECT 19.010 80.890 19.270 81.060 ;
        RECT 19.440 80.890 19.710 81.060 ;
        RECT 19.880 80.890 20.120 81.060 ;
        RECT 20.290 80.890 20.520 81.060 ;
        RECT 6.340 77.690 9.070 78.690 ;
        RECT 10.180 77.690 12.910 78.690 ;
      LAYER li1 ;
        RECT 15.000 77.830 15.250 79.510 ;
      LAYER li1 ;
        RECT 15.560 78.620 15.890 79.080 ;
      LAYER li1 ;
        RECT 16.350 78.800 16.680 80.590 ;
      LAYER li1 ;
        RECT 16.860 78.620 17.110 80.340 ;
        RECT 17.780 80.010 20.520 80.890 ;
        RECT 21.370 81.060 22.820 81.090 ;
        RECT 21.370 80.890 21.620 81.060 ;
        RECT 21.790 80.890 21.980 81.060 ;
        RECT 22.150 80.890 22.420 81.060 ;
        RECT 22.590 80.890 22.820 81.060 ;
        RECT 21.370 80.020 22.820 80.890 ;
        RECT 23.670 81.010 24.260 81.040 ;
        RECT 23.670 80.840 23.700 81.010 ;
        RECT 23.870 80.840 24.060 81.010 ;
        RECT 24.230 80.840 24.260 81.010 ;
        RECT 18.020 78.690 18.350 79.360 ;
        RECT 18.750 79.030 19.080 80.010 ;
        RECT 19.300 78.690 19.630 79.360 ;
        RECT 20.030 79.030 20.360 80.010 ;
        RECT 15.560 78.450 17.110 78.620 ;
        RECT 15.430 77.700 16.680 78.270 ;
        RECT 16.860 77.830 17.110 78.450 ;
        RECT 17.860 77.690 20.590 78.690 ;
        RECT 21.600 78.580 21.930 79.360 ;
        RECT 22.140 79.030 22.470 80.020 ;
        RECT 23.150 79.860 23.480 80.790 ;
        RECT 23.670 80.060 24.260 80.840 ;
        RECT 24.440 80.970 25.880 81.140 ;
        RECT 24.440 79.860 24.610 80.970 ;
        RECT 23.150 79.690 24.610 79.860 ;
        RECT 21.600 78.180 22.900 78.580 ;
        RECT 21.290 77.700 22.900 78.180 ;
        RECT 23.150 77.830 23.420 79.690 ;
        RECT 24.280 79.190 24.610 79.690 ;
        RECT 24.790 79.480 25.040 80.790 ;
        RECT 25.280 80.170 25.530 80.790 ;
        RECT 25.710 80.520 25.880 80.970 ;
        RECT 26.060 81.010 26.390 81.040 ;
        RECT 26.060 80.840 26.090 81.010 ;
        RECT 26.260 80.840 26.390 81.010 ;
        RECT 26.060 80.700 26.390 80.840 ;
        RECT 26.570 80.970 28.310 81.140 ;
        RECT 26.570 80.520 26.740 80.970 ;
        RECT 25.710 80.350 26.740 80.520 ;
        RECT 26.920 80.170 27.090 80.790 ;
        RECT 27.620 80.530 27.950 80.790 ;
        RECT 25.280 80.000 27.090 80.170 ;
        RECT 27.270 80.000 27.490 80.330 ;
        RECT 26.920 79.820 27.090 80.000 ;
        RECT 24.790 79.250 25.320 79.480 ;
        RECT 24.790 78.330 25.060 79.250 ;
      LAYER li1 ;
        RECT 25.740 78.950 26.280 79.820 ;
      LAYER li1 ;
        RECT 26.920 79.650 27.140 79.820 ;
        RECT 23.600 77.700 24.550 78.330 ;
        RECT 24.730 77.830 25.060 78.330 ;
        RECT 25.240 77.700 25.830 78.580 ;
      LAYER li1 ;
        RECT 26.110 78.340 26.280 78.950 ;
        RECT 26.070 78.170 26.280 78.340 ;
        RECT 26.110 77.960 26.280 78.170 ;
        RECT 26.460 78.140 26.790 79.440 ;
      LAYER li1 ;
        RECT 26.970 78.660 27.140 79.650 ;
        RECT 27.320 79.480 27.490 80.000 ;
        RECT 27.670 79.830 27.840 80.530 ;
        RECT 28.140 80.380 28.310 80.970 ;
        RECT 28.490 81.010 29.440 81.040 ;
        RECT 28.490 80.840 28.520 81.010 ;
        RECT 28.690 80.840 28.880 81.010 ;
        RECT 29.050 80.840 29.240 81.010 ;
        RECT 29.410 80.840 29.440 81.010 ;
        RECT 28.490 80.560 29.440 80.840 ;
        RECT 29.620 80.970 30.650 81.140 ;
        RECT 29.620 80.380 29.790 80.970 ;
        RECT 28.140 80.330 29.790 80.380 ;
        RECT 28.020 80.210 29.790 80.330 ;
        RECT 28.020 80.010 28.350 80.210 ;
        RECT 29.970 80.030 30.300 80.790 ;
        RECT 30.480 80.610 30.650 80.970 ;
        RECT 30.830 81.010 31.780 81.090 ;
        RECT 30.830 80.840 30.860 81.010 ;
        RECT 31.030 80.840 31.220 81.010 ;
        RECT 31.390 80.840 31.580 81.010 ;
        RECT 31.750 80.840 31.780 81.010 ;
        RECT 30.830 80.790 31.780 80.840 ;
        RECT 30.480 80.440 32.290 80.610 ;
        RECT 28.530 79.860 30.300 80.030 ;
        RECT 28.530 79.830 28.700 79.860 ;
        RECT 27.670 79.660 28.700 79.830 ;
        RECT 31.610 79.680 31.940 80.260 ;
        RECT 27.320 79.250 28.350 79.480 ;
        RECT 28.020 78.760 28.350 79.250 ;
        RECT 28.530 78.980 28.700 79.660 ;
        RECT 28.880 79.510 31.940 79.680 ;
        RECT 28.880 79.160 29.210 79.510 ;
      LAYER li1 ;
        RECT 29.650 79.160 31.500 79.330 ;
      LAYER li1 ;
        RECT 28.530 78.810 31.150 78.980 ;
        RECT 26.970 78.160 27.240 78.660 ;
        RECT 28.530 78.580 28.700 78.810 ;
      LAYER li1 ;
        RECT 31.330 78.630 31.500 79.160 ;
      LAYER li1 ;
        RECT 27.690 78.410 28.700 78.580 ;
      LAYER li1 ;
        RECT 28.880 78.460 31.500 78.630 ;
      LAYER li1 ;
        RECT 27.690 78.160 28.020 78.410 ;
      LAYER li1 ;
        RECT 28.880 77.960 29.050 78.460 ;
        RECT 26.110 77.790 29.050 77.960 ;
      LAYER li1 ;
        RECT 30.200 77.700 31.150 78.280 ;
      LAYER li1 ;
        RECT 31.330 77.770 31.500 78.460 ;
      LAYER li1 ;
        RECT 31.680 78.660 31.940 79.510 ;
        RECT 32.120 79.090 32.290 80.440 ;
        RECT 32.470 80.180 32.720 81.090 ;
        RECT 33.530 81.010 34.480 81.040 ;
        RECT 35.310 81.010 36.210 81.040 ;
        RECT 33.530 80.840 33.560 81.010 ;
        RECT 33.730 80.840 33.920 81.010 ;
        RECT 34.090 80.840 34.280 81.010 ;
        RECT 34.450 80.840 34.480 81.010 ;
        RECT 35.480 80.840 35.670 81.010 ;
        RECT 35.840 80.840 36.030 81.010 ;
        RECT 36.200 80.840 36.210 81.010 ;
        RECT 32.470 80.010 33.350 80.180 ;
        RECT 33.530 80.010 34.480 80.840 ;
        RECT 34.880 80.040 35.130 80.510 ;
        RECT 35.310 80.220 36.210 80.840 ;
        RECT 36.820 81.010 37.760 81.070 ;
        RECT 36.820 80.840 36.840 81.010 ;
        RECT 37.010 80.840 37.200 81.010 ;
        RECT 37.370 80.840 37.560 81.010 ;
        RECT 37.730 80.840 37.760 81.010 ;
        RECT 32.670 79.270 33.000 79.770 ;
        RECT 33.180 79.690 33.350 80.010 ;
        RECT 34.880 79.870 35.890 80.040 ;
        RECT 33.180 79.520 35.540 79.690 ;
        RECT 32.120 78.920 33.290 79.090 ;
        RECT 31.680 77.950 32.010 78.660 ;
        RECT 32.470 78.120 32.800 78.660 ;
        RECT 33.010 78.420 33.290 78.920 ;
        RECT 33.470 78.120 33.640 79.520 ;
        RECT 35.720 79.340 35.890 79.870 ;
        RECT 33.850 79.170 35.890 79.340 ;
        RECT 33.850 78.780 34.180 79.170 ;
      LAYER li1 ;
        RECT 34.500 78.600 34.830 78.990 ;
      LAYER li1 ;
        RECT 32.470 77.950 33.640 78.120 ;
      LAYER li1 ;
        RECT 33.820 78.430 34.830 78.600 ;
        RECT 33.820 77.770 33.990 78.430 ;
      LAYER li1 ;
        RECT 35.660 78.330 35.890 79.170 ;
        RECT 36.390 79.340 36.640 80.340 ;
        RECT 36.820 79.530 37.760 80.840 ;
        RECT 36.390 79.010 37.760 79.340 ;
        RECT 36.390 78.830 36.600 79.010 ;
        RECT 36.270 78.330 36.600 78.830 ;
      LAYER li1 ;
        RECT 31.330 77.600 33.990 77.770 ;
      LAYER li1 ;
        RECT 34.170 77.700 35.120 78.250 ;
        RECT 35.660 77.830 35.990 78.330 ;
        RECT 36.780 77.700 37.730 78.830 ;
      LAYER li1 ;
        RECT 37.940 78.000 38.280 81.070 ;
      LAYER li1 ;
        RECT 38.900 81.060 41.640 81.080 ;
        RECT 38.900 80.890 39.110 81.060 ;
        RECT 39.280 80.890 39.550 81.060 ;
        RECT 39.720 80.890 39.960 81.060 ;
        RECT 40.130 80.890 40.390 81.060 ;
        RECT 40.560 80.890 40.830 81.060 ;
        RECT 41.000 80.890 41.240 81.060 ;
        RECT 41.410 80.890 41.640 81.060 ;
        RECT 38.900 80.010 41.640 80.890 ;
        RECT 42.870 81.010 43.460 81.040 ;
        RECT 42.870 80.840 42.900 81.010 ;
        RECT 43.070 80.840 43.260 81.010 ;
        RECT 43.430 80.840 43.460 81.010 ;
        RECT 39.140 78.690 39.470 79.360 ;
        RECT 39.870 79.030 40.200 80.010 ;
        RECT 40.420 78.690 40.750 79.360 ;
        RECT 41.150 79.030 41.480 80.010 ;
        RECT 42.350 79.860 42.680 80.790 ;
        RECT 42.870 80.060 43.460 80.840 ;
        RECT 43.640 80.970 45.080 81.140 ;
        RECT 43.640 79.860 43.810 80.970 ;
        RECT 42.350 79.690 43.810 79.860 ;
        RECT 38.980 77.690 41.710 78.690 ;
        RECT 42.350 77.830 42.620 79.690 ;
        RECT 43.480 79.190 43.810 79.690 ;
        RECT 43.990 79.480 44.240 80.790 ;
        RECT 44.480 80.170 44.730 80.790 ;
        RECT 44.910 80.520 45.080 80.970 ;
        RECT 45.260 81.010 45.590 81.040 ;
        RECT 45.260 80.840 45.290 81.010 ;
        RECT 45.460 80.840 45.590 81.010 ;
        RECT 45.260 80.700 45.590 80.840 ;
        RECT 45.770 80.970 47.510 81.140 ;
        RECT 45.770 80.520 45.940 80.970 ;
        RECT 44.910 80.350 45.940 80.520 ;
        RECT 46.120 80.170 46.290 80.790 ;
        RECT 46.820 80.530 47.150 80.790 ;
        RECT 44.480 80.000 46.290 80.170 ;
        RECT 46.470 80.000 46.690 80.330 ;
        RECT 46.120 79.820 46.290 80.000 ;
        RECT 43.990 79.250 44.520 79.480 ;
        RECT 43.990 78.330 44.260 79.250 ;
      LAYER li1 ;
        RECT 44.940 78.950 45.480 79.820 ;
      LAYER li1 ;
        RECT 46.120 79.650 46.340 79.820 ;
      LAYER li1 ;
        RECT 45.270 78.910 45.480 78.950 ;
      LAYER li1 ;
        RECT 42.800 77.700 43.750 78.330 ;
        RECT 43.930 77.830 44.260 78.330 ;
        RECT 44.440 77.700 45.030 78.580 ;
      LAYER li1 ;
        RECT 45.310 77.960 45.480 78.910 ;
        RECT 45.660 78.140 45.990 79.440 ;
      LAYER li1 ;
        RECT 46.170 78.660 46.340 79.650 ;
        RECT 46.520 79.480 46.690 80.000 ;
        RECT 46.870 79.830 47.040 80.530 ;
        RECT 47.340 80.380 47.510 80.970 ;
        RECT 47.690 81.010 48.640 81.040 ;
        RECT 47.690 80.840 47.720 81.010 ;
        RECT 47.890 80.840 48.080 81.010 ;
        RECT 48.250 80.840 48.440 81.010 ;
        RECT 48.610 80.840 48.640 81.010 ;
        RECT 47.690 80.560 48.640 80.840 ;
        RECT 48.820 80.970 49.850 81.140 ;
        RECT 48.820 80.380 48.990 80.970 ;
        RECT 47.340 80.330 48.990 80.380 ;
        RECT 47.220 80.210 48.990 80.330 ;
        RECT 47.220 80.010 47.550 80.210 ;
        RECT 49.170 80.030 49.500 80.790 ;
        RECT 49.680 80.610 49.850 80.970 ;
        RECT 50.030 81.010 50.980 81.090 ;
        RECT 50.030 80.840 50.060 81.010 ;
        RECT 50.230 80.840 50.420 81.010 ;
        RECT 50.590 80.840 50.780 81.010 ;
        RECT 50.950 80.840 50.980 81.010 ;
        RECT 50.030 80.790 50.980 80.840 ;
        RECT 49.680 80.440 51.490 80.610 ;
        RECT 47.730 79.860 49.500 80.030 ;
        RECT 47.730 79.830 47.900 79.860 ;
        RECT 46.870 79.660 47.900 79.830 ;
        RECT 50.810 79.680 51.140 80.260 ;
        RECT 46.520 79.250 47.550 79.480 ;
        RECT 47.220 78.760 47.550 79.250 ;
        RECT 47.730 78.980 47.900 79.660 ;
        RECT 48.080 79.510 51.140 79.680 ;
        RECT 48.080 79.160 48.410 79.510 ;
      LAYER li1 ;
        RECT 48.850 79.160 50.700 79.330 ;
      LAYER li1 ;
        RECT 47.730 78.810 50.350 78.980 ;
        RECT 46.170 78.160 46.440 78.660 ;
        RECT 47.730 78.580 47.900 78.810 ;
      LAYER li1 ;
        RECT 50.530 78.630 50.700 79.160 ;
      LAYER li1 ;
        RECT 46.890 78.410 47.900 78.580 ;
      LAYER li1 ;
        RECT 48.080 78.460 50.700 78.630 ;
      LAYER li1 ;
        RECT 46.890 78.160 47.220 78.410 ;
      LAYER li1 ;
        RECT 48.080 77.960 48.250 78.460 ;
        RECT 45.310 77.790 48.250 77.960 ;
      LAYER li1 ;
        RECT 49.400 77.700 50.350 78.280 ;
      LAYER li1 ;
        RECT 50.530 77.770 50.700 78.460 ;
      LAYER li1 ;
        RECT 50.880 78.660 51.140 79.510 ;
        RECT 51.320 79.090 51.490 80.440 ;
        RECT 51.670 80.180 51.920 81.090 ;
        RECT 52.730 81.010 53.680 81.040 ;
        RECT 54.510 81.010 55.410 81.040 ;
        RECT 52.730 80.840 52.760 81.010 ;
        RECT 52.930 80.840 53.120 81.010 ;
        RECT 53.290 80.840 53.480 81.010 ;
        RECT 53.650 80.840 53.680 81.010 ;
        RECT 54.680 80.840 54.870 81.010 ;
        RECT 55.040 80.840 55.230 81.010 ;
        RECT 55.400 80.840 55.410 81.010 ;
        RECT 51.670 80.010 52.550 80.180 ;
        RECT 52.730 80.010 53.680 80.840 ;
        RECT 54.080 80.040 54.330 80.510 ;
        RECT 54.510 80.220 55.410 80.840 ;
        RECT 56.020 81.010 56.960 81.070 ;
        RECT 56.020 80.840 56.040 81.010 ;
        RECT 56.210 80.840 56.400 81.010 ;
        RECT 56.570 80.840 56.760 81.010 ;
        RECT 56.930 80.840 56.960 81.010 ;
        RECT 51.870 79.270 52.200 79.770 ;
        RECT 52.380 79.690 52.550 80.010 ;
        RECT 54.080 79.870 55.090 80.040 ;
        RECT 52.380 79.520 54.740 79.690 ;
        RECT 51.320 78.920 52.490 79.090 ;
        RECT 50.880 77.950 51.210 78.660 ;
        RECT 51.670 78.120 52.000 78.660 ;
        RECT 52.210 78.420 52.490 78.920 ;
        RECT 52.670 78.120 52.840 79.520 ;
        RECT 54.920 79.340 55.090 79.870 ;
        RECT 53.050 79.170 55.090 79.340 ;
        RECT 53.050 78.780 53.380 79.170 ;
      LAYER li1 ;
        RECT 53.700 78.600 54.030 78.990 ;
      LAYER li1 ;
        RECT 51.670 77.950 52.840 78.120 ;
      LAYER li1 ;
        RECT 53.020 78.430 54.030 78.600 ;
        RECT 53.020 77.770 53.190 78.430 ;
      LAYER li1 ;
        RECT 54.860 78.330 55.090 79.170 ;
        RECT 55.590 79.340 55.840 80.340 ;
        RECT 56.020 79.530 56.960 80.840 ;
        RECT 55.590 79.010 56.960 79.340 ;
        RECT 55.590 78.830 55.800 79.010 ;
        RECT 55.470 78.330 55.800 78.830 ;
      LAYER li1 ;
        RECT 50.530 77.600 53.190 77.770 ;
      LAYER li1 ;
        RECT 53.370 77.700 54.320 78.250 ;
        RECT 54.860 77.830 55.190 78.330 ;
        RECT 55.980 77.700 56.930 78.830 ;
      LAYER li1 ;
        RECT 57.140 78.000 57.480 81.070 ;
      LAYER li1 ;
        RECT 58.100 81.060 60.840 81.080 ;
        RECT 58.100 80.890 58.310 81.060 ;
        RECT 58.480 80.890 58.750 81.060 ;
        RECT 58.920 80.890 59.160 81.060 ;
        RECT 59.330 80.890 59.590 81.060 ;
        RECT 59.760 80.890 60.030 81.060 ;
        RECT 60.200 80.890 60.440 81.060 ;
        RECT 60.610 80.890 60.840 81.060 ;
        RECT 58.100 80.010 60.840 80.890 ;
        RECT 61.530 81.010 62.480 81.090 ;
        RECT 61.530 80.840 61.560 81.010 ;
        RECT 61.730 80.840 61.920 81.010 ;
        RECT 62.090 80.840 62.280 81.010 ;
        RECT 62.450 80.840 62.480 81.010 ;
        RECT 58.340 78.690 58.670 79.360 ;
        RECT 59.070 79.030 59.400 80.010 ;
        RECT 59.620 78.690 59.950 79.360 ;
        RECT 60.350 79.030 60.680 80.010 ;
        RECT 61.530 79.510 62.480 80.840 ;
      LAYER li1 ;
        RECT 62.660 79.410 62.910 81.090 ;
      LAYER li1 ;
        RECT 63.090 81.010 64.040 81.090 ;
        RECT 63.090 80.840 63.120 81.010 ;
        RECT 63.290 80.840 63.480 81.010 ;
        RECT 63.650 80.840 63.840 81.010 ;
        RECT 64.010 80.840 64.040 81.010 ;
        RECT 63.090 79.590 64.040 80.840 ;
      LAYER li1 ;
        RECT 64.220 79.410 64.550 81.090 ;
      LAYER li1 ;
        RECT 64.730 81.010 65.680 81.090 ;
        RECT 64.730 80.840 64.760 81.010 ;
        RECT 64.930 80.840 65.120 81.010 ;
        RECT 65.290 80.840 65.480 81.010 ;
        RECT 65.650 80.840 65.680 81.010 ;
        RECT 64.730 79.630 65.680 80.840 ;
      LAYER li1 ;
        RECT 62.660 79.240 64.550 79.410 ;
        RECT 62.660 79.110 62.830 79.240 ;
        RECT 65.330 79.110 65.660 79.450 ;
        RECT 61.570 78.880 62.830 79.110 ;
      LAYER li1 ;
        RECT 63.010 78.930 65.040 79.060 ;
        RECT 65.860 78.930 66.110 81.090 ;
        RECT 66.740 81.060 69.480 81.080 ;
        RECT 66.740 80.890 66.950 81.060 ;
        RECT 67.120 80.890 67.390 81.060 ;
        RECT 67.560 80.890 67.800 81.060 ;
        RECT 67.970 80.890 68.230 81.060 ;
        RECT 68.400 80.890 68.670 81.060 ;
        RECT 68.840 80.890 69.080 81.060 ;
        RECT 69.250 80.890 69.480 81.060 ;
        RECT 66.740 80.010 69.480 80.890 ;
        RECT 63.010 78.890 66.110 78.930 ;
      LAYER li1 ;
        RECT 62.660 78.710 62.830 78.880 ;
      LAYER li1 ;
        RECT 64.870 78.760 66.110 78.890 ;
        RECT 58.180 77.690 60.910 78.690 ;
        RECT 61.530 77.700 62.480 78.660 ;
      LAYER li1 ;
        RECT 62.660 78.540 64.470 78.710 ;
        RECT 62.660 77.830 62.910 78.540 ;
      LAYER li1 ;
        RECT 63.090 77.700 64.040 78.360 ;
      LAYER li1 ;
        RECT 64.220 77.830 64.470 78.540 ;
      LAYER li1 ;
        RECT 64.650 77.700 65.600 78.580 ;
        RECT 65.780 77.830 66.110 78.760 ;
        RECT 66.980 78.690 67.310 79.360 ;
        RECT 67.710 79.030 68.040 80.010 ;
        RECT 68.260 78.690 68.590 79.360 ;
        RECT 68.990 79.030 69.320 80.010 ;
      LAYER li1 ;
        RECT 71.650 79.260 72.020 81.090 ;
      LAYER li1 ;
        RECT 72.200 81.010 72.780 81.090 ;
        RECT 77.300 81.060 80.040 81.080 ;
        RECT 72.200 80.840 72.220 81.010 ;
        RECT 72.390 80.840 72.580 81.010 ;
        RECT 72.750 80.840 72.780 81.010 ;
        RECT 72.200 79.510 72.780 80.840 ;
        RECT 74.930 81.010 76.240 81.040 ;
        RECT 74.930 80.840 74.960 81.010 ;
        RECT 75.130 80.840 75.320 81.010 ;
        RECT 75.490 80.840 75.680 81.010 ;
        RECT 75.850 80.840 76.040 81.010 ;
        RECT 76.210 80.840 76.240 81.010 ;
      LAYER li1 ;
        RECT 72.960 80.430 74.750 80.600 ;
      LAYER li1 ;
        RECT 66.820 77.690 69.550 78.690 ;
      LAYER li1 ;
        RECT 71.650 77.830 71.940 79.260 ;
      LAYER li1 ;
        RECT 72.140 78.860 72.470 79.080 ;
      LAYER li1 ;
        RECT 72.960 79.040 73.290 80.430 ;
        RECT 74.550 80.390 74.750 80.430 ;
      LAYER li1 ;
        RECT 74.070 79.920 74.400 80.250 ;
        RECT 73.470 79.750 74.400 79.920 ;
        RECT 73.470 78.860 73.640 79.750 ;
      LAYER li1 ;
        RECT 74.580 79.640 74.750 80.390 ;
      LAYER li1 ;
        RECT 74.930 79.830 76.240 80.840 ;
        RECT 77.300 80.890 77.510 81.060 ;
        RECT 77.680 80.890 77.950 81.060 ;
        RECT 78.120 80.890 78.360 81.060 ;
        RECT 78.530 80.890 78.790 81.060 ;
        RECT 78.960 80.890 79.230 81.060 ;
        RECT 79.400 80.890 79.640 81.060 ;
        RECT 79.810 80.890 80.040 81.060 ;
      LAYER li1 ;
        RECT 73.820 79.290 74.150 79.570 ;
        RECT 74.580 79.470 76.200 79.640 ;
        RECT 73.820 79.120 74.430 79.290 ;
      LAYER li1 ;
        RECT 72.140 78.690 74.080 78.860 ;
        RECT 72.120 77.700 73.730 78.510 ;
        RECT 73.910 78.250 74.080 78.690 ;
      LAYER li1 ;
        RECT 74.260 78.720 74.430 79.120 ;
        RECT 74.260 78.430 75.210 78.720 ;
      LAYER li1 ;
        RECT 75.390 78.610 75.640 79.110 ;
      LAYER li1 ;
        RECT 75.890 78.880 76.200 79.470 ;
      LAYER li1 ;
        RECT 76.420 78.610 76.670 80.250 ;
        RECT 77.300 80.010 80.040 80.890 ;
        RECT 81.210 81.010 82.160 81.090 ;
        RECT 81.210 80.840 81.240 81.010 ;
        RECT 81.410 80.840 81.600 81.010 ;
        RECT 81.770 80.840 81.960 81.010 ;
        RECT 82.130 80.840 82.160 81.010 ;
        RECT 77.540 78.690 77.870 79.360 ;
        RECT 78.270 79.030 78.600 80.010 ;
        RECT 78.820 78.690 79.150 79.360 ;
        RECT 79.550 79.030 79.880 80.010 ;
        RECT 81.210 79.510 82.160 80.840 ;
      LAYER li1 ;
        RECT 82.340 79.410 82.590 81.090 ;
      LAYER li1 ;
        RECT 82.770 81.010 83.720 81.090 ;
        RECT 82.770 80.840 82.800 81.010 ;
        RECT 82.970 80.840 83.160 81.010 ;
        RECT 83.330 80.840 83.520 81.010 ;
        RECT 83.690 80.840 83.720 81.010 ;
        RECT 82.770 79.590 83.720 80.840 ;
      LAYER li1 ;
        RECT 83.900 79.410 84.230 81.090 ;
      LAYER li1 ;
        RECT 84.410 81.010 85.360 81.090 ;
        RECT 84.410 80.840 84.440 81.010 ;
        RECT 84.610 80.840 84.800 81.010 ;
        RECT 84.970 80.840 85.160 81.010 ;
        RECT 85.330 80.840 85.360 81.010 ;
        RECT 84.410 79.630 85.360 80.840 ;
      LAYER li1 ;
        RECT 82.340 79.240 84.230 79.410 ;
        RECT 82.340 79.110 82.510 79.240 ;
        RECT 85.010 79.110 85.340 79.450 ;
        RECT 81.250 78.880 82.510 79.110 ;
      LAYER li1 ;
        RECT 82.690 78.930 84.720 79.060 ;
        RECT 85.540 78.930 85.790 81.090 ;
        RECT 86.170 81.060 87.620 81.090 ;
        RECT 86.170 80.890 86.420 81.060 ;
        RECT 86.590 80.890 86.780 81.060 ;
        RECT 86.950 80.890 87.220 81.060 ;
        RECT 87.390 80.890 87.620 81.060 ;
        RECT 86.170 80.020 87.620 80.890 ;
        RECT 87.930 81.010 88.880 81.090 ;
        RECT 87.930 80.840 87.960 81.010 ;
        RECT 88.130 80.840 88.320 81.010 ;
        RECT 88.490 80.840 88.680 81.010 ;
        RECT 88.850 80.840 88.880 81.010 ;
        RECT 82.690 78.890 85.790 78.930 ;
      LAYER li1 ;
        RECT 82.340 78.710 82.510 78.880 ;
      LAYER li1 ;
        RECT 84.550 78.760 85.790 78.890 ;
        RECT 75.390 78.440 76.670 78.610 ;
        RECT 73.910 77.830 74.400 78.250 ;
        RECT 74.580 77.700 76.240 78.250 ;
        RECT 76.420 77.830 76.670 78.440 ;
        RECT 77.380 77.690 80.110 78.690 ;
        RECT 81.210 77.700 82.160 78.660 ;
      LAYER li1 ;
        RECT 82.340 78.540 84.150 78.710 ;
        RECT 82.340 77.830 82.590 78.540 ;
      LAYER li1 ;
        RECT 82.770 77.700 83.720 78.360 ;
      LAYER li1 ;
        RECT 83.900 77.830 84.150 78.540 ;
      LAYER li1 ;
        RECT 84.330 77.700 85.280 78.580 ;
        RECT 85.460 77.830 85.790 78.760 ;
        RECT 86.400 78.580 86.730 79.360 ;
        RECT 86.940 79.030 87.270 80.020 ;
        RECT 87.930 79.510 88.880 80.840 ;
      LAYER li1 ;
        RECT 89.060 79.410 89.310 81.090 ;
      LAYER li1 ;
        RECT 89.490 81.010 90.440 81.090 ;
        RECT 89.490 80.840 89.520 81.010 ;
        RECT 89.690 80.840 89.880 81.010 ;
        RECT 90.050 80.840 90.240 81.010 ;
        RECT 90.410 80.840 90.440 81.010 ;
        RECT 89.490 79.590 90.440 80.840 ;
      LAYER li1 ;
        RECT 90.620 79.410 90.950 81.090 ;
      LAYER li1 ;
        RECT 91.130 81.010 92.080 81.090 ;
        RECT 91.130 80.840 91.160 81.010 ;
        RECT 91.330 80.840 91.520 81.010 ;
        RECT 91.690 80.840 91.880 81.010 ;
        RECT 92.050 80.840 92.080 81.010 ;
        RECT 91.130 79.630 92.080 80.840 ;
      LAYER li1 ;
        RECT 89.060 79.240 90.950 79.410 ;
        RECT 89.060 79.110 89.230 79.240 ;
        RECT 91.730 79.110 92.060 79.450 ;
        RECT 87.970 78.880 89.230 79.110 ;
      LAYER li1 ;
        RECT 89.410 78.930 91.440 79.060 ;
        RECT 92.260 78.930 92.510 81.090 ;
        RECT 92.890 81.060 94.340 81.090 ;
        RECT 92.890 80.890 93.140 81.060 ;
        RECT 93.310 80.890 93.500 81.060 ;
        RECT 93.670 80.890 93.940 81.060 ;
        RECT 94.110 80.890 94.340 81.060 ;
        RECT 95.390 81.010 97.360 81.090 ;
        RECT 92.890 80.020 94.340 80.890 ;
        RECT 95.560 80.840 95.750 81.010 ;
        RECT 95.920 80.840 96.110 81.010 ;
        RECT 96.280 80.840 96.470 81.010 ;
        RECT 96.640 80.840 96.830 81.010 ;
        RECT 97.000 80.840 97.190 81.010 ;
        RECT 89.410 78.890 92.510 78.930 ;
      LAYER li1 ;
        RECT 89.060 78.710 89.230 78.880 ;
      LAYER li1 ;
        RECT 91.270 78.760 92.510 78.890 ;
        RECT 86.400 78.180 87.700 78.580 ;
        RECT 86.090 77.700 87.700 78.180 ;
        RECT 87.930 77.700 88.880 78.660 ;
      LAYER li1 ;
        RECT 89.060 78.540 90.870 78.710 ;
        RECT 89.060 77.830 89.310 78.540 ;
      LAYER li1 ;
        RECT 89.490 77.700 90.440 78.360 ;
      LAYER li1 ;
        RECT 90.620 77.830 90.870 78.540 ;
      LAYER li1 ;
        RECT 91.050 77.700 92.000 78.580 ;
        RECT 92.180 77.830 92.510 78.760 ;
        RECT 93.120 78.580 93.450 79.360 ;
        RECT 93.660 79.030 93.990 80.020 ;
        RECT 94.960 79.410 95.210 80.010 ;
        RECT 95.390 79.590 97.360 80.840 ;
        RECT 94.960 79.240 97.340 79.410 ;
        RECT 93.120 78.180 94.420 78.580 ;
      LAYER li1 ;
        RECT 95.170 78.510 95.500 79.060 ;
      LAYER li1 ;
        RECT 95.740 78.330 95.910 79.240 ;
        RECT 97.010 79.060 97.340 79.240 ;
      LAYER li1 ;
        RECT 96.090 78.510 96.420 79.060 ;
      LAYER li1 ;
        RECT 92.810 77.700 94.420 78.180 ;
        RECT 94.650 77.700 95.560 78.330 ;
        RECT 95.740 77.830 96.070 78.330 ;
        RECT 96.600 77.700 97.190 78.660 ;
      LAYER li1 ;
        RECT 97.540 77.830 97.800 81.090 ;
      LAYER li1 ;
        RECT 98.170 81.060 99.620 81.090 ;
        RECT 98.170 80.890 98.420 81.060 ;
        RECT 98.590 80.890 98.780 81.060 ;
        RECT 98.950 80.890 99.220 81.060 ;
        RECT 99.390 80.890 99.620 81.060 ;
        RECT 100.670 81.010 102.640 81.090 ;
        RECT 98.170 80.020 99.620 80.890 ;
        RECT 100.840 80.840 101.030 81.010 ;
        RECT 101.200 80.840 101.390 81.010 ;
        RECT 101.560 80.840 101.750 81.010 ;
        RECT 101.920 80.840 102.110 81.010 ;
        RECT 102.280 80.840 102.470 81.010 ;
        RECT 98.400 78.580 98.730 79.360 ;
        RECT 98.940 79.030 99.270 80.020 ;
        RECT 100.240 79.410 100.490 80.010 ;
        RECT 100.670 79.590 102.640 80.840 ;
        RECT 100.240 79.240 102.620 79.410 ;
        RECT 98.400 78.180 99.700 78.580 ;
      LAYER li1 ;
        RECT 100.450 78.510 100.780 79.060 ;
      LAYER li1 ;
        RECT 101.020 78.330 101.190 79.240 ;
        RECT 102.290 79.060 102.620 79.240 ;
      LAYER li1 ;
        RECT 101.370 78.510 101.700 79.060 ;
      LAYER li1 ;
        RECT 98.090 77.700 99.700 78.180 ;
        RECT 99.930 77.700 100.840 78.330 ;
        RECT 101.020 77.830 101.350 78.330 ;
        RECT 101.880 77.700 102.470 78.660 ;
      LAYER li1 ;
        RECT 102.820 77.830 103.080 81.090 ;
      LAYER li1 ;
        RECT 103.450 81.060 104.900 81.090 ;
        RECT 103.450 80.890 103.700 81.060 ;
        RECT 103.870 80.890 104.060 81.060 ;
        RECT 104.230 80.890 104.500 81.060 ;
        RECT 104.670 80.890 104.900 81.060 ;
        RECT 105.950 81.010 107.920 81.090 ;
        RECT 103.450 80.020 104.900 80.890 ;
        RECT 106.120 80.840 106.310 81.010 ;
        RECT 106.480 80.840 106.670 81.010 ;
        RECT 106.840 80.840 107.030 81.010 ;
        RECT 107.200 80.840 107.390 81.010 ;
        RECT 107.560 80.840 107.750 81.010 ;
        RECT 103.680 78.580 104.010 79.360 ;
        RECT 104.220 79.030 104.550 80.020 ;
        RECT 105.520 79.410 105.770 80.010 ;
        RECT 105.950 79.590 107.920 80.840 ;
        RECT 105.520 79.240 107.900 79.410 ;
        RECT 103.680 78.180 104.980 78.580 ;
      LAYER li1 ;
        RECT 105.730 78.510 106.060 79.060 ;
      LAYER li1 ;
        RECT 106.300 78.330 106.470 79.240 ;
        RECT 107.570 79.060 107.900 79.240 ;
      LAYER li1 ;
        RECT 106.650 78.510 106.980 79.060 ;
      LAYER li1 ;
        RECT 103.370 77.700 104.980 78.180 ;
        RECT 105.210 77.700 106.120 78.330 ;
        RECT 106.300 77.830 106.630 78.330 ;
        RECT 107.160 77.700 107.750 78.660 ;
      LAYER li1 ;
        RECT 108.100 77.830 108.360 81.090 ;
      LAYER li1 ;
        RECT 108.730 81.060 110.180 81.090 ;
        RECT 108.730 80.890 108.980 81.060 ;
        RECT 109.150 80.890 109.340 81.060 ;
        RECT 109.510 80.890 109.780 81.060 ;
        RECT 109.950 80.890 110.180 81.060 ;
        RECT 108.730 80.020 110.180 80.890 ;
        RECT 108.960 78.580 109.290 79.360 ;
        RECT 109.500 79.030 109.830 80.020 ;
      LAYER li1 ;
        RECT 110.520 79.510 110.950 81.090 ;
      LAYER li1 ;
        RECT 111.130 81.010 111.690 81.090 ;
        RECT 111.130 80.840 111.140 81.010 ;
        RECT 111.310 80.840 111.500 81.010 ;
        RECT 111.670 80.840 111.690 81.010 ;
        RECT 111.130 79.510 111.690 80.840 ;
        RECT 113.050 81.060 114.500 81.090 ;
        RECT 113.050 80.890 113.300 81.060 ;
        RECT 113.470 80.890 113.660 81.060 ;
        RECT 113.830 80.890 114.100 81.060 ;
        RECT 114.270 80.890 114.500 81.060 ;
        RECT 108.960 78.180 110.260 78.580 ;
        RECT 108.650 77.700 110.260 78.180 ;
      LAYER li1 ;
        RECT 110.520 77.830 110.770 79.510 ;
      LAYER li1 ;
        RECT 111.080 78.620 111.410 79.080 ;
      LAYER li1 ;
        RECT 111.870 78.800 112.200 80.590 ;
      LAYER li1 ;
        RECT 112.380 78.620 112.630 80.340 ;
        RECT 113.050 80.020 114.500 80.890 ;
        RECT 111.080 78.450 112.630 78.620 ;
        RECT 110.950 77.700 112.200 78.270 ;
        RECT 112.380 77.830 112.630 78.450 ;
        RECT 113.280 78.580 113.610 79.360 ;
        RECT 113.820 79.030 114.150 80.020 ;
      LAYER li1 ;
        RECT 114.840 79.510 115.270 81.090 ;
      LAYER li1 ;
        RECT 115.450 81.010 116.010 81.090 ;
        RECT 115.450 80.840 115.460 81.010 ;
        RECT 115.630 80.840 115.820 81.010 ;
        RECT 115.990 80.840 116.010 81.010 ;
        RECT 115.450 79.510 116.010 80.840 ;
        RECT 117.370 81.060 118.820 81.090 ;
        RECT 117.370 80.890 117.620 81.060 ;
        RECT 117.790 80.890 117.980 81.060 ;
        RECT 118.150 80.890 118.420 81.060 ;
        RECT 118.590 80.890 118.820 81.060 ;
        RECT 113.280 78.180 114.580 78.580 ;
        RECT 112.970 77.700 114.580 78.180 ;
      LAYER li1 ;
        RECT 114.840 77.830 115.090 79.510 ;
      LAYER li1 ;
        RECT 115.400 78.620 115.730 79.080 ;
      LAYER li1 ;
        RECT 116.190 78.800 116.520 80.590 ;
      LAYER li1 ;
        RECT 116.700 78.620 116.950 80.340 ;
        RECT 117.370 80.020 118.820 80.890 ;
        RECT 115.400 78.450 116.950 78.620 ;
        RECT 115.270 77.700 116.520 78.270 ;
        RECT 116.700 77.830 116.950 78.450 ;
        RECT 117.600 78.580 117.930 79.360 ;
        RECT 118.140 79.030 118.470 80.020 ;
      LAYER li1 ;
        RECT 119.160 79.510 119.590 81.090 ;
      LAYER li1 ;
        RECT 119.770 81.010 120.330 81.090 ;
        RECT 119.770 80.840 119.780 81.010 ;
        RECT 119.950 80.840 120.140 81.010 ;
        RECT 120.310 80.840 120.330 81.010 ;
        RECT 119.770 79.510 120.330 80.840 ;
        RECT 121.690 81.060 123.140 81.090 ;
        RECT 121.690 80.890 121.940 81.060 ;
        RECT 122.110 80.890 122.300 81.060 ;
        RECT 122.470 80.890 122.740 81.060 ;
        RECT 122.910 80.890 123.140 81.060 ;
        RECT 117.600 78.180 118.900 78.580 ;
        RECT 117.290 77.700 118.900 78.180 ;
      LAYER li1 ;
        RECT 119.160 77.830 119.410 79.510 ;
      LAYER li1 ;
        RECT 119.720 78.620 120.050 79.080 ;
      LAYER li1 ;
        RECT 120.510 78.800 120.840 80.590 ;
      LAYER li1 ;
        RECT 121.020 78.620 121.270 80.340 ;
        RECT 121.690 80.020 123.140 80.890 ;
        RECT 119.720 78.450 121.270 78.620 ;
        RECT 119.590 77.700 120.840 78.270 ;
        RECT 121.020 77.830 121.270 78.450 ;
        RECT 121.920 78.580 122.250 79.360 ;
        RECT 122.460 79.030 122.790 80.020 ;
      LAYER li1 ;
        RECT 123.480 79.510 123.910 81.090 ;
      LAYER li1 ;
        RECT 124.090 81.010 124.650 81.090 ;
        RECT 124.090 80.840 124.100 81.010 ;
        RECT 124.270 80.840 124.460 81.010 ;
        RECT 124.630 80.840 124.650 81.010 ;
        RECT 124.090 79.510 124.650 80.840 ;
        RECT 126.260 81.060 129.000 81.080 ;
        RECT 126.260 80.890 126.470 81.060 ;
        RECT 126.640 80.890 126.910 81.060 ;
        RECT 127.080 80.890 127.320 81.060 ;
        RECT 127.490 80.890 127.750 81.060 ;
        RECT 127.920 80.890 128.190 81.060 ;
        RECT 128.360 80.890 128.600 81.060 ;
        RECT 128.770 80.890 129.000 81.060 ;
        RECT 121.920 78.180 123.220 78.580 ;
        RECT 121.610 77.700 123.220 78.180 ;
      LAYER li1 ;
        RECT 123.480 77.830 123.730 79.510 ;
      LAYER li1 ;
        RECT 124.040 78.620 124.370 79.080 ;
      LAYER li1 ;
        RECT 124.830 78.800 125.160 80.590 ;
      LAYER li1 ;
        RECT 125.340 78.620 125.590 80.340 ;
        RECT 126.260 80.010 129.000 80.890 ;
        RECT 130.100 81.060 132.840 81.080 ;
        RECT 130.100 80.890 130.310 81.060 ;
        RECT 130.480 80.890 130.750 81.060 ;
        RECT 130.920 80.890 131.160 81.060 ;
        RECT 131.330 80.890 131.590 81.060 ;
        RECT 131.760 80.890 132.030 81.060 ;
        RECT 132.200 80.890 132.440 81.060 ;
        RECT 132.610 80.890 132.840 81.060 ;
        RECT 130.100 80.010 132.840 80.890 ;
        RECT 133.940 81.060 136.680 81.080 ;
        RECT 133.940 80.890 134.150 81.060 ;
        RECT 134.320 80.890 134.590 81.060 ;
        RECT 134.760 80.890 135.000 81.060 ;
        RECT 135.170 80.890 135.430 81.060 ;
        RECT 135.600 80.890 135.870 81.060 ;
        RECT 136.040 80.890 136.280 81.060 ;
        RECT 136.450 80.890 136.680 81.060 ;
        RECT 133.940 80.010 136.680 80.890 ;
        RECT 137.780 81.060 140.520 81.080 ;
        RECT 137.780 80.890 137.990 81.060 ;
        RECT 138.160 80.890 138.430 81.060 ;
        RECT 138.600 80.890 138.840 81.060 ;
        RECT 139.010 80.890 139.270 81.060 ;
        RECT 139.440 80.890 139.710 81.060 ;
        RECT 139.880 80.890 140.120 81.060 ;
        RECT 140.290 80.890 140.520 81.060 ;
        RECT 137.780 80.010 140.520 80.890 ;
        RECT 126.500 78.690 126.830 79.360 ;
        RECT 127.230 79.030 127.560 80.010 ;
        RECT 127.780 78.690 128.110 79.360 ;
        RECT 128.510 79.030 128.840 80.010 ;
        RECT 130.340 78.690 130.670 79.360 ;
        RECT 131.070 79.030 131.400 80.010 ;
        RECT 131.620 78.690 131.950 79.360 ;
        RECT 132.350 79.030 132.680 80.010 ;
        RECT 134.180 78.690 134.510 79.360 ;
        RECT 134.910 79.030 135.240 80.010 ;
        RECT 135.460 78.690 135.790 79.360 ;
        RECT 136.190 79.030 136.520 80.010 ;
        RECT 138.020 78.690 138.350 79.360 ;
        RECT 138.750 79.030 139.080 80.010 ;
        RECT 139.300 78.690 139.630 79.360 ;
        RECT 140.030 79.030 140.360 80.010 ;
        RECT 124.040 78.450 125.590 78.620 ;
        RECT 123.910 77.700 125.160 78.270 ;
        RECT 125.340 77.830 125.590 78.450 ;
        RECT 126.340 77.690 129.070 78.690 ;
        RECT 130.180 77.690 132.910 78.690 ;
        RECT 134.020 77.690 136.750 78.690 ;
        RECT 137.860 77.690 140.590 78.690 ;
        RECT 5.760 77.240 5.920 77.420 ;
        RECT 6.090 77.240 6.400 77.420 ;
        RECT 6.570 77.240 6.880 77.420 ;
        RECT 7.050 77.240 7.360 77.420 ;
        RECT 7.530 77.240 7.840 77.420 ;
        RECT 8.010 77.240 8.320 77.420 ;
        RECT 8.490 77.240 8.800 77.420 ;
        RECT 8.970 77.240 9.280 77.420 ;
        RECT 9.450 77.240 9.760 77.420 ;
        RECT 9.930 77.240 10.240 77.420 ;
        RECT 10.410 77.240 10.720 77.420 ;
        RECT 10.890 77.240 11.200 77.420 ;
        RECT 11.370 77.240 11.680 77.420 ;
        RECT 11.850 77.240 12.160 77.420 ;
        RECT 12.330 77.240 12.640 77.420 ;
        RECT 12.810 77.240 13.120 77.420 ;
        RECT 13.290 77.240 13.600 77.420 ;
        RECT 13.770 77.240 14.080 77.420 ;
        RECT 14.250 77.240 14.400 77.420 ;
        RECT 14.880 77.240 15.040 77.420 ;
        RECT 15.210 77.240 15.520 77.420 ;
        RECT 15.690 77.240 16.000 77.420 ;
        RECT 16.170 77.240 16.480 77.420 ;
        RECT 16.650 77.240 16.960 77.420 ;
        RECT 17.130 77.240 17.440 77.420 ;
        RECT 17.610 77.240 17.920 77.420 ;
        RECT 18.090 77.240 18.400 77.420 ;
        RECT 18.570 77.240 18.880 77.420 ;
        RECT 19.050 77.240 19.360 77.420 ;
        RECT 19.530 77.240 19.840 77.420 ;
        RECT 20.010 77.240 20.320 77.420 ;
        RECT 20.490 77.240 20.800 77.420 ;
        RECT 20.970 77.240 21.280 77.420 ;
        RECT 21.450 77.240 21.760 77.420 ;
        RECT 21.930 77.240 22.240 77.420 ;
        RECT 22.410 77.240 22.720 77.420 ;
        RECT 22.890 77.240 23.200 77.420 ;
        RECT 23.370 77.240 23.680 77.420 ;
        RECT 23.850 77.240 24.160 77.420 ;
        RECT 24.330 77.240 24.640 77.420 ;
        RECT 24.810 77.240 25.120 77.420 ;
        RECT 25.290 77.240 25.600 77.420 ;
        RECT 25.770 77.240 26.080 77.420 ;
        RECT 26.250 77.240 26.560 77.420 ;
        RECT 26.730 77.240 27.040 77.420 ;
        RECT 27.210 77.240 27.520 77.420 ;
        RECT 27.690 77.240 28.000 77.420 ;
        RECT 28.170 77.240 28.480 77.420 ;
        RECT 28.650 77.240 28.960 77.420 ;
        RECT 29.130 77.240 29.440 77.420 ;
        RECT 29.610 77.240 29.920 77.420 ;
        RECT 30.090 77.240 30.400 77.420 ;
        RECT 30.570 77.240 30.880 77.420 ;
        RECT 31.050 77.240 31.360 77.420 ;
        RECT 31.530 77.240 31.840 77.420 ;
        RECT 32.010 77.240 32.320 77.420 ;
        RECT 32.490 77.240 32.800 77.420 ;
        RECT 32.970 77.240 33.280 77.420 ;
        RECT 33.450 77.240 33.760 77.420 ;
        RECT 33.930 77.240 34.240 77.420 ;
        RECT 34.410 77.240 34.720 77.420 ;
        RECT 34.890 77.240 35.200 77.420 ;
        RECT 35.370 77.240 35.680 77.420 ;
        RECT 35.850 77.240 36.160 77.420 ;
        RECT 36.330 77.240 36.640 77.420 ;
        RECT 36.810 77.240 37.120 77.420 ;
        RECT 37.290 77.240 37.600 77.420 ;
        RECT 37.770 77.240 38.080 77.420 ;
        RECT 38.250 77.240 38.560 77.420 ;
        RECT 38.730 77.240 39.040 77.420 ;
        RECT 39.210 77.240 39.520 77.420 ;
        RECT 39.690 77.240 40.000 77.420 ;
        RECT 40.170 77.240 40.480 77.420 ;
        RECT 40.650 77.240 40.960 77.420 ;
        RECT 41.130 77.240 41.440 77.420 ;
        RECT 41.610 77.240 41.920 77.420 ;
        RECT 42.090 77.240 42.400 77.420 ;
        RECT 42.570 77.240 42.880 77.420 ;
        RECT 43.050 77.240 43.360 77.420 ;
        RECT 43.530 77.240 43.840 77.420 ;
        RECT 44.010 77.240 44.320 77.420 ;
        RECT 44.490 77.240 44.800 77.420 ;
        RECT 44.970 77.240 45.280 77.420 ;
        RECT 45.450 77.240 45.760 77.420 ;
        RECT 45.930 77.240 46.240 77.420 ;
        RECT 46.410 77.240 46.720 77.420 ;
        RECT 46.890 77.240 47.200 77.420 ;
        RECT 47.370 77.240 47.680 77.420 ;
        RECT 47.850 77.240 48.160 77.420 ;
        RECT 48.330 77.240 48.640 77.420 ;
        RECT 48.810 77.240 49.120 77.420 ;
        RECT 49.290 77.240 49.600 77.420 ;
        RECT 49.770 77.240 50.080 77.420 ;
        RECT 50.250 77.240 50.560 77.420 ;
        RECT 50.730 77.240 51.040 77.420 ;
        RECT 51.210 77.240 51.520 77.420 ;
        RECT 51.690 77.240 52.000 77.420 ;
        RECT 52.170 77.240 52.480 77.420 ;
        RECT 52.650 77.240 52.960 77.420 ;
        RECT 53.130 77.240 53.440 77.420 ;
        RECT 53.610 77.240 53.920 77.420 ;
        RECT 54.090 77.240 54.400 77.420 ;
        RECT 54.570 77.240 54.880 77.420 ;
        RECT 55.050 77.240 55.360 77.420 ;
        RECT 55.530 77.240 55.840 77.420 ;
        RECT 56.010 77.240 56.320 77.420 ;
        RECT 56.490 77.240 56.800 77.420 ;
        RECT 56.970 77.240 57.280 77.420 ;
        RECT 57.450 77.240 57.760 77.420 ;
        RECT 57.930 77.240 58.240 77.420 ;
        RECT 58.410 77.240 58.720 77.420 ;
        RECT 58.890 77.240 59.200 77.420 ;
        RECT 59.370 77.240 59.680 77.420 ;
        RECT 59.850 77.240 60.160 77.420 ;
        RECT 60.330 77.240 60.640 77.420 ;
        RECT 60.810 77.240 61.120 77.420 ;
        RECT 61.290 77.240 61.600 77.420 ;
        RECT 61.770 77.240 62.080 77.420 ;
        RECT 62.250 77.240 62.560 77.420 ;
        RECT 62.730 77.240 63.040 77.420 ;
        RECT 63.210 77.240 63.520 77.420 ;
        RECT 63.690 77.240 64.000 77.420 ;
        RECT 64.170 77.240 64.480 77.420 ;
        RECT 64.650 77.240 64.960 77.420 ;
        RECT 65.130 77.240 65.440 77.420 ;
        RECT 65.610 77.240 65.920 77.420 ;
        RECT 66.090 77.240 66.400 77.420 ;
        RECT 66.570 77.240 66.880 77.420 ;
        RECT 67.050 77.240 67.360 77.420 ;
        RECT 67.530 77.240 67.840 77.420 ;
        RECT 68.010 77.240 68.320 77.420 ;
        RECT 68.490 77.240 68.800 77.420 ;
        RECT 68.970 77.240 69.280 77.420 ;
        RECT 69.450 77.240 69.760 77.420 ;
        RECT 69.930 77.240 70.240 77.420 ;
        RECT 70.410 77.240 70.720 77.420 ;
        RECT 70.890 77.240 71.040 77.420 ;
        RECT 71.520 77.240 71.680 77.420 ;
        RECT 71.850 77.240 72.160 77.420 ;
        RECT 72.330 77.240 72.640 77.420 ;
        RECT 72.810 77.240 73.120 77.420 ;
        RECT 73.290 77.240 73.600 77.420 ;
        RECT 73.770 77.240 74.080 77.420 ;
        RECT 74.250 77.240 74.560 77.420 ;
        RECT 74.730 77.240 75.040 77.420 ;
        RECT 75.210 77.240 75.520 77.420 ;
        RECT 75.690 77.240 76.000 77.420 ;
        RECT 76.170 77.240 76.480 77.420 ;
        RECT 76.650 77.240 76.960 77.420 ;
        RECT 77.130 77.240 77.440 77.420 ;
        RECT 77.610 77.240 77.920 77.420 ;
        RECT 78.090 77.240 78.400 77.420 ;
        RECT 78.570 77.240 78.880 77.420 ;
        RECT 79.050 77.240 79.360 77.420 ;
        RECT 79.530 77.240 79.840 77.420 ;
        RECT 80.010 77.240 80.320 77.420 ;
        RECT 80.490 77.240 80.640 77.420 ;
        RECT 81.120 77.240 81.280 77.420 ;
        RECT 81.450 77.240 81.760 77.420 ;
        RECT 81.930 77.240 82.240 77.420 ;
        RECT 82.410 77.240 82.720 77.420 ;
        RECT 82.890 77.240 83.200 77.420 ;
        RECT 83.370 77.240 83.680 77.420 ;
        RECT 83.850 77.240 84.160 77.420 ;
        RECT 84.330 77.240 84.640 77.420 ;
        RECT 84.810 77.240 85.120 77.420 ;
        RECT 85.290 77.240 85.600 77.420 ;
        RECT 85.770 77.240 86.080 77.420 ;
        RECT 86.250 77.240 86.560 77.420 ;
        RECT 86.730 77.240 87.040 77.420 ;
        RECT 87.210 77.240 87.520 77.420 ;
        RECT 87.690 77.240 88.000 77.420 ;
        RECT 88.170 77.240 88.480 77.420 ;
        RECT 88.650 77.240 88.960 77.420 ;
        RECT 89.130 77.240 89.440 77.420 ;
        RECT 89.610 77.240 89.920 77.420 ;
        RECT 90.090 77.240 90.400 77.420 ;
        RECT 90.570 77.240 90.880 77.420 ;
        RECT 91.050 77.240 91.360 77.420 ;
        RECT 91.530 77.240 91.840 77.420 ;
        RECT 92.010 77.240 92.320 77.420 ;
        RECT 92.490 77.240 92.800 77.420 ;
        RECT 92.970 77.240 93.280 77.420 ;
        RECT 93.450 77.240 93.760 77.420 ;
        RECT 93.930 77.240 94.240 77.420 ;
        RECT 94.410 77.240 94.720 77.420 ;
        RECT 94.890 77.240 95.200 77.420 ;
        RECT 95.370 77.240 95.680 77.420 ;
        RECT 95.850 77.240 96.160 77.420 ;
        RECT 96.330 77.240 96.640 77.420 ;
        RECT 96.810 77.240 97.120 77.420 ;
        RECT 97.290 77.240 97.600 77.420 ;
        RECT 97.770 77.240 98.080 77.420 ;
        RECT 98.250 77.240 98.560 77.420 ;
        RECT 98.730 77.240 99.040 77.420 ;
        RECT 99.210 77.240 99.520 77.420 ;
        RECT 99.690 77.240 100.000 77.420 ;
        RECT 100.170 77.240 100.480 77.420 ;
        RECT 100.650 77.240 100.960 77.420 ;
        RECT 101.130 77.240 101.440 77.420 ;
        RECT 101.610 77.240 101.920 77.420 ;
        RECT 102.090 77.240 102.400 77.420 ;
        RECT 102.570 77.240 102.880 77.420 ;
        RECT 103.050 77.240 103.360 77.420 ;
        RECT 103.530 77.240 103.840 77.420 ;
        RECT 104.010 77.240 104.320 77.420 ;
        RECT 104.490 77.240 104.800 77.420 ;
        RECT 104.970 77.240 105.280 77.420 ;
        RECT 105.450 77.240 105.760 77.420 ;
        RECT 105.930 77.240 106.240 77.420 ;
        RECT 106.410 77.240 106.720 77.420 ;
        RECT 106.890 77.240 107.200 77.420 ;
        RECT 107.370 77.240 107.680 77.420 ;
        RECT 107.850 77.240 108.160 77.420 ;
        RECT 108.330 77.240 108.640 77.420 ;
        RECT 108.810 77.240 109.120 77.420 ;
        RECT 109.290 77.240 109.600 77.420 ;
        RECT 109.770 77.240 110.080 77.420 ;
        RECT 110.250 77.240 110.560 77.420 ;
        RECT 110.730 77.240 111.040 77.420 ;
        RECT 111.210 77.240 111.520 77.420 ;
        RECT 111.690 77.240 112.000 77.420 ;
        RECT 112.170 77.240 112.480 77.420 ;
        RECT 112.650 77.240 112.960 77.420 ;
        RECT 113.130 77.240 113.440 77.420 ;
        RECT 113.610 77.240 113.920 77.420 ;
        RECT 114.090 77.240 114.400 77.420 ;
        RECT 114.570 77.240 114.880 77.420 ;
        RECT 115.050 77.240 115.360 77.420 ;
        RECT 115.530 77.240 115.840 77.420 ;
        RECT 116.010 77.240 116.320 77.420 ;
        RECT 116.490 77.240 116.800 77.420 ;
        RECT 116.970 77.240 117.280 77.420 ;
        RECT 117.450 77.240 117.760 77.420 ;
        RECT 117.930 77.240 118.240 77.420 ;
        RECT 118.410 77.240 118.720 77.420 ;
        RECT 118.890 77.240 119.200 77.420 ;
        RECT 119.370 77.240 119.680 77.420 ;
        RECT 119.850 77.240 120.160 77.420 ;
        RECT 120.330 77.240 120.640 77.420 ;
        RECT 120.810 77.240 121.120 77.420 ;
        RECT 121.290 77.240 121.600 77.420 ;
        RECT 121.770 77.240 122.080 77.420 ;
        RECT 122.250 77.240 122.560 77.420 ;
        RECT 122.730 77.240 123.040 77.420 ;
        RECT 123.210 77.240 123.520 77.420 ;
        RECT 123.690 77.240 124.000 77.420 ;
        RECT 124.170 77.240 124.480 77.420 ;
        RECT 124.650 77.240 124.960 77.420 ;
        RECT 125.130 77.240 125.440 77.420 ;
        RECT 125.610 77.240 125.920 77.420 ;
        RECT 126.090 77.240 126.400 77.420 ;
        RECT 126.570 77.240 126.880 77.420 ;
        RECT 127.050 77.240 127.360 77.420 ;
        RECT 127.530 77.240 127.840 77.420 ;
        RECT 128.010 77.240 128.320 77.420 ;
        RECT 128.490 77.240 128.800 77.420 ;
        RECT 128.970 77.240 129.280 77.420 ;
        RECT 129.450 77.240 129.760 77.420 ;
        RECT 129.930 77.240 130.240 77.420 ;
        RECT 130.410 77.240 130.720 77.420 ;
        RECT 130.890 77.240 131.200 77.420 ;
        RECT 131.370 77.240 131.680 77.420 ;
        RECT 131.850 77.240 132.160 77.420 ;
        RECT 132.330 77.240 132.640 77.420 ;
        RECT 132.810 77.240 133.120 77.420 ;
        RECT 133.290 77.240 133.600 77.420 ;
        RECT 133.770 77.240 134.080 77.420 ;
        RECT 134.250 77.240 134.560 77.420 ;
        RECT 134.730 77.240 135.040 77.420 ;
        RECT 135.210 77.240 135.520 77.420 ;
        RECT 135.690 77.240 136.000 77.420 ;
        RECT 136.170 77.240 136.480 77.420 ;
        RECT 136.650 77.240 136.960 77.420 ;
        RECT 137.130 77.240 137.440 77.420 ;
        RECT 137.610 77.240 137.920 77.420 ;
        RECT 138.090 77.240 138.400 77.420 ;
        RECT 138.570 77.240 138.880 77.420 ;
        RECT 139.050 77.240 139.360 77.420 ;
        RECT 139.530 77.240 139.840 77.420 ;
        RECT 140.010 77.240 140.320 77.420 ;
        RECT 140.490 77.240 140.800 77.420 ;
        RECT 140.970 77.240 141.280 77.420 ;
        RECT 141.450 77.240 141.760 77.420 ;
        RECT 141.930 77.240 142.080 77.420 ;
        RECT 6.340 76.940 9.070 76.970 ;
        RECT 6.340 76.770 6.510 76.940 ;
        RECT 6.680 76.770 6.950 76.940 ;
        RECT 7.120 76.770 7.360 76.940 ;
        RECT 7.530 76.770 7.790 76.940 ;
        RECT 7.960 76.770 8.230 76.940 ;
        RECT 8.400 76.770 8.640 76.940 ;
        RECT 8.810 76.770 9.070 76.940 ;
        RECT 6.340 75.970 9.070 76.770 ;
        RECT 10.180 76.940 12.910 76.970 ;
        RECT 10.180 76.770 10.350 76.940 ;
        RECT 10.520 76.770 10.790 76.940 ;
        RECT 10.960 76.770 11.200 76.940 ;
        RECT 11.370 76.770 11.630 76.940 ;
        RECT 11.800 76.770 12.070 76.940 ;
        RECT 12.240 76.770 12.480 76.940 ;
        RECT 12.650 76.770 12.910 76.940 ;
        RECT 10.180 75.970 12.910 76.770 ;
        RECT 14.020 76.940 16.750 76.970 ;
        RECT 14.020 76.770 14.190 76.940 ;
        RECT 14.360 76.770 14.630 76.940 ;
        RECT 14.800 76.770 15.040 76.940 ;
        RECT 15.210 76.770 15.470 76.940 ;
        RECT 15.640 76.770 15.910 76.940 ;
        RECT 16.080 76.770 16.320 76.940 ;
        RECT 16.490 76.770 16.750 76.940 ;
        RECT 17.830 76.930 19.080 76.960 ;
        RECT 19.850 76.930 21.460 76.960 ;
        RECT 22.150 76.930 23.400 76.960 ;
        RECT 24.170 76.930 25.780 76.960 ;
        RECT 14.020 75.970 16.750 76.770 ;
        RECT 6.500 75.300 6.830 75.970 ;
        RECT 7.230 74.650 7.560 75.630 ;
        RECT 7.780 75.300 8.110 75.970 ;
        RECT 8.510 74.650 8.840 75.630 ;
        RECT 10.340 75.300 10.670 75.970 ;
        RECT 11.070 74.650 11.400 75.630 ;
        RECT 11.620 75.300 11.950 75.970 ;
        RECT 12.350 74.650 12.680 75.630 ;
        RECT 14.180 75.300 14.510 75.970 ;
        RECT 14.910 74.650 15.240 75.630 ;
        RECT 15.460 75.300 15.790 75.970 ;
        RECT 16.190 74.650 16.520 75.630 ;
      LAYER li1 ;
        RECT 17.400 75.150 17.650 76.830 ;
      LAYER li1 ;
        RECT 18.000 76.760 18.190 76.930 ;
        RECT 18.360 76.760 18.550 76.930 ;
        RECT 18.720 76.760 18.910 76.930 ;
        RECT 17.830 76.390 19.080 76.760 ;
        RECT 19.260 76.210 19.510 76.830 ;
        RECT 19.850 76.760 19.900 76.930 ;
        RECT 20.070 76.760 20.340 76.930 ;
        RECT 20.510 76.760 20.780 76.930 ;
        RECT 20.950 76.760 21.190 76.930 ;
        RECT 21.360 76.760 21.460 76.930 ;
        RECT 19.850 76.480 21.460 76.760 ;
        RECT 17.960 76.040 19.510 76.210 ;
        RECT 17.960 75.580 18.290 76.040 ;
        RECT 6.260 73.770 9.000 74.650 ;
        RECT 6.260 73.600 6.470 73.770 ;
        RECT 6.640 73.600 6.910 73.770 ;
        RECT 7.080 73.600 7.320 73.770 ;
        RECT 7.490 73.600 7.750 73.770 ;
        RECT 7.920 73.600 8.190 73.770 ;
        RECT 8.360 73.600 8.600 73.770 ;
        RECT 8.770 73.600 9.000 73.770 ;
        RECT 6.260 73.580 9.000 73.600 ;
        RECT 10.100 73.770 12.840 74.650 ;
        RECT 10.100 73.600 10.310 73.770 ;
        RECT 10.480 73.600 10.750 73.770 ;
        RECT 10.920 73.600 11.160 73.770 ;
        RECT 11.330 73.600 11.590 73.770 ;
        RECT 11.760 73.600 12.030 73.770 ;
        RECT 12.200 73.600 12.440 73.770 ;
        RECT 12.610 73.600 12.840 73.770 ;
        RECT 10.100 73.580 12.840 73.600 ;
        RECT 13.940 73.770 16.680 74.650 ;
        RECT 13.940 73.600 14.150 73.770 ;
        RECT 14.320 73.600 14.590 73.770 ;
        RECT 14.760 73.600 15.000 73.770 ;
        RECT 15.170 73.600 15.430 73.770 ;
        RECT 15.600 73.600 15.870 73.770 ;
        RECT 16.040 73.600 16.280 73.770 ;
        RECT 16.450 73.600 16.680 73.770 ;
        RECT 13.940 73.580 16.680 73.600 ;
      LAYER li1 ;
        RECT 17.400 73.570 17.830 75.150 ;
      LAYER li1 ;
        RECT 18.010 73.820 18.570 75.150 ;
      LAYER li1 ;
        RECT 18.750 74.070 19.080 75.860 ;
      LAYER li1 ;
        RECT 19.260 74.320 19.510 76.040 ;
        RECT 20.160 76.080 21.460 76.480 ;
        RECT 20.160 75.300 20.490 76.080 ;
        RECT 20.700 74.640 21.030 75.630 ;
      LAYER li1 ;
        RECT 21.720 75.150 21.970 76.830 ;
      LAYER li1 ;
        RECT 22.320 76.760 22.510 76.930 ;
        RECT 22.680 76.760 22.870 76.930 ;
        RECT 23.040 76.760 23.230 76.930 ;
        RECT 22.150 76.390 23.400 76.760 ;
        RECT 23.580 76.210 23.830 76.830 ;
        RECT 24.170 76.760 24.220 76.930 ;
        RECT 24.390 76.760 24.660 76.930 ;
        RECT 24.830 76.760 25.100 76.930 ;
        RECT 25.270 76.760 25.510 76.930 ;
        RECT 25.680 76.760 25.780 76.930 ;
        RECT 24.170 76.480 25.780 76.760 ;
        RECT 22.280 76.040 23.830 76.210 ;
        RECT 22.280 75.580 22.610 76.040 ;
        RECT 18.010 73.650 18.020 73.820 ;
        RECT 18.190 73.650 18.380 73.820 ;
        RECT 18.550 73.650 18.570 73.820 ;
        RECT 18.010 73.570 18.570 73.650 ;
        RECT 19.930 73.770 21.380 74.640 ;
        RECT 19.930 73.600 20.180 73.770 ;
        RECT 20.350 73.600 20.540 73.770 ;
        RECT 20.710 73.600 20.980 73.770 ;
        RECT 21.150 73.600 21.380 73.770 ;
        RECT 19.930 73.570 21.380 73.600 ;
      LAYER li1 ;
        RECT 21.720 73.570 22.150 75.150 ;
      LAYER li1 ;
        RECT 22.330 73.820 22.890 75.150 ;
      LAYER li1 ;
        RECT 23.070 74.070 23.400 75.860 ;
      LAYER li1 ;
        RECT 23.580 74.320 23.830 76.040 ;
        RECT 24.480 76.080 25.780 76.480 ;
        RECT 26.010 76.930 26.960 76.960 ;
        RECT 26.010 76.760 26.040 76.930 ;
        RECT 26.210 76.760 26.400 76.930 ;
        RECT 26.570 76.760 26.760 76.930 ;
        RECT 26.930 76.760 26.960 76.930 ;
        RECT 27.570 76.930 28.520 76.960 ;
        RECT 24.480 75.300 24.810 76.080 ;
        RECT 26.010 76.000 26.960 76.760 ;
      LAYER li1 ;
        RECT 27.140 76.120 27.390 76.830 ;
      LAYER li1 ;
        RECT 27.570 76.760 27.600 76.930 ;
        RECT 27.770 76.760 27.960 76.930 ;
        RECT 28.130 76.760 28.320 76.930 ;
        RECT 28.490 76.760 28.520 76.930 ;
        RECT 29.130 76.930 30.080 76.960 ;
        RECT 27.570 76.300 28.520 76.760 ;
      LAYER li1 ;
        RECT 28.700 76.120 28.950 76.830 ;
        RECT 27.140 75.950 28.950 76.120 ;
      LAYER li1 ;
        RECT 29.130 76.760 29.160 76.930 ;
        RECT 29.330 76.760 29.520 76.930 ;
        RECT 29.690 76.760 29.880 76.930 ;
        RECT 30.050 76.760 30.080 76.930 ;
        RECT 30.890 76.930 32.500 76.960 ;
        RECT 29.130 76.080 30.080 76.760 ;
      LAYER li1 ;
        RECT 27.140 75.780 27.310 75.950 ;
      LAYER li1 ;
        RECT 30.260 75.900 30.590 76.830 ;
        RECT 30.890 76.760 30.940 76.930 ;
        RECT 31.110 76.760 31.380 76.930 ;
        RECT 31.550 76.760 31.820 76.930 ;
        RECT 31.990 76.760 32.230 76.930 ;
        RECT 32.400 76.760 32.500 76.930 ;
        RECT 30.890 76.480 32.500 76.760 ;
        RECT 25.020 74.640 25.350 75.630 ;
      LAYER li1 ;
        RECT 26.050 75.550 27.310 75.780 ;
      LAYER li1 ;
        RECT 29.350 75.770 30.590 75.900 ;
        RECT 27.490 75.730 30.590 75.770 ;
        RECT 27.490 75.600 29.520 75.730 ;
      LAYER li1 ;
        RECT 27.140 75.420 27.310 75.550 ;
        RECT 27.140 75.250 29.030 75.420 ;
      LAYER li1 ;
        RECT 22.330 73.650 22.340 73.820 ;
        RECT 22.510 73.650 22.700 73.820 ;
        RECT 22.870 73.650 22.890 73.820 ;
        RECT 22.330 73.570 22.890 73.650 ;
        RECT 24.250 73.770 25.700 74.640 ;
        RECT 24.250 73.600 24.500 73.770 ;
        RECT 24.670 73.600 24.860 73.770 ;
        RECT 25.030 73.600 25.300 73.770 ;
        RECT 25.470 73.600 25.700 73.770 ;
        RECT 24.250 73.570 25.700 73.600 ;
        RECT 26.010 73.820 26.960 75.150 ;
        RECT 26.010 73.650 26.040 73.820 ;
        RECT 26.210 73.650 26.400 73.820 ;
        RECT 26.570 73.650 26.760 73.820 ;
        RECT 26.930 73.650 26.960 73.820 ;
        RECT 26.010 73.570 26.960 73.650 ;
      LAYER li1 ;
        RECT 27.140 73.570 27.390 75.250 ;
      LAYER li1 ;
        RECT 27.570 73.820 28.520 75.070 ;
        RECT 27.570 73.650 27.600 73.820 ;
        RECT 27.770 73.650 27.960 73.820 ;
        RECT 28.130 73.650 28.320 73.820 ;
        RECT 28.490 73.650 28.520 73.820 ;
        RECT 27.570 73.570 28.520 73.650 ;
      LAYER li1 ;
        RECT 28.700 73.570 29.030 75.250 ;
        RECT 29.810 75.210 30.140 75.550 ;
      LAYER li1 ;
        RECT 29.210 73.820 30.160 75.030 ;
        RECT 29.210 73.650 29.240 73.820 ;
        RECT 29.410 73.650 29.600 73.820 ;
        RECT 29.770 73.650 29.960 73.820 ;
        RECT 30.130 73.650 30.160 73.820 ;
        RECT 29.210 73.570 30.160 73.650 ;
        RECT 30.340 73.570 30.590 75.730 ;
        RECT 31.200 76.080 32.500 76.480 ;
        RECT 32.730 76.930 33.680 76.960 ;
        RECT 32.730 76.760 32.760 76.930 ;
        RECT 32.930 76.760 33.120 76.930 ;
        RECT 33.290 76.760 33.480 76.930 ;
        RECT 33.650 76.760 33.680 76.930 ;
        RECT 34.290 76.930 35.240 76.960 ;
        RECT 31.200 75.300 31.530 76.080 ;
        RECT 32.730 76.000 33.680 76.760 ;
      LAYER li1 ;
        RECT 33.860 76.120 34.110 76.830 ;
      LAYER li1 ;
        RECT 34.290 76.760 34.320 76.930 ;
        RECT 34.490 76.760 34.680 76.930 ;
        RECT 34.850 76.760 35.040 76.930 ;
        RECT 35.210 76.760 35.240 76.930 ;
        RECT 35.850 76.930 36.800 76.960 ;
        RECT 34.290 76.300 35.240 76.760 ;
      LAYER li1 ;
        RECT 35.420 76.120 35.670 76.830 ;
        RECT 33.860 75.950 35.670 76.120 ;
      LAYER li1 ;
        RECT 35.850 76.760 35.880 76.930 ;
        RECT 36.050 76.760 36.240 76.930 ;
        RECT 36.410 76.760 36.600 76.930 ;
        RECT 36.770 76.760 36.800 76.930 ;
        RECT 37.610 76.930 39.220 76.960 ;
        RECT 35.850 76.080 36.800 76.760 ;
      LAYER li1 ;
        RECT 33.860 75.780 34.030 75.950 ;
      LAYER li1 ;
        RECT 36.980 75.900 37.310 76.830 ;
        RECT 37.610 76.760 37.660 76.930 ;
        RECT 37.830 76.760 38.100 76.930 ;
        RECT 38.270 76.760 38.540 76.930 ;
        RECT 38.710 76.760 38.950 76.930 ;
        RECT 39.120 76.760 39.220 76.930 ;
        RECT 37.610 76.480 39.220 76.760 ;
        RECT 31.740 74.640 32.070 75.630 ;
      LAYER li1 ;
        RECT 32.770 75.550 34.030 75.780 ;
      LAYER li1 ;
        RECT 36.070 75.770 37.310 75.900 ;
        RECT 34.210 75.730 37.310 75.770 ;
        RECT 34.210 75.600 36.240 75.730 ;
      LAYER li1 ;
        RECT 33.860 75.420 34.030 75.550 ;
        RECT 33.860 75.250 35.750 75.420 ;
      LAYER li1 ;
        RECT 30.970 73.770 32.420 74.640 ;
        RECT 30.970 73.600 31.220 73.770 ;
        RECT 31.390 73.600 31.580 73.770 ;
        RECT 31.750 73.600 32.020 73.770 ;
        RECT 32.190 73.600 32.420 73.770 ;
        RECT 30.970 73.570 32.420 73.600 ;
        RECT 32.730 73.820 33.680 75.150 ;
        RECT 32.730 73.650 32.760 73.820 ;
        RECT 32.930 73.650 33.120 73.820 ;
        RECT 33.290 73.650 33.480 73.820 ;
        RECT 33.650 73.650 33.680 73.820 ;
        RECT 32.730 73.570 33.680 73.650 ;
      LAYER li1 ;
        RECT 33.860 73.570 34.110 75.250 ;
      LAYER li1 ;
        RECT 34.290 73.820 35.240 75.070 ;
        RECT 34.290 73.650 34.320 73.820 ;
        RECT 34.490 73.650 34.680 73.820 ;
        RECT 34.850 73.650 35.040 73.820 ;
        RECT 35.210 73.650 35.240 73.820 ;
        RECT 34.290 73.570 35.240 73.650 ;
      LAYER li1 ;
        RECT 35.420 73.570 35.750 75.250 ;
        RECT 36.530 75.210 36.860 75.550 ;
      LAYER li1 ;
        RECT 35.930 73.820 36.880 75.030 ;
        RECT 35.930 73.650 35.960 73.820 ;
        RECT 36.130 73.650 36.320 73.820 ;
        RECT 36.490 73.650 36.680 73.820 ;
        RECT 36.850 73.650 36.880 73.820 ;
        RECT 35.930 73.570 36.880 73.650 ;
        RECT 37.060 73.570 37.310 75.730 ;
        RECT 37.920 76.080 39.220 76.480 ;
        RECT 39.450 76.930 40.400 76.960 ;
        RECT 39.450 76.760 39.480 76.930 ;
        RECT 39.650 76.760 39.840 76.930 ;
        RECT 40.010 76.760 40.200 76.930 ;
        RECT 40.370 76.760 40.400 76.930 ;
        RECT 41.010 76.930 41.960 76.960 ;
        RECT 37.920 75.300 38.250 76.080 ;
        RECT 39.450 76.000 40.400 76.760 ;
      LAYER li1 ;
        RECT 40.580 76.120 40.830 76.830 ;
      LAYER li1 ;
        RECT 41.010 76.760 41.040 76.930 ;
        RECT 41.210 76.760 41.400 76.930 ;
        RECT 41.570 76.760 41.760 76.930 ;
        RECT 41.930 76.760 41.960 76.930 ;
        RECT 42.570 76.930 43.520 76.960 ;
        RECT 41.010 76.300 41.960 76.760 ;
      LAYER li1 ;
        RECT 42.140 76.120 42.390 76.830 ;
        RECT 40.580 75.950 42.390 76.120 ;
      LAYER li1 ;
        RECT 42.570 76.760 42.600 76.930 ;
        RECT 42.770 76.760 42.960 76.930 ;
        RECT 43.130 76.760 43.320 76.930 ;
        RECT 43.490 76.760 43.520 76.930 ;
        RECT 44.330 76.930 45.940 76.960 ;
        RECT 42.570 76.080 43.520 76.760 ;
      LAYER li1 ;
        RECT 40.580 75.780 40.750 75.950 ;
      LAYER li1 ;
        RECT 43.700 75.900 44.030 76.830 ;
        RECT 44.330 76.760 44.380 76.930 ;
        RECT 44.550 76.760 44.820 76.930 ;
        RECT 44.990 76.760 45.260 76.930 ;
        RECT 45.430 76.760 45.670 76.930 ;
        RECT 45.840 76.760 45.940 76.930 ;
        RECT 44.330 76.480 45.940 76.760 ;
        RECT 38.460 74.640 38.790 75.630 ;
      LAYER li1 ;
        RECT 39.490 75.550 40.750 75.780 ;
      LAYER li1 ;
        RECT 42.790 75.770 44.030 75.900 ;
        RECT 40.930 75.730 44.030 75.770 ;
        RECT 40.930 75.600 42.960 75.730 ;
      LAYER li1 ;
        RECT 40.580 75.420 40.750 75.550 ;
        RECT 40.580 75.250 42.470 75.420 ;
      LAYER li1 ;
        RECT 37.690 73.770 39.140 74.640 ;
        RECT 37.690 73.600 37.940 73.770 ;
        RECT 38.110 73.600 38.300 73.770 ;
        RECT 38.470 73.600 38.740 73.770 ;
        RECT 38.910 73.600 39.140 73.770 ;
        RECT 37.690 73.570 39.140 73.600 ;
        RECT 39.450 73.820 40.400 75.150 ;
        RECT 39.450 73.650 39.480 73.820 ;
        RECT 39.650 73.650 39.840 73.820 ;
        RECT 40.010 73.650 40.200 73.820 ;
        RECT 40.370 73.650 40.400 73.820 ;
        RECT 39.450 73.570 40.400 73.650 ;
      LAYER li1 ;
        RECT 40.580 73.570 40.830 75.250 ;
      LAYER li1 ;
        RECT 41.010 73.820 41.960 75.070 ;
        RECT 41.010 73.650 41.040 73.820 ;
        RECT 41.210 73.650 41.400 73.820 ;
        RECT 41.570 73.650 41.760 73.820 ;
        RECT 41.930 73.650 41.960 73.820 ;
        RECT 41.010 73.570 41.960 73.650 ;
      LAYER li1 ;
        RECT 42.140 73.570 42.470 75.250 ;
        RECT 43.250 75.210 43.580 75.550 ;
      LAYER li1 ;
        RECT 42.650 73.820 43.600 75.030 ;
        RECT 42.650 73.650 42.680 73.820 ;
        RECT 42.850 73.650 43.040 73.820 ;
        RECT 43.210 73.650 43.400 73.820 ;
        RECT 43.570 73.650 43.600 73.820 ;
        RECT 42.650 73.570 43.600 73.650 ;
        RECT 43.780 73.570 44.030 75.730 ;
        RECT 44.640 76.080 45.940 76.480 ;
        RECT 47.610 76.930 48.560 76.960 ;
        RECT 47.610 76.760 47.640 76.930 ;
        RECT 47.810 76.760 48.000 76.930 ;
        RECT 48.170 76.760 48.360 76.930 ;
        RECT 48.530 76.760 48.560 76.930 ;
        RECT 49.170 76.930 50.120 76.960 ;
        RECT 44.640 75.300 44.970 76.080 ;
        RECT 47.610 76.000 48.560 76.760 ;
      LAYER li1 ;
        RECT 48.740 76.120 48.990 76.830 ;
      LAYER li1 ;
        RECT 49.170 76.760 49.200 76.930 ;
        RECT 49.370 76.760 49.560 76.930 ;
        RECT 49.730 76.760 49.920 76.930 ;
        RECT 50.090 76.760 50.120 76.930 ;
        RECT 50.730 76.930 51.680 76.960 ;
        RECT 49.170 76.300 50.120 76.760 ;
      LAYER li1 ;
        RECT 50.300 76.120 50.550 76.830 ;
        RECT 48.740 75.950 50.550 76.120 ;
      LAYER li1 ;
        RECT 50.730 76.760 50.760 76.930 ;
        RECT 50.930 76.760 51.120 76.930 ;
        RECT 51.290 76.760 51.480 76.930 ;
        RECT 51.650 76.760 51.680 76.930 ;
        RECT 52.490 76.930 54.100 76.960 ;
        RECT 54.840 76.930 56.450 76.960 ;
        RECT 57.300 76.930 58.960 76.960 ;
        RECT 50.730 76.080 51.680 76.760 ;
      LAYER li1 ;
        RECT 48.740 75.780 48.910 75.950 ;
      LAYER li1 ;
        RECT 51.860 75.900 52.190 76.830 ;
        RECT 52.490 76.760 52.540 76.930 ;
        RECT 52.710 76.760 52.980 76.930 ;
        RECT 53.150 76.760 53.420 76.930 ;
        RECT 53.590 76.760 53.830 76.930 ;
        RECT 54.000 76.760 54.100 76.930 ;
        RECT 52.490 76.480 54.100 76.760 ;
        RECT 45.180 74.640 45.510 75.630 ;
      LAYER li1 ;
        RECT 47.650 75.550 48.910 75.780 ;
      LAYER li1 ;
        RECT 50.950 75.770 52.190 75.900 ;
        RECT 49.090 75.730 52.190 75.770 ;
        RECT 49.090 75.600 51.120 75.730 ;
      LAYER li1 ;
        RECT 48.740 75.420 48.910 75.550 ;
        RECT 48.740 75.250 50.630 75.420 ;
      LAYER li1 ;
        RECT 44.410 73.770 45.860 74.640 ;
        RECT 44.410 73.600 44.660 73.770 ;
        RECT 44.830 73.600 45.020 73.770 ;
        RECT 45.190 73.600 45.460 73.770 ;
        RECT 45.630 73.600 45.860 73.770 ;
        RECT 44.410 73.570 45.860 73.600 ;
        RECT 47.610 73.820 48.560 75.150 ;
        RECT 47.610 73.650 47.640 73.820 ;
        RECT 47.810 73.650 48.000 73.820 ;
        RECT 48.170 73.650 48.360 73.820 ;
        RECT 48.530 73.650 48.560 73.820 ;
        RECT 47.610 73.570 48.560 73.650 ;
      LAYER li1 ;
        RECT 48.740 73.570 48.990 75.250 ;
      LAYER li1 ;
        RECT 49.170 73.820 50.120 75.070 ;
        RECT 49.170 73.650 49.200 73.820 ;
        RECT 49.370 73.650 49.560 73.820 ;
        RECT 49.730 73.650 49.920 73.820 ;
        RECT 50.090 73.650 50.120 73.820 ;
        RECT 49.170 73.570 50.120 73.650 ;
      LAYER li1 ;
        RECT 50.300 73.570 50.630 75.250 ;
        RECT 51.410 75.210 51.740 75.550 ;
      LAYER li1 ;
        RECT 50.810 73.820 51.760 75.030 ;
        RECT 50.810 73.650 50.840 73.820 ;
        RECT 51.010 73.650 51.200 73.820 ;
        RECT 51.370 73.650 51.560 73.820 ;
        RECT 51.730 73.650 51.760 73.820 ;
        RECT 50.810 73.570 51.760 73.650 ;
        RECT 51.940 73.570 52.190 75.730 ;
        RECT 52.800 76.080 54.100 76.480 ;
        RECT 52.800 75.300 53.130 76.080 ;
        RECT 53.340 74.640 53.670 75.630 ;
      LAYER li1 ;
        RECT 54.370 75.400 54.660 76.830 ;
      LAYER li1 ;
        RECT 55.010 76.760 55.200 76.930 ;
        RECT 55.370 76.760 55.560 76.930 ;
        RECT 55.730 76.760 55.920 76.930 ;
        RECT 56.090 76.760 56.280 76.930 ;
        RECT 54.840 76.150 56.450 76.760 ;
        RECT 56.630 76.410 57.120 76.830 ;
        RECT 57.300 76.760 57.330 76.930 ;
        RECT 57.500 76.760 57.690 76.930 ;
        RECT 57.860 76.760 58.050 76.930 ;
        RECT 58.220 76.760 58.410 76.930 ;
        RECT 58.580 76.760 58.770 76.930 ;
        RECT 58.940 76.760 58.960 76.930 ;
        RECT 59.690 76.930 61.300 76.960 ;
        RECT 57.300 76.410 58.960 76.760 ;
        RECT 56.630 75.970 56.800 76.410 ;
        RECT 54.860 75.800 56.800 75.970 ;
      LAYER li1 ;
        RECT 56.980 75.940 57.930 76.230 ;
      LAYER li1 ;
        RECT 59.140 76.220 59.390 76.830 ;
        RECT 59.690 76.760 59.740 76.930 ;
        RECT 59.910 76.760 60.180 76.930 ;
        RECT 60.350 76.760 60.620 76.930 ;
        RECT 60.790 76.760 61.030 76.930 ;
        RECT 61.200 76.760 61.300 76.930 ;
        RECT 62.000 76.930 62.950 76.960 ;
        RECT 59.690 76.480 61.300 76.760 ;
        RECT 58.110 76.050 59.390 76.220 ;
        RECT 54.860 75.580 55.190 75.800 ;
        RECT 52.570 73.770 54.020 74.640 ;
        RECT 52.570 73.600 52.820 73.770 ;
        RECT 52.990 73.600 53.180 73.770 ;
        RECT 53.350 73.600 53.620 73.770 ;
        RECT 53.790 73.600 54.020 73.770 ;
        RECT 52.570 73.570 54.020 73.600 ;
      LAYER li1 ;
        RECT 54.370 73.570 54.740 75.400 ;
      LAYER li1 ;
        RECT 54.920 73.820 55.500 75.150 ;
      LAYER li1 ;
        RECT 55.680 74.230 56.010 75.620 ;
      LAYER li1 ;
        RECT 56.190 74.910 56.360 75.800 ;
      LAYER li1 ;
        RECT 56.980 75.540 57.150 75.940 ;
        RECT 56.540 75.370 57.150 75.540 ;
        RECT 57.330 75.370 57.930 75.760 ;
      LAYER li1 ;
        RECT 58.110 75.550 58.360 76.050 ;
      LAYER li1 ;
        RECT 56.540 75.090 56.870 75.370 ;
        RECT 58.610 75.190 58.920 75.780 ;
        RECT 57.300 75.020 58.920 75.190 ;
      LAYER li1 ;
        RECT 56.190 74.740 57.120 74.910 ;
        RECT 56.790 74.410 57.120 74.740 ;
      LAYER li1 ;
        RECT 57.300 74.230 57.470 75.020 ;
        RECT 55.680 74.060 57.470 74.230 ;
      LAYER li1 ;
        RECT 54.920 73.650 54.940 73.820 ;
        RECT 55.110 73.650 55.300 73.820 ;
        RECT 55.470 73.650 55.500 73.820 ;
        RECT 54.920 73.570 55.500 73.650 ;
        RECT 57.650 73.820 58.960 74.830 ;
        RECT 59.140 74.410 59.390 76.050 ;
        RECT 60.000 76.080 61.300 76.480 ;
        RECT 60.000 75.300 60.330 76.080 ;
        RECT 60.540 74.640 60.870 75.630 ;
        RECT 61.550 74.970 61.820 76.830 ;
        RECT 62.000 76.760 62.030 76.930 ;
        RECT 62.200 76.760 62.390 76.930 ;
        RECT 62.560 76.760 62.750 76.930 ;
        RECT 62.920 76.760 62.950 76.930 ;
        RECT 63.640 76.930 64.230 76.960 ;
        RECT 62.000 76.330 62.950 76.760 ;
        RECT 63.130 76.330 63.460 76.830 ;
        RECT 62.680 74.970 63.010 75.470 ;
        RECT 61.550 74.800 63.010 74.970 ;
        RECT 57.650 73.650 57.680 73.820 ;
        RECT 57.850 73.650 58.040 73.820 ;
        RECT 58.210 73.650 58.400 73.820 ;
        RECT 58.570 73.650 58.760 73.820 ;
        RECT 58.930 73.650 58.960 73.820 ;
        RECT 57.650 73.620 58.960 73.650 ;
        RECT 59.770 73.770 61.220 74.640 ;
        RECT 61.550 73.870 61.880 74.800 ;
        RECT 59.770 73.600 60.020 73.770 ;
        RECT 60.190 73.600 60.380 73.770 ;
        RECT 60.550 73.600 60.820 73.770 ;
        RECT 60.990 73.600 61.220 73.770 ;
        RECT 62.070 73.820 62.660 74.600 ;
        RECT 62.070 73.650 62.100 73.820 ;
        RECT 62.270 73.650 62.460 73.820 ;
        RECT 62.630 73.650 62.660 73.820 ;
        RECT 62.070 73.620 62.660 73.650 ;
        RECT 62.840 73.690 63.010 74.800 ;
        RECT 63.190 75.410 63.460 76.330 ;
        RECT 63.640 76.760 63.670 76.930 ;
        RECT 63.840 76.760 64.030 76.930 ;
        RECT 64.200 76.760 64.230 76.930 ;
        RECT 68.600 76.930 69.550 76.960 ;
        RECT 63.640 76.080 64.230 76.760 ;
      LAYER li1 ;
        RECT 64.510 76.700 67.450 76.870 ;
        RECT 64.510 75.710 64.680 76.700 ;
      LAYER li1 ;
        RECT 63.190 75.180 63.720 75.410 ;
        RECT 63.190 73.870 63.440 75.180 ;
      LAYER li1 ;
        RECT 64.140 74.840 64.680 75.710 ;
        RECT 64.860 75.220 65.190 76.520 ;
      LAYER li1 ;
        RECT 65.370 76.000 65.640 76.500 ;
        RECT 66.090 76.250 66.420 76.500 ;
        RECT 66.090 76.080 67.100 76.250 ;
        RECT 65.370 75.010 65.540 76.000 ;
        RECT 66.420 75.410 66.750 75.900 ;
        RECT 65.320 74.840 65.540 75.010 ;
        RECT 65.720 75.180 66.750 75.410 ;
        RECT 66.930 75.850 67.100 76.080 ;
      LAYER li1 ;
        RECT 67.280 76.200 67.450 76.700 ;
      LAYER li1 ;
        RECT 68.600 76.760 68.630 76.930 ;
        RECT 68.800 76.760 68.990 76.930 ;
        RECT 69.160 76.760 69.350 76.930 ;
        RECT 69.520 76.760 69.550 76.930 ;
        RECT 68.600 76.380 69.550 76.760 ;
      LAYER li1 ;
        RECT 69.730 76.890 72.390 77.060 ;
        RECT 69.730 76.200 69.900 76.890 ;
        RECT 67.280 76.030 69.900 76.200 ;
      LAYER li1 ;
        RECT 66.930 75.680 69.550 75.850 ;
        RECT 65.320 74.660 65.490 74.840 ;
        RECT 65.720 74.660 65.890 75.180 ;
        RECT 66.930 75.000 67.100 75.680 ;
      LAYER li1 ;
        RECT 69.730 75.500 69.900 76.030 ;
      LAYER li1 ;
        RECT 63.680 74.490 65.490 74.660 ;
        RECT 63.680 73.870 63.930 74.490 ;
        RECT 64.110 74.140 65.140 74.310 ;
        RECT 64.110 73.690 64.280 74.140 ;
        RECT 59.770 73.570 61.220 73.600 ;
        RECT 62.840 73.520 64.280 73.690 ;
        RECT 64.460 73.820 64.790 73.960 ;
        RECT 64.460 73.650 64.490 73.820 ;
        RECT 64.660 73.650 64.790 73.820 ;
        RECT 64.460 73.620 64.790 73.650 ;
        RECT 64.970 73.690 65.140 74.140 ;
        RECT 65.320 73.870 65.490 74.490 ;
        RECT 65.670 74.330 65.890 74.660 ;
        RECT 66.070 74.830 67.100 75.000 ;
        RECT 67.280 75.150 67.610 75.500 ;
      LAYER li1 ;
        RECT 68.050 75.330 69.900 75.500 ;
      LAYER li1 ;
        RECT 70.080 76.000 70.410 76.710 ;
        RECT 70.870 76.540 72.040 76.710 ;
        RECT 70.870 76.000 71.200 76.540 ;
        RECT 70.080 75.150 70.340 76.000 ;
        RECT 71.410 75.740 71.690 76.240 ;
        RECT 67.280 74.980 70.340 75.150 ;
        RECT 66.070 74.130 66.240 74.830 ;
        RECT 66.930 74.800 67.100 74.830 ;
        RECT 66.420 74.450 66.750 74.650 ;
        RECT 66.930 74.630 68.700 74.800 ;
        RECT 66.420 74.330 68.190 74.450 ;
        RECT 66.540 74.280 68.190 74.330 ;
        RECT 66.020 73.870 66.350 74.130 ;
        RECT 66.540 73.690 66.710 74.280 ;
        RECT 64.970 73.520 66.710 73.690 ;
        RECT 66.890 73.820 67.840 74.100 ;
        RECT 66.890 73.650 66.920 73.820 ;
        RECT 67.090 73.650 67.280 73.820 ;
        RECT 67.450 73.650 67.640 73.820 ;
        RECT 67.810 73.650 67.840 73.820 ;
        RECT 66.890 73.620 67.840 73.650 ;
        RECT 68.020 73.690 68.190 74.280 ;
        RECT 68.370 73.870 68.700 74.630 ;
        RECT 70.010 74.400 70.340 74.980 ;
        RECT 70.520 75.570 71.690 75.740 ;
        RECT 70.520 74.220 70.690 75.570 ;
        RECT 71.070 74.890 71.400 75.390 ;
        RECT 71.870 75.140 72.040 76.540 ;
      LAYER li1 ;
        RECT 72.220 76.230 72.390 76.890 ;
      LAYER li1 ;
        RECT 72.570 76.930 73.520 76.960 ;
        RECT 72.570 76.760 72.600 76.930 ;
        RECT 72.770 76.760 72.960 76.930 ;
        RECT 73.130 76.760 73.320 76.930 ;
        RECT 73.490 76.760 73.520 76.930 ;
        RECT 75.180 76.930 76.130 76.960 ;
        RECT 72.570 76.410 73.520 76.760 ;
        RECT 74.060 76.330 74.390 76.830 ;
        RECT 75.180 76.760 75.210 76.930 ;
        RECT 75.380 76.760 75.570 76.930 ;
        RECT 75.740 76.760 75.930 76.930 ;
        RECT 76.100 76.760 76.130 76.930 ;
      LAYER li1 ;
        RECT 72.220 76.120 73.230 76.230 ;
        RECT 72.220 76.060 73.280 76.120 ;
        RECT 72.900 75.950 73.280 76.060 ;
      LAYER li1 ;
        RECT 72.250 75.490 72.580 75.880 ;
      LAYER li1 ;
        RECT 72.900 75.670 73.230 75.950 ;
      LAYER li1 ;
        RECT 74.060 75.490 74.290 76.330 ;
        RECT 74.670 75.830 75.000 76.330 ;
        RECT 75.180 75.830 76.130 76.760 ;
        RECT 76.970 76.930 78.580 76.960 ;
        RECT 76.970 76.760 77.020 76.930 ;
        RECT 77.190 76.760 77.460 76.930 ;
        RECT 77.630 76.760 77.900 76.930 ;
        RECT 78.070 76.760 78.310 76.930 ;
        RECT 78.480 76.760 78.580 76.930 ;
        RECT 76.970 76.480 78.580 76.760 ;
        RECT 77.280 76.080 78.580 76.480 ;
        RECT 79.290 76.930 79.880 76.960 ;
        RECT 79.290 76.760 79.320 76.930 ;
        RECT 79.490 76.760 79.680 76.930 ;
        RECT 79.850 76.760 79.880 76.930 ;
        RECT 80.810 76.930 82.420 76.960 ;
        RECT 83.120 76.930 84.010 76.960 ;
        RECT 72.250 75.320 74.290 75.490 ;
        RECT 71.580 74.970 73.940 75.140 ;
        RECT 71.580 74.650 71.750 74.970 ;
        RECT 74.120 74.790 74.290 75.320 ;
        RECT 68.880 74.050 70.690 74.220 ;
        RECT 70.870 74.480 71.750 74.650 ;
        RECT 68.880 73.690 69.050 74.050 ;
        RECT 68.020 73.520 69.050 73.690 ;
        RECT 69.230 73.820 70.180 73.870 ;
        RECT 69.230 73.650 69.260 73.820 ;
        RECT 69.430 73.650 69.620 73.820 ;
        RECT 69.790 73.650 69.980 73.820 ;
        RECT 70.150 73.650 70.180 73.820 ;
        RECT 69.230 73.570 70.180 73.650 ;
        RECT 70.870 73.570 71.120 74.480 ;
        RECT 71.930 73.820 72.880 74.650 ;
        RECT 73.280 74.620 74.290 74.790 ;
        RECT 74.790 75.650 75.000 75.830 ;
        RECT 74.790 75.320 76.160 75.650 ;
        RECT 73.280 74.150 73.530 74.620 ;
        RECT 73.710 73.820 74.610 74.440 ;
        RECT 74.790 74.320 75.040 75.320 ;
        RECT 77.280 75.300 77.610 76.080 ;
        RECT 79.290 76.000 79.880 76.760 ;
        RECT 71.930 73.650 71.960 73.820 ;
        RECT 72.130 73.650 72.320 73.820 ;
        RECT 72.490 73.650 72.680 73.820 ;
        RECT 72.850 73.650 72.880 73.820 ;
        RECT 73.880 73.650 74.070 73.820 ;
        RECT 74.240 73.650 74.430 73.820 ;
        RECT 74.600 73.650 74.610 73.820 ;
        RECT 71.930 73.620 72.880 73.650 ;
        RECT 73.710 73.620 74.610 73.650 ;
        RECT 75.220 73.820 76.160 75.130 ;
        RECT 77.820 74.640 78.150 75.630 ;
      LAYER li1 ;
        RECT 79.330 75.390 80.040 75.780 ;
        RECT 80.220 75.150 80.550 76.830 ;
      LAYER li1 ;
        RECT 80.810 76.760 80.860 76.930 ;
        RECT 81.030 76.760 81.300 76.930 ;
        RECT 81.470 76.760 81.740 76.930 ;
        RECT 81.910 76.760 82.150 76.930 ;
        RECT 82.320 76.760 82.420 76.930 ;
        RECT 80.810 76.480 82.420 76.760 ;
        RECT 81.120 76.080 82.420 76.480 ;
        RECT 81.120 75.300 81.450 76.080 ;
        RECT 75.220 73.650 75.240 73.820 ;
        RECT 75.410 73.650 75.600 73.820 ;
        RECT 75.770 73.650 75.960 73.820 ;
        RECT 76.130 73.650 76.160 73.820 ;
        RECT 75.220 73.590 76.160 73.650 ;
        RECT 77.050 73.770 78.500 74.640 ;
        RECT 77.050 73.600 77.300 73.770 ;
        RECT 77.470 73.600 77.660 73.770 ;
        RECT 77.830 73.600 78.100 73.770 ;
        RECT 78.270 73.600 78.500 73.770 ;
        RECT 77.050 73.570 78.500 73.600 ;
        RECT 79.290 73.820 79.880 75.150 ;
        RECT 79.290 73.650 79.320 73.820 ;
        RECT 79.490 73.650 79.680 73.820 ;
        RECT 79.850 73.650 79.880 73.820 ;
        RECT 79.290 73.570 79.880 73.650 ;
      LAYER li1 ;
        RECT 80.160 73.570 80.550 75.150 ;
      LAYER li1 ;
        RECT 81.660 74.640 81.990 75.630 ;
        RECT 80.890 73.770 82.340 74.640 ;
        RECT 80.890 73.600 81.140 73.770 ;
        RECT 81.310 73.600 81.500 73.770 ;
        RECT 81.670 73.600 81.940 73.770 ;
        RECT 82.110 73.600 82.340 73.770 ;
        RECT 80.890 73.570 82.340 73.600 ;
      LAYER li1 ;
        RECT 82.690 73.570 82.940 76.830 ;
      LAYER li1 ;
        RECT 83.290 76.760 83.480 76.930 ;
        RECT 83.650 76.760 83.840 76.930 ;
        RECT 84.310 76.890 86.240 77.060 ;
        RECT 83.120 76.080 84.010 76.760 ;
        RECT 84.310 76.460 84.640 76.890 ;
        RECT 85.090 76.450 85.420 76.710 ;
        RECT 84.820 76.280 85.420 76.450 ;
        RECT 85.910 76.300 86.240 76.890 ;
        RECT 86.450 76.930 87.750 76.960 ;
        RECT 86.450 76.760 86.480 76.930 ;
        RECT 86.650 76.760 86.840 76.930 ;
        RECT 87.010 76.760 87.200 76.930 ;
        RECT 87.370 76.760 87.560 76.930 ;
        RECT 87.730 76.760 87.750 76.930 ;
        RECT 86.450 76.280 87.750 76.760 ;
        RECT 88.010 76.930 89.620 76.960 ;
        RECT 88.010 76.760 88.060 76.930 ;
        RECT 88.230 76.760 88.500 76.930 ;
        RECT 88.670 76.760 88.940 76.930 ;
        RECT 89.110 76.760 89.350 76.930 ;
        RECT 89.520 76.760 89.620 76.930 ;
        RECT 90.310 76.930 91.080 76.960 ;
        RECT 92.550 76.930 93.440 76.960 ;
        RECT 94.250 76.930 95.860 76.960 ;
        RECT 96.640 76.930 97.530 76.960 ;
        RECT 99.530 76.930 101.140 76.960 ;
        RECT 101.880 76.930 103.490 76.960 ;
        RECT 104.340 76.930 106.000 76.960 ;
        RECT 88.010 76.480 89.620 76.760 ;
        RECT 84.190 76.110 84.990 76.280 ;
        RECT 84.190 75.900 84.360 76.110 ;
      LAYER li1 ;
        RECT 85.600 76.100 86.270 76.120 ;
        RECT 85.170 75.930 87.440 76.100 ;
      LAYER li1 ;
        RECT 83.150 75.730 84.360 75.900 ;
      LAYER li1 ;
        RECT 84.540 75.760 85.340 75.930 ;
      LAYER li1 ;
        RECT 83.150 75.030 83.480 75.730 ;
      LAYER li1 ;
        RECT 84.540 75.550 84.710 75.760 ;
        RECT 87.110 75.750 87.440 75.930 ;
        RECT 83.980 75.270 84.710 75.550 ;
        RECT 84.890 75.210 85.320 75.580 ;
        RECT 85.520 75.210 85.810 75.750 ;
        RECT 86.050 75.420 86.760 75.750 ;
        RECT 87.030 75.580 87.440 75.750 ;
        RECT 87.110 75.310 87.440 75.580 ;
      LAYER li1 ;
        RECT 88.320 76.080 89.620 76.480 ;
        RECT 88.320 75.300 88.650 76.080 ;
        RECT 85.990 75.030 86.240 75.150 ;
        RECT 83.150 74.860 86.240 75.030 ;
        RECT 83.120 73.820 85.810 74.680 ;
        RECT 83.290 73.650 83.480 73.820 ;
        RECT 83.650 73.650 83.840 73.820 ;
        RECT 84.010 73.650 84.200 73.820 ;
        RECT 84.370 73.650 84.560 73.820 ;
        RECT 84.730 73.650 84.920 73.820 ;
        RECT 85.090 73.650 85.280 73.820 ;
        RECT 85.450 73.650 85.640 73.820 ;
        RECT 83.120 73.570 85.810 73.650 ;
        RECT 85.990 73.570 86.240 74.860 ;
        RECT 86.420 73.820 87.730 75.130 ;
        RECT 88.860 74.640 89.190 75.630 ;
      LAYER li1 ;
        RECT 89.890 75.350 90.140 76.800 ;
      LAYER li1 ;
        RECT 90.310 76.760 90.360 76.930 ;
        RECT 90.530 76.760 90.870 76.930 ;
        RECT 91.040 76.760 91.080 76.930 ;
        RECT 90.310 76.050 91.080 76.760 ;
        RECT 91.260 75.870 91.590 76.830 ;
        RECT 92.040 76.220 92.370 76.830 ;
        RECT 92.720 76.760 92.910 76.930 ;
        RECT 93.080 76.760 93.270 76.930 ;
        RECT 92.550 76.400 93.440 76.760 ;
        RECT 93.620 76.220 93.950 76.830 ;
        RECT 94.250 76.760 94.300 76.930 ;
        RECT 94.470 76.760 94.740 76.930 ;
        RECT 94.910 76.760 95.180 76.930 ;
        RECT 95.350 76.760 95.590 76.930 ;
        RECT 95.760 76.760 95.860 76.930 ;
        RECT 94.250 76.480 95.860 76.760 ;
        RECT 92.040 76.050 93.950 76.220 ;
        RECT 93.620 76.000 93.950 76.050 ;
        RECT 94.560 76.080 95.860 76.480 ;
        RECT 96.130 76.220 96.460 76.830 ;
        RECT 96.810 76.760 97.000 76.930 ;
        RECT 97.170 76.760 97.360 76.930 ;
        RECT 96.640 76.400 97.530 76.760 ;
        RECT 97.710 76.220 98.040 76.830 ;
        RECT 90.310 75.700 92.140 75.870 ;
        RECT 90.310 75.530 90.600 75.700 ;
        RECT 86.420 73.650 86.450 73.820 ;
        RECT 86.620 73.650 86.810 73.820 ;
        RECT 86.980 73.650 87.170 73.820 ;
        RECT 87.340 73.650 87.530 73.820 ;
        RECT 87.700 73.650 87.730 73.820 ;
        RECT 86.420 73.590 87.730 73.650 ;
        RECT 88.090 73.770 89.540 74.640 ;
        RECT 88.090 73.600 88.340 73.770 ;
        RECT 88.510 73.600 88.700 73.770 ;
        RECT 88.870 73.600 89.140 73.770 ;
        RECT 89.310 73.600 89.540 73.770 ;
        RECT 88.090 73.570 89.540 73.600 ;
      LAYER li1 ;
        RECT 89.890 73.570 90.360 75.350 ;
        RECT 90.850 75.210 91.760 75.520 ;
      LAYER li1 ;
        RECT 90.540 73.820 91.790 75.030 ;
        RECT 90.710 73.650 90.900 73.820 ;
        RECT 91.070 73.650 91.260 73.820 ;
        RECT 91.430 73.650 91.620 73.820 ;
        RECT 90.540 73.570 91.790 73.650 ;
        RECT 91.970 73.570 92.140 75.700 ;
      LAYER li1 ;
        RECT 92.320 75.010 92.550 75.780 ;
        RECT 92.770 75.490 93.960 75.820 ;
      LAYER li1 ;
        RECT 94.560 75.300 94.890 76.080 ;
        RECT 96.130 76.050 98.040 76.220 ;
        RECT 96.130 76.000 96.460 76.050 ;
      LAYER li1 ;
        RECT 98.490 75.870 98.820 76.830 ;
      LAYER li1 ;
        RECT 99.530 76.760 99.580 76.930 ;
        RECT 99.750 76.760 100.020 76.930 ;
        RECT 100.190 76.760 100.460 76.930 ;
        RECT 100.630 76.760 100.870 76.930 ;
        RECT 101.040 76.760 101.140 76.930 ;
        RECT 99.530 76.480 101.140 76.760 ;
      LAYER li1 ;
        RECT 92.310 74.840 92.550 75.010 ;
        RECT 92.320 74.070 92.550 74.840 ;
      LAYER li1 ;
        RECT 92.730 73.820 93.990 75.150 ;
        RECT 95.100 74.640 95.430 75.630 ;
      LAYER li1 ;
        RECT 97.070 75.570 97.800 75.820 ;
        RECT 97.980 75.700 98.820 75.870 ;
      LAYER li1 ;
        RECT 99.840 76.080 101.140 76.480 ;
      LAYER li1 ;
        RECT 97.980 75.390 98.150 75.700 ;
        RECT 97.570 75.220 98.150 75.390 ;
      LAYER li1 ;
        RECT 92.900 73.650 93.090 73.820 ;
        RECT 93.260 73.650 93.450 73.820 ;
        RECT 93.620 73.650 93.810 73.820 ;
        RECT 93.980 73.650 93.990 73.820 ;
        RECT 92.730 73.570 93.990 73.650 ;
        RECT 94.330 73.770 95.780 74.640 ;
        RECT 94.330 73.600 94.580 73.770 ;
        RECT 94.750 73.600 94.940 73.770 ;
        RECT 95.110 73.600 95.380 73.770 ;
        RECT 95.550 73.600 95.780 73.770 ;
        RECT 94.330 73.570 95.780 73.600 ;
        RECT 96.090 73.820 97.040 75.150 ;
        RECT 96.090 73.650 96.120 73.820 ;
        RECT 96.290 73.650 96.480 73.820 ;
        RECT 96.650 73.650 96.840 73.820 ;
        RECT 97.010 73.650 97.040 73.820 ;
        RECT 96.090 73.570 97.040 73.650 ;
      LAYER li1 ;
        RECT 97.570 73.570 98.040 75.220 ;
        RECT 98.330 75.210 99.240 75.520 ;
      LAYER li1 ;
        RECT 99.840 75.300 100.170 76.080 ;
        RECT 98.220 73.820 99.170 75.030 ;
        RECT 100.380 74.640 100.710 75.630 ;
      LAYER li1 ;
        RECT 101.410 75.400 101.700 76.830 ;
      LAYER li1 ;
        RECT 102.050 76.760 102.240 76.930 ;
        RECT 102.410 76.760 102.600 76.930 ;
        RECT 102.770 76.760 102.960 76.930 ;
        RECT 103.130 76.760 103.320 76.930 ;
        RECT 101.880 76.150 103.490 76.760 ;
        RECT 103.670 76.410 104.160 76.830 ;
        RECT 104.340 76.760 104.370 76.930 ;
        RECT 104.540 76.760 104.730 76.930 ;
        RECT 104.900 76.760 105.090 76.930 ;
        RECT 105.260 76.760 105.450 76.930 ;
        RECT 105.620 76.760 105.810 76.930 ;
        RECT 105.980 76.760 106.000 76.930 ;
        RECT 106.730 76.930 108.340 76.960 ;
        RECT 104.340 76.410 106.000 76.760 ;
        RECT 103.670 75.970 103.840 76.410 ;
        RECT 101.900 75.800 103.840 75.970 ;
      LAYER li1 ;
        RECT 104.020 75.940 104.970 76.230 ;
      LAYER li1 ;
        RECT 106.180 76.220 106.430 76.830 ;
        RECT 106.730 76.760 106.780 76.930 ;
        RECT 106.950 76.760 107.220 76.930 ;
        RECT 107.390 76.760 107.660 76.930 ;
        RECT 107.830 76.760 108.070 76.930 ;
        RECT 108.240 76.760 108.340 76.930 ;
        RECT 106.730 76.480 108.340 76.760 ;
        RECT 105.150 76.050 106.430 76.220 ;
        RECT 101.900 75.580 102.230 75.800 ;
        RECT 98.220 73.650 98.250 73.820 ;
        RECT 98.420 73.650 98.610 73.820 ;
        RECT 98.780 73.650 98.970 73.820 ;
        RECT 99.140 73.650 99.170 73.820 ;
        RECT 98.220 73.570 99.170 73.650 ;
        RECT 99.610 73.770 101.060 74.640 ;
        RECT 99.610 73.600 99.860 73.770 ;
        RECT 100.030 73.600 100.220 73.770 ;
        RECT 100.390 73.600 100.660 73.770 ;
        RECT 100.830 73.600 101.060 73.770 ;
        RECT 99.610 73.570 101.060 73.600 ;
      LAYER li1 ;
        RECT 101.410 73.570 101.780 75.400 ;
      LAYER li1 ;
        RECT 101.960 73.820 102.540 75.150 ;
      LAYER li1 ;
        RECT 102.720 74.230 103.050 75.620 ;
      LAYER li1 ;
        RECT 103.230 74.910 103.400 75.800 ;
      LAYER li1 ;
        RECT 104.020 75.540 104.190 75.940 ;
      LAYER li1 ;
        RECT 105.150 75.550 105.400 76.050 ;
      LAYER li1 ;
        RECT 103.580 75.370 104.190 75.540 ;
        RECT 103.580 75.090 103.910 75.370 ;
        RECT 105.650 75.190 105.960 75.780 ;
        RECT 104.340 75.020 105.960 75.190 ;
      LAYER li1 ;
        RECT 103.230 74.740 104.160 74.910 ;
        RECT 103.830 74.410 104.160 74.740 ;
      LAYER li1 ;
        RECT 104.340 74.230 104.510 75.020 ;
        RECT 102.720 74.060 104.510 74.230 ;
      LAYER li1 ;
        RECT 101.960 73.650 101.980 73.820 ;
        RECT 102.150 73.650 102.340 73.820 ;
        RECT 102.510 73.650 102.540 73.820 ;
        RECT 101.960 73.570 102.540 73.650 ;
        RECT 104.690 73.820 106.000 74.830 ;
        RECT 106.180 74.410 106.430 76.050 ;
        RECT 107.040 76.080 108.340 76.480 ;
        RECT 109.530 76.930 110.840 76.960 ;
        RECT 109.530 76.760 109.560 76.930 ;
        RECT 109.730 76.760 109.920 76.930 ;
        RECT 110.090 76.760 110.280 76.930 ;
        RECT 110.450 76.760 110.640 76.930 ;
        RECT 110.810 76.760 110.840 76.930 ;
        RECT 112.010 76.930 113.620 76.960 ;
        RECT 107.040 75.300 107.370 76.080 ;
        RECT 109.530 75.980 110.840 76.760 ;
      LAYER li1 ;
        RECT 111.290 76.150 111.620 76.810 ;
      LAYER li1 ;
        RECT 112.010 76.760 112.060 76.930 ;
        RECT 112.230 76.760 112.500 76.930 ;
        RECT 112.670 76.760 112.940 76.930 ;
        RECT 113.110 76.760 113.350 76.930 ;
        RECT 113.520 76.760 113.620 76.930 ;
        RECT 114.320 76.930 115.270 76.960 ;
        RECT 112.010 76.480 113.620 76.760 ;
      LAYER li1 ;
        RECT 111.020 75.980 111.620 76.150 ;
      LAYER li1 ;
        RECT 112.320 76.080 113.620 76.480 ;
      LAYER li1 ;
        RECT 111.020 75.800 111.240 75.980 ;
      LAYER li1 ;
        RECT 107.580 74.640 107.910 75.630 ;
      LAYER li1 ;
        RECT 109.570 75.390 110.460 75.780 ;
        RECT 110.660 75.630 111.240 75.800 ;
      LAYER li1 ;
        RECT 104.690 73.650 104.720 73.820 ;
        RECT 104.890 73.650 105.080 73.820 ;
        RECT 105.250 73.650 105.440 73.820 ;
        RECT 105.610 73.650 105.800 73.820 ;
        RECT 105.970 73.650 106.000 73.820 ;
        RECT 104.690 73.620 106.000 73.650 ;
        RECT 106.810 73.770 108.260 74.640 ;
        RECT 106.810 73.600 107.060 73.770 ;
        RECT 107.230 73.600 107.420 73.770 ;
        RECT 107.590 73.600 107.860 73.770 ;
        RECT 108.030 73.600 108.260 73.770 ;
        RECT 106.810 73.570 108.260 73.600 ;
        RECT 109.530 73.820 110.480 75.150 ;
        RECT 109.530 73.650 109.560 73.820 ;
        RECT 109.730 73.650 109.920 73.820 ;
        RECT 110.090 73.650 110.280 73.820 ;
        RECT 110.450 73.650 110.480 73.820 ;
        RECT 109.530 73.570 110.480 73.650 ;
      LAYER li1 ;
        RECT 110.660 73.570 110.910 75.630 ;
        RECT 111.420 75.470 111.720 75.800 ;
      LAYER li1 ;
        RECT 112.320 75.300 112.650 76.080 ;
        RECT 111.100 73.820 111.690 75.150 ;
        RECT 112.860 74.640 113.190 75.630 ;
      LAYER li1 ;
        RECT 113.430 74.840 113.600 75.750 ;
      LAYER li1 ;
        RECT 113.870 74.970 114.140 76.830 ;
        RECT 114.320 76.760 114.350 76.930 ;
        RECT 114.520 76.760 114.710 76.930 ;
        RECT 114.880 76.760 115.070 76.930 ;
        RECT 115.240 76.760 115.270 76.930 ;
        RECT 115.960 76.930 116.550 76.960 ;
        RECT 114.320 76.330 115.270 76.760 ;
        RECT 115.450 76.330 115.780 76.830 ;
        RECT 115.000 74.970 115.330 75.470 ;
        RECT 113.870 74.800 115.330 74.970 ;
        RECT 111.100 73.650 111.130 73.820 ;
        RECT 111.300 73.650 111.490 73.820 ;
        RECT 111.660 73.650 111.690 73.820 ;
        RECT 111.100 73.570 111.690 73.650 ;
        RECT 112.090 73.770 113.540 74.640 ;
        RECT 113.870 73.870 114.200 74.800 ;
        RECT 112.090 73.600 112.340 73.770 ;
        RECT 112.510 73.600 112.700 73.770 ;
        RECT 112.870 73.600 113.140 73.770 ;
        RECT 113.310 73.600 113.540 73.770 ;
        RECT 114.390 73.820 114.980 74.600 ;
        RECT 114.390 73.650 114.420 73.820 ;
        RECT 114.590 73.650 114.780 73.820 ;
        RECT 114.950 73.650 114.980 73.820 ;
        RECT 114.390 73.620 114.980 73.650 ;
        RECT 115.160 73.690 115.330 74.800 ;
        RECT 115.510 75.410 115.780 76.330 ;
        RECT 115.960 76.760 115.990 76.930 ;
        RECT 116.160 76.760 116.350 76.930 ;
        RECT 116.520 76.760 116.550 76.930 ;
        RECT 120.920 76.930 121.870 76.960 ;
        RECT 115.960 76.080 116.550 76.760 ;
      LAYER li1 ;
        RECT 116.830 76.700 119.770 76.870 ;
        RECT 116.830 76.490 117.000 76.700 ;
        RECT 116.790 76.320 117.000 76.490 ;
        RECT 116.830 75.710 117.000 76.320 ;
      LAYER li1 ;
        RECT 115.510 75.180 116.040 75.410 ;
        RECT 115.510 73.870 115.760 75.180 ;
      LAYER li1 ;
        RECT 116.460 74.840 117.000 75.710 ;
        RECT 117.180 75.220 117.510 76.520 ;
      LAYER li1 ;
        RECT 117.690 76.000 117.960 76.500 ;
        RECT 118.410 76.250 118.740 76.500 ;
        RECT 118.410 76.080 119.420 76.250 ;
        RECT 117.690 75.010 117.860 76.000 ;
        RECT 118.740 75.410 119.070 75.900 ;
        RECT 117.640 74.840 117.860 75.010 ;
        RECT 118.040 75.180 119.070 75.410 ;
        RECT 119.250 75.850 119.420 76.080 ;
      LAYER li1 ;
        RECT 119.600 76.200 119.770 76.700 ;
      LAYER li1 ;
        RECT 120.920 76.760 120.950 76.930 ;
        RECT 121.120 76.760 121.310 76.930 ;
        RECT 121.480 76.760 121.670 76.930 ;
        RECT 121.840 76.760 121.870 76.930 ;
        RECT 120.920 76.380 121.870 76.760 ;
      LAYER li1 ;
        RECT 122.050 76.890 124.710 77.060 ;
        RECT 122.050 76.200 122.220 76.890 ;
        RECT 119.600 76.030 122.220 76.200 ;
      LAYER li1 ;
        RECT 119.250 75.680 121.870 75.850 ;
        RECT 117.640 74.660 117.810 74.840 ;
        RECT 118.040 74.660 118.210 75.180 ;
        RECT 119.250 75.000 119.420 75.680 ;
      LAYER li1 ;
        RECT 122.050 75.500 122.220 76.030 ;
      LAYER li1 ;
        RECT 116.000 74.490 117.810 74.660 ;
        RECT 116.000 73.870 116.250 74.490 ;
        RECT 116.430 74.140 117.460 74.310 ;
        RECT 116.430 73.690 116.600 74.140 ;
        RECT 112.090 73.570 113.540 73.600 ;
        RECT 115.160 73.520 116.600 73.690 ;
        RECT 116.780 73.820 117.110 73.960 ;
        RECT 116.780 73.650 116.810 73.820 ;
        RECT 116.980 73.650 117.110 73.820 ;
        RECT 116.780 73.620 117.110 73.650 ;
        RECT 117.290 73.690 117.460 74.140 ;
        RECT 117.640 73.870 117.810 74.490 ;
        RECT 117.990 74.330 118.210 74.660 ;
        RECT 118.390 74.830 119.420 75.000 ;
        RECT 119.600 75.150 119.930 75.500 ;
      LAYER li1 ;
        RECT 120.370 75.330 122.220 75.500 ;
      LAYER li1 ;
        RECT 122.400 76.000 122.730 76.710 ;
        RECT 123.190 76.540 124.360 76.710 ;
        RECT 123.190 76.000 123.520 76.540 ;
        RECT 122.400 75.150 122.660 76.000 ;
        RECT 123.730 75.740 124.010 76.240 ;
        RECT 119.600 74.980 122.660 75.150 ;
        RECT 118.390 74.130 118.560 74.830 ;
        RECT 119.250 74.800 119.420 74.830 ;
        RECT 118.740 74.450 119.070 74.650 ;
        RECT 119.250 74.630 121.020 74.800 ;
        RECT 118.740 74.330 120.510 74.450 ;
        RECT 118.860 74.280 120.510 74.330 ;
        RECT 118.340 73.870 118.670 74.130 ;
        RECT 118.860 73.690 119.030 74.280 ;
        RECT 117.290 73.520 119.030 73.690 ;
        RECT 119.210 73.820 120.160 74.100 ;
        RECT 119.210 73.650 119.240 73.820 ;
        RECT 119.410 73.650 119.600 73.820 ;
        RECT 119.770 73.650 119.960 73.820 ;
        RECT 120.130 73.650 120.160 73.820 ;
        RECT 119.210 73.620 120.160 73.650 ;
        RECT 120.340 73.690 120.510 74.280 ;
        RECT 120.690 73.870 121.020 74.630 ;
        RECT 122.330 74.400 122.660 74.980 ;
        RECT 122.840 75.570 124.010 75.740 ;
        RECT 122.840 74.220 123.010 75.570 ;
        RECT 123.390 74.890 123.720 75.390 ;
        RECT 124.190 75.140 124.360 76.540 ;
      LAYER li1 ;
        RECT 124.540 76.230 124.710 76.890 ;
      LAYER li1 ;
        RECT 124.890 76.930 125.840 76.960 ;
        RECT 124.890 76.760 124.920 76.930 ;
        RECT 125.090 76.760 125.280 76.930 ;
        RECT 125.450 76.760 125.640 76.930 ;
        RECT 125.810 76.760 125.840 76.930 ;
        RECT 127.500 76.930 128.450 76.960 ;
        RECT 124.890 76.410 125.840 76.760 ;
        RECT 126.380 76.330 126.710 76.830 ;
        RECT 127.500 76.760 127.530 76.930 ;
        RECT 127.700 76.760 127.890 76.930 ;
        RECT 128.060 76.760 128.250 76.930 ;
        RECT 128.420 76.760 128.450 76.930 ;
      LAYER li1 ;
        RECT 124.540 76.060 125.550 76.230 ;
      LAYER li1 ;
        RECT 124.570 75.490 124.900 75.880 ;
      LAYER li1 ;
        RECT 125.220 75.670 125.550 76.060 ;
      LAYER li1 ;
        RECT 126.380 75.490 126.610 76.330 ;
        RECT 126.990 75.830 127.320 76.330 ;
        RECT 127.500 75.830 128.450 76.760 ;
        RECT 129.700 76.940 132.430 76.970 ;
        RECT 129.700 76.770 129.870 76.940 ;
        RECT 130.040 76.770 130.310 76.940 ;
        RECT 130.480 76.770 130.720 76.940 ;
        RECT 130.890 76.770 131.150 76.940 ;
        RECT 131.320 76.770 131.590 76.940 ;
        RECT 131.760 76.770 132.000 76.940 ;
        RECT 132.170 76.770 132.430 76.940 ;
        RECT 135.940 76.930 136.590 77.040 ;
        RECT 129.700 75.970 132.430 76.770 ;
      LAYER li1 ;
        RECT 134.690 76.260 135.270 76.900 ;
      LAYER li1 ;
        RECT 135.940 76.760 136.000 76.930 ;
        RECT 136.170 76.760 136.360 76.930 ;
        RECT 136.530 76.760 136.590 76.930 ;
        RECT 135.940 76.700 136.590 76.760 ;
        RECT 136.180 76.260 136.590 76.700 ;
        RECT 137.380 76.940 140.110 76.970 ;
        RECT 137.380 76.770 137.550 76.940 ;
        RECT 137.720 76.770 137.990 76.940 ;
        RECT 138.160 76.770 138.400 76.940 ;
        RECT 138.570 76.770 138.830 76.940 ;
        RECT 139.000 76.770 139.270 76.940 ;
        RECT 139.440 76.770 139.680 76.940 ;
        RECT 139.850 76.770 140.110 76.940 ;
        RECT 124.570 75.320 126.610 75.490 ;
        RECT 123.900 74.970 126.260 75.140 ;
        RECT 123.900 74.650 124.070 74.970 ;
        RECT 126.440 74.790 126.610 75.320 ;
        RECT 121.200 74.050 123.010 74.220 ;
        RECT 123.190 74.480 124.070 74.650 ;
        RECT 121.200 73.690 121.370 74.050 ;
        RECT 120.340 73.520 121.370 73.690 ;
        RECT 121.550 73.820 122.500 73.870 ;
        RECT 121.550 73.650 121.580 73.820 ;
        RECT 121.750 73.650 121.940 73.820 ;
        RECT 122.110 73.650 122.300 73.820 ;
        RECT 122.470 73.650 122.500 73.820 ;
        RECT 121.550 73.570 122.500 73.650 ;
        RECT 123.190 73.570 123.440 74.480 ;
        RECT 124.250 73.820 125.200 74.650 ;
        RECT 125.600 74.620 126.610 74.790 ;
        RECT 127.110 75.650 127.320 75.830 ;
        RECT 127.110 75.320 128.480 75.650 ;
        RECT 125.600 74.150 125.850 74.620 ;
        RECT 126.030 73.820 126.930 74.440 ;
        RECT 127.110 74.320 127.360 75.320 ;
        RECT 129.860 75.300 130.190 75.970 ;
        RECT 124.250 73.650 124.280 73.820 ;
        RECT 124.450 73.650 124.640 73.820 ;
        RECT 124.810 73.650 125.000 73.820 ;
        RECT 125.170 73.650 125.200 73.820 ;
        RECT 126.200 73.650 126.390 73.820 ;
        RECT 126.560 73.650 126.750 73.820 ;
        RECT 126.920 73.650 126.930 73.820 ;
        RECT 124.250 73.620 125.200 73.650 ;
        RECT 126.030 73.620 126.930 73.650 ;
        RECT 127.540 73.820 128.480 75.130 ;
        RECT 130.590 74.650 130.920 75.630 ;
        RECT 131.140 75.300 131.470 75.970 ;
        RECT 131.870 74.650 132.200 75.630 ;
      LAYER li1 ;
        RECT 135.020 75.390 135.270 76.260 ;
      LAYER li1 ;
        RECT 137.380 75.970 140.110 76.770 ;
      LAYER li1 ;
        RECT 135.020 75.140 135.730 75.390 ;
      LAYER li1 ;
        RECT 137.540 75.300 137.870 75.970 ;
        RECT 127.540 73.650 127.560 73.820 ;
        RECT 127.730 73.650 127.920 73.820 ;
        RECT 128.090 73.650 128.280 73.820 ;
        RECT 128.450 73.650 128.480 73.820 ;
        RECT 127.540 73.590 128.480 73.650 ;
        RECT 129.620 73.770 132.360 74.650 ;
        RECT 129.620 73.600 129.830 73.770 ;
        RECT 130.000 73.600 130.270 73.770 ;
        RECT 130.440 73.600 130.680 73.770 ;
        RECT 130.850 73.600 131.110 73.770 ;
        RECT 131.280 73.600 131.550 73.770 ;
        RECT 131.720 73.600 131.960 73.770 ;
        RECT 132.130 73.600 132.360 73.770 ;
        RECT 129.620 73.580 132.360 73.600 ;
        RECT 134.620 73.880 135.020 74.150 ;
        RECT 134.620 73.820 135.270 73.880 ;
        RECT 134.620 73.650 134.680 73.820 ;
        RECT 134.850 73.650 135.040 73.820 ;
        RECT 135.210 73.650 135.270 73.820 ;
      LAYER li1 ;
        RECT 135.480 73.800 135.730 75.140 ;
      LAYER li1 ;
        RECT 138.270 74.650 138.600 75.630 ;
        RECT 138.820 75.300 139.150 75.970 ;
        RECT 139.550 74.650 139.880 75.630 ;
        RECT 134.620 73.540 135.270 73.650 ;
        RECT 137.300 73.770 140.040 74.650 ;
        RECT 137.300 73.600 137.510 73.770 ;
        RECT 137.680 73.600 137.950 73.770 ;
        RECT 138.120 73.600 138.360 73.770 ;
        RECT 138.530 73.600 138.790 73.770 ;
        RECT 138.960 73.600 139.230 73.770 ;
        RECT 139.400 73.600 139.640 73.770 ;
        RECT 139.810 73.600 140.040 73.770 ;
        RECT 137.300 73.580 140.040 73.600 ;
        RECT 5.760 73.170 5.920 73.350 ;
        RECT 6.090 73.170 6.400 73.350 ;
        RECT 6.570 73.170 6.880 73.350 ;
        RECT 7.050 73.170 7.360 73.350 ;
        RECT 7.530 73.170 7.840 73.350 ;
        RECT 8.010 73.170 8.320 73.350 ;
        RECT 8.490 73.170 8.800 73.350 ;
        RECT 8.970 73.170 9.280 73.350 ;
        RECT 9.450 73.170 9.760 73.350 ;
        RECT 9.930 73.170 10.240 73.350 ;
        RECT 10.410 73.170 10.720 73.350 ;
        RECT 10.890 73.170 11.200 73.350 ;
        RECT 11.370 73.170 11.680 73.350 ;
        RECT 11.850 73.170 12.160 73.350 ;
        RECT 12.330 73.170 12.640 73.350 ;
        RECT 12.810 73.170 13.120 73.350 ;
        RECT 13.290 73.170 13.600 73.350 ;
        RECT 13.770 73.170 14.080 73.350 ;
        RECT 14.250 73.170 14.560 73.350 ;
        RECT 14.730 73.170 15.040 73.350 ;
        RECT 15.210 73.170 15.520 73.350 ;
        RECT 15.690 73.170 16.000 73.350 ;
        RECT 16.170 73.170 16.480 73.350 ;
        RECT 16.650 73.170 16.960 73.350 ;
        RECT 17.130 73.170 17.440 73.350 ;
        RECT 17.610 73.170 17.920 73.350 ;
        RECT 18.090 73.170 18.400 73.350 ;
        RECT 18.570 73.170 18.880 73.350 ;
        RECT 19.050 73.170 19.360 73.350 ;
        RECT 19.530 73.170 19.840 73.350 ;
        RECT 20.010 73.170 20.320 73.350 ;
        RECT 20.490 73.170 20.800 73.350 ;
        RECT 20.970 73.170 21.280 73.350 ;
        RECT 21.450 73.170 21.760 73.350 ;
        RECT 21.930 73.170 22.240 73.350 ;
        RECT 22.410 73.170 22.720 73.350 ;
        RECT 22.890 73.170 23.200 73.350 ;
        RECT 23.370 73.170 23.680 73.350 ;
        RECT 23.850 73.170 24.160 73.350 ;
        RECT 24.330 73.170 24.640 73.350 ;
        RECT 24.810 73.170 25.120 73.350 ;
        RECT 25.290 73.170 25.600 73.350 ;
        RECT 25.770 73.170 26.080 73.350 ;
        RECT 26.250 73.170 26.560 73.350 ;
        RECT 26.730 73.170 27.040 73.350 ;
        RECT 27.210 73.170 27.520 73.350 ;
        RECT 27.690 73.170 28.000 73.350 ;
        RECT 28.170 73.170 28.480 73.350 ;
        RECT 28.650 73.170 28.960 73.350 ;
        RECT 29.130 73.170 29.440 73.350 ;
        RECT 29.610 73.170 29.920 73.350 ;
        RECT 30.090 73.170 30.400 73.350 ;
        RECT 30.570 73.170 30.880 73.350 ;
        RECT 31.050 73.170 31.360 73.350 ;
        RECT 31.530 73.170 31.840 73.350 ;
        RECT 32.010 73.170 32.320 73.350 ;
        RECT 32.490 73.170 32.800 73.350 ;
        RECT 32.970 73.170 33.280 73.350 ;
        RECT 33.450 73.170 33.760 73.350 ;
        RECT 33.930 73.170 34.240 73.350 ;
        RECT 34.410 73.170 34.720 73.350 ;
        RECT 34.890 73.170 35.200 73.350 ;
        RECT 35.370 73.170 35.680 73.350 ;
        RECT 35.850 73.170 36.160 73.350 ;
        RECT 36.330 73.170 36.640 73.350 ;
        RECT 36.810 73.170 37.120 73.350 ;
        RECT 37.290 73.170 37.600 73.350 ;
        RECT 37.770 73.170 38.080 73.350 ;
        RECT 38.250 73.170 38.560 73.350 ;
        RECT 38.730 73.170 39.040 73.350 ;
        RECT 39.210 73.170 39.520 73.350 ;
        RECT 39.690 73.170 40.000 73.350 ;
        RECT 40.170 73.170 40.480 73.350 ;
        RECT 40.650 73.170 40.960 73.350 ;
        RECT 41.130 73.170 41.440 73.350 ;
        RECT 41.610 73.170 41.920 73.350 ;
        RECT 42.090 73.170 42.400 73.350 ;
        RECT 42.570 73.170 42.880 73.350 ;
        RECT 43.050 73.170 43.360 73.350 ;
        RECT 43.530 73.170 43.840 73.350 ;
        RECT 44.010 73.170 44.320 73.350 ;
        RECT 44.490 73.170 44.800 73.350 ;
        RECT 44.970 73.170 45.280 73.350 ;
        RECT 45.450 73.170 45.760 73.350 ;
        RECT 45.930 73.170 46.240 73.350 ;
        RECT 46.410 73.170 46.720 73.350 ;
        RECT 46.890 73.340 47.200 73.350 ;
        RECT 47.370 73.340 47.520 73.350 ;
        RECT 48.000 73.340 48.160 73.350 ;
        RECT 46.890 73.170 47.040 73.340 ;
        RECT 47.520 73.170 47.680 73.340 ;
        RECT 47.850 73.170 48.160 73.340 ;
        RECT 48.330 73.170 48.640 73.350 ;
        RECT 48.810 73.170 49.120 73.350 ;
        RECT 49.290 73.170 49.600 73.350 ;
        RECT 49.770 73.170 50.080 73.350 ;
        RECT 50.250 73.170 50.560 73.350 ;
        RECT 50.730 73.170 51.040 73.350 ;
        RECT 51.210 73.170 51.520 73.350 ;
        RECT 51.690 73.170 52.000 73.350 ;
        RECT 52.170 73.170 52.480 73.350 ;
        RECT 52.650 73.170 52.960 73.350 ;
        RECT 53.130 73.170 53.440 73.350 ;
        RECT 53.610 73.170 53.920 73.350 ;
        RECT 54.090 73.170 54.400 73.350 ;
        RECT 54.570 73.170 54.880 73.350 ;
        RECT 55.050 73.170 55.360 73.350 ;
        RECT 55.530 73.170 55.840 73.350 ;
        RECT 56.010 73.170 56.320 73.350 ;
        RECT 56.490 73.170 56.800 73.350 ;
        RECT 56.970 73.170 57.280 73.350 ;
        RECT 57.450 73.170 57.760 73.350 ;
        RECT 57.930 73.170 58.240 73.350 ;
        RECT 58.410 73.170 58.720 73.350 ;
        RECT 58.890 73.340 59.040 73.350 ;
        RECT 59.520 73.340 59.680 73.350 ;
        RECT 58.890 73.170 59.200 73.340 ;
        RECT 59.370 73.170 59.680 73.340 ;
        RECT 59.850 73.170 60.160 73.350 ;
        RECT 60.330 73.170 60.640 73.350 ;
        RECT 60.810 73.170 61.120 73.350 ;
        RECT 61.290 73.170 61.600 73.350 ;
        RECT 61.770 73.170 62.080 73.350 ;
        RECT 62.250 73.170 62.560 73.350 ;
        RECT 62.730 73.170 63.040 73.350 ;
        RECT 63.210 73.170 63.520 73.350 ;
        RECT 63.690 73.170 64.000 73.350 ;
        RECT 64.170 73.170 64.480 73.350 ;
        RECT 64.650 73.170 64.960 73.350 ;
        RECT 65.130 73.170 65.440 73.350 ;
        RECT 65.610 73.170 65.920 73.350 ;
        RECT 66.090 73.170 66.400 73.350 ;
        RECT 66.570 73.170 66.880 73.350 ;
        RECT 67.050 73.170 67.360 73.350 ;
        RECT 67.530 73.170 67.840 73.350 ;
        RECT 68.010 73.170 68.320 73.350 ;
        RECT 68.490 73.170 68.800 73.350 ;
        RECT 68.970 73.170 69.280 73.350 ;
        RECT 69.450 73.170 69.760 73.350 ;
        RECT 69.930 73.170 70.240 73.350 ;
        RECT 70.410 73.170 70.720 73.350 ;
        RECT 70.890 73.170 71.200 73.350 ;
        RECT 71.370 73.170 71.680 73.350 ;
        RECT 71.850 73.170 72.160 73.350 ;
        RECT 72.330 73.170 72.640 73.350 ;
        RECT 72.810 73.170 73.120 73.350 ;
        RECT 73.290 73.170 73.600 73.350 ;
        RECT 73.770 73.170 74.080 73.350 ;
        RECT 74.250 73.170 74.560 73.350 ;
        RECT 74.730 73.170 75.040 73.350 ;
        RECT 75.210 73.170 75.520 73.350 ;
        RECT 75.690 73.170 76.000 73.350 ;
        RECT 76.170 73.340 76.320 73.350 ;
        RECT 76.800 73.340 76.960 73.350 ;
        RECT 76.170 73.170 76.480 73.340 ;
        RECT 76.650 73.170 76.960 73.340 ;
        RECT 77.130 73.170 77.440 73.350 ;
        RECT 77.610 73.170 77.920 73.350 ;
        RECT 78.090 73.170 78.400 73.350 ;
        RECT 78.570 73.340 78.880 73.350 ;
        RECT 79.050 73.340 79.360 73.350 ;
        RECT 78.570 73.170 78.720 73.340 ;
        RECT 79.200 73.170 79.360 73.340 ;
        RECT 79.530 73.170 79.840 73.350 ;
        RECT 80.010 73.170 80.320 73.350 ;
        RECT 80.490 73.170 80.800 73.350 ;
        RECT 80.970 73.170 81.280 73.350 ;
        RECT 81.450 73.170 81.760 73.350 ;
        RECT 81.930 73.170 82.240 73.350 ;
        RECT 82.410 73.170 82.720 73.350 ;
        RECT 82.890 73.170 83.200 73.350 ;
        RECT 83.370 73.170 83.680 73.350 ;
        RECT 83.850 73.170 84.160 73.350 ;
        RECT 84.330 73.170 84.640 73.350 ;
        RECT 84.810 73.170 85.120 73.350 ;
        RECT 85.290 73.170 85.600 73.350 ;
        RECT 85.770 73.170 86.080 73.350 ;
        RECT 86.250 73.170 86.560 73.350 ;
        RECT 86.730 73.170 87.040 73.350 ;
        RECT 87.210 73.170 87.520 73.350 ;
        RECT 87.690 73.170 88.000 73.350 ;
        RECT 88.170 73.170 88.480 73.350 ;
        RECT 88.650 73.170 88.960 73.350 ;
        RECT 89.130 73.170 89.440 73.350 ;
        RECT 89.610 73.170 89.920 73.350 ;
        RECT 90.090 73.170 90.400 73.350 ;
        RECT 90.570 73.170 90.880 73.350 ;
        RECT 91.050 73.170 91.360 73.350 ;
        RECT 91.530 73.170 91.840 73.350 ;
        RECT 92.010 73.170 92.320 73.350 ;
        RECT 92.490 73.170 92.800 73.350 ;
        RECT 92.970 73.170 93.280 73.350 ;
        RECT 93.450 73.170 93.760 73.350 ;
        RECT 93.930 73.170 94.240 73.350 ;
        RECT 94.410 73.170 94.720 73.350 ;
        RECT 94.890 73.170 95.200 73.350 ;
        RECT 95.370 73.170 95.680 73.350 ;
        RECT 95.850 73.170 96.160 73.350 ;
        RECT 96.330 73.170 96.640 73.350 ;
        RECT 96.810 73.170 97.120 73.350 ;
        RECT 97.290 73.170 97.600 73.350 ;
        RECT 97.770 73.170 98.080 73.350 ;
        RECT 98.250 73.170 98.560 73.350 ;
        RECT 98.730 73.170 99.040 73.350 ;
        RECT 99.210 73.170 99.520 73.350 ;
        RECT 99.690 73.170 100.000 73.350 ;
        RECT 100.170 73.170 100.480 73.350 ;
        RECT 100.650 73.170 100.960 73.350 ;
        RECT 101.130 73.170 101.440 73.350 ;
        RECT 101.610 73.170 101.920 73.350 ;
        RECT 102.090 73.170 102.400 73.350 ;
        RECT 102.570 73.170 102.880 73.350 ;
        RECT 103.050 73.170 103.360 73.350 ;
        RECT 103.530 73.170 103.840 73.350 ;
        RECT 104.010 73.170 104.320 73.350 ;
        RECT 104.490 73.170 104.800 73.350 ;
        RECT 104.970 73.170 105.280 73.350 ;
        RECT 105.450 73.170 105.760 73.350 ;
        RECT 105.930 73.170 106.240 73.350 ;
        RECT 106.410 73.170 106.720 73.350 ;
        RECT 106.890 73.170 107.200 73.350 ;
        RECT 107.370 73.170 107.680 73.350 ;
        RECT 107.850 73.170 108.160 73.350 ;
        RECT 108.330 73.170 108.640 73.350 ;
        RECT 108.810 73.170 109.120 73.350 ;
        RECT 109.290 73.170 109.600 73.350 ;
        RECT 109.770 73.170 110.080 73.350 ;
        RECT 110.250 73.170 110.560 73.350 ;
        RECT 110.730 73.170 111.040 73.350 ;
        RECT 111.210 73.170 111.520 73.350 ;
        RECT 111.690 73.170 112.000 73.350 ;
        RECT 112.170 73.170 112.480 73.350 ;
        RECT 112.650 73.170 112.960 73.350 ;
        RECT 113.130 73.170 113.440 73.350 ;
        RECT 113.610 73.170 113.920 73.350 ;
        RECT 114.090 73.170 114.400 73.350 ;
        RECT 114.570 73.170 114.880 73.350 ;
        RECT 115.050 73.170 115.360 73.350 ;
        RECT 115.530 73.170 115.840 73.350 ;
        RECT 116.010 73.170 116.320 73.350 ;
        RECT 116.490 73.170 116.800 73.350 ;
        RECT 116.970 73.170 117.280 73.350 ;
        RECT 117.450 73.170 117.760 73.350 ;
        RECT 117.930 73.170 118.240 73.350 ;
        RECT 118.410 73.170 118.720 73.350 ;
        RECT 118.890 73.170 119.200 73.350 ;
        RECT 119.370 73.170 119.680 73.350 ;
        RECT 119.850 73.170 120.160 73.350 ;
        RECT 120.330 73.170 120.640 73.350 ;
        RECT 120.810 73.170 121.120 73.350 ;
        RECT 121.290 73.170 121.600 73.350 ;
        RECT 121.770 73.170 122.080 73.350 ;
        RECT 122.250 73.170 122.560 73.350 ;
        RECT 122.730 73.170 123.040 73.350 ;
        RECT 123.210 73.170 123.520 73.350 ;
        RECT 123.690 73.170 124.000 73.350 ;
        RECT 124.170 73.170 124.480 73.350 ;
        RECT 124.650 73.170 124.960 73.350 ;
        RECT 125.130 73.170 125.440 73.350 ;
        RECT 125.610 73.170 125.920 73.350 ;
        RECT 126.090 73.170 126.400 73.350 ;
        RECT 126.570 73.170 126.880 73.350 ;
        RECT 127.050 73.170 127.360 73.350 ;
        RECT 127.530 73.170 127.840 73.350 ;
        RECT 128.010 73.170 128.320 73.350 ;
        RECT 128.490 73.170 128.800 73.350 ;
        RECT 128.970 73.170 129.280 73.350 ;
        RECT 129.450 73.170 129.760 73.350 ;
        RECT 129.930 73.170 130.240 73.350 ;
        RECT 130.410 73.170 130.720 73.350 ;
        RECT 130.890 73.170 131.200 73.350 ;
        RECT 131.370 73.170 131.680 73.350 ;
        RECT 131.850 73.170 132.160 73.350 ;
        RECT 132.330 73.170 132.640 73.350 ;
        RECT 132.810 73.170 133.120 73.350 ;
        RECT 133.290 73.170 133.600 73.350 ;
        RECT 133.770 73.340 134.080 73.350 ;
        RECT 134.250 73.340 134.560 73.350 ;
        RECT 133.770 73.170 133.920 73.340 ;
        RECT 134.400 73.170 134.560 73.340 ;
        RECT 134.730 73.170 135.040 73.350 ;
        RECT 135.210 73.170 135.520 73.350 ;
        RECT 135.690 73.170 136.000 73.350 ;
        RECT 136.170 73.170 136.480 73.350 ;
        RECT 136.650 73.170 136.960 73.350 ;
        RECT 137.130 73.170 137.440 73.350 ;
        RECT 137.610 73.170 137.920 73.350 ;
        RECT 138.090 73.170 138.400 73.350 ;
        RECT 138.570 73.170 138.880 73.350 ;
        RECT 139.050 73.170 139.360 73.350 ;
        RECT 139.530 73.170 139.840 73.350 ;
        RECT 140.010 73.170 140.320 73.350 ;
        RECT 140.490 73.170 140.800 73.350 ;
        RECT 140.970 73.170 141.280 73.350 ;
        RECT 141.450 73.340 141.760 73.350 ;
        RECT 141.930 73.340 142.080 73.350 ;
        RECT 141.450 73.170 141.600 73.340 ;
        RECT 6.260 72.920 9.000 72.940 ;
        RECT 6.260 72.750 6.470 72.920 ;
        RECT 6.640 72.750 6.910 72.920 ;
        RECT 7.080 72.750 7.320 72.920 ;
        RECT 7.490 72.750 7.750 72.920 ;
        RECT 7.920 72.750 8.190 72.920 ;
        RECT 8.360 72.750 8.600 72.920 ;
        RECT 8.770 72.750 9.000 72.920 ;
        RECT 6.260 71.870 9.000 72.750 ;
        RECT 9.850 72.920 11.300 72.950 ;
        RECT 9.850 72.750 10.100 72.920 ;
        RECT 10.270 72.750 10.460 72.920 ;
        RECT 10.630 72.750 10.900 72.920 ;
        RECT 11.070 72.750 11.300 72.920 ;
        RECT 9.850 71.880 11.300 72.750 ;
        RECT 6.500 70.550 6.830 71.220 ;
        RECT 7.230 70.890 7.560 71.870 ;
        RECT 7.780 70.550 8.110 71.220 ;
        RECT 8.510 70.890 8.840 71.870 ;
        RECT 6.340 69.550 9.070 70.550 ;
        RECT 10.080 70.440 10.410 71.220 ;
        RECT 10.620 70.890 10.950 71.880 ;
      LAYER li1 ;
        RECT 12.600 71.370 13.030 72.950 ;
      LAYER li1 ;
        RECT 13.210 72.870 13.770 72.950 ;
        RECT 13.210 72.700 13.220 72.870 ;
        RECT 13.390 72.700 13.580 72.870 ;
        RECT 13.750 72.700 13.770 72.870 ;
        RECT 13.210 71.370 13.770 72.700 ;
        RECT 15.130 72.920 16.580 72.950 ;
        RECT 15.130 72.750 15.380 72.920 ;
        RECT 15.550 72.750 15.740 72.920 ;
        RECT 15.910 72.750 16.180 72.920 ;
        RECT 16.350 72.750 16.580 72.920 ;
        RECT 10.080 70.040 11.380 70.440 ;
        RECT 9.770 69.560 11.380 70.040 ;
      LAYER li1 ;
        RECT 12.600 69.690 12.850 71.370 ;
      LAYER li1 ;
        RECT 13.160 70.480 13.490 70.940 ;
      LAYER li1 ;
        RECT 13.950 70.660 14.280 72.450 ;
      LAYER li1 ;
        RECT 14.460 70.480 14.710 72.200 ;
        RECT 15.130 71.880 16.580 72.750 ;
        RECT 13.160 70.310 14.710 70.480 ;
        RECT 13.030 69.560 14.280 70.130 ;
        RECT 14.460 69.690 14.710 70.310 ;
        RECT 15.360 70.440 15.690 71.220 ;
        RECT 15.900 70.890 16.230 71.880 ;
      LAYER li1 ;
        RECT 16.920 71.370 17.350 72.950 ;
      LAYER li1 ;
        RECT 17.530 72.870 18.090 72.950 ;
        RECT 17.530 72.700 17.540 72.870 ;
        RECT 17.710 72.700 17.900 72.870 ;
        RECT 18.070 72.700 18.090 72.870 ;
        RECT 17.530 71.370 18.090 72.700 ;
        RECT 19.450 72.920 20.900 72.950 ;
        RECT 19.450 72.750 19.700 72.920 ;
        RECT 19.870 72.750 20.060 72.920 ;
        RECT 20.230 72.750 20.500 72.920 ;
        RECT 20.670 72.750 20.900 72.920 ;
        RECT 15.360 70.040 16.660 70.440 ;
        RECT 15.050 69.560 16.660 70.040 ;
      LAYER li1 ;
        RECT 16.920 69.690 17.170 71.370 ;
      LAYER li1 ;
        RECT 17.480 70.480 17.810 70.940 ;
      LAYER li1 ;
        RECT 18.270 70.660 18.600 72.450 ;
      LAYER li1 ;
        RECT 18.780 70.480 19.030 72.200 ;
        RECT 19.450 71.880 20.900 72.750 ;
        RECT 17.480 70.310 19.030 70.480 ;
        RECT 17.350 69.560 18.600 70.130 ;
        RECT 18.780 69.690 19.030 70.310 ;
        RECT 19.680 70.440 20.010 71.220 ;
        RECT 20.220 70.890 20.550 71.880 ;
        RECT 21.380 71.290 21.630 72.950 ;
        RECT 21.810 72.870 23.060 72.950 ;
        RECT 21.980 72.700 22.170 72.870 ;
        RECT 22.340 72.700 22.530 72.870 ;
        RECT 22.700 72.700 22.890 72.870 ;
        RECT 21.810 71.470 23.060 72.700 ;
        RECT 23.240 71.290 23.410 72.950 ;
        RECT 21.380 71.120 23.410 71.290 ;
      LAYER li1 ;
        RECT 23.590 71.000 23.920 72.450 ;
        RECT 21.250 70.700 22.440 70.940 ;
        RECT 22.690 70.700 23.040 70.940 ;
        RECT 24.100 70.820 24.360 72.950 ;
      LAYER li1 ;
        RECT 24.730 72.920 26.180 72.950 ;
        RECT 24.730 72.750 24.980 72.920 ;
        RECT 25.150 72.750 25.340 72.920 ;
        RECT 25.510 72.750 25.780 72.920 ;
        RECT 25.950 72.750 26.180 72.920 ;
        RECT 24.730 71.880 26.180 72.750 ;
        RECT 26.490 72.870 27.440 72.950 ;
        RECT 26.490 72.700 26.520 72.870 ;
        RECT 26.690 72.700 26.880 72.870 ;
        RECT 27.050 72.700 27.240 72.870 ;
        RECT 27.410 72.700 27.440 72.870 ;
      LAYER li1 ;
        RECT 23.340 70.650 24.360 70.820 ;
      LAYER li1 ;
        RECT 19.680 70.040 20.980 70.440 ;
        RECT 19.370 69.560 20.980 70.040 ;
        RECT 21.450 69.560 23.160 70.520 ;
      LAYER li1 ;
        RECT 23.340 69.690 23.590 70.650 ;
      LAYER li1 ;
        RECT 23.800 69.560 24.390 70.470 ;
        RECT 24.960 70.440 25.290 71.220 ;
        RECT 25.500 70.890 25.830 71.880 ;
        RECT 26.490 71.370 27.440 72.700 ;
      LAYER li1 ;
        RECT 27.620 71.270 27.870 72.950 ;
      LAYER li1 ;
        RECT 28.050 72.870 29.000 72.950 ;
        RECT 28.050 72.700 28.080 72.870 ;
        RECT 28.250 72.700 28.440 72.870 ;
        RECT 28.610 72.700 28.800 72.870 ;
        RECT 28.970 72.700 29.000 72.870 ;
        RECT 28.050 71.450 29.000 72.700 ;
      LAYER li1 ;
        RECT 29.180 71.270 29.510 72.950 ;
      LAYER li1 ;
        RECT 29.690 72.870 30.640 72.950 ;
        RECT 29.690 72.700 29.720 72.870 ;
        RECT 29.890 72.700 30.080 72.870 ;
        RECT 30.250 72.700 30.440 72.870 ;
        RECT 30.610 72.700 30.640 72.870 ;
        RECT 29.690 71.490 30.640 72.700 ;
      LAYER li1 ;
        RECT 27.620 71.100 29.510 71.270 ;
        RECT 27.620 70.970 27.790 71.100 ;
        RECT 30.290 70.970 30.620 71.310 ;
        RECT 26.530 70.740 27.790 70.970 ;
      LAYER li1 ;
        RECT 27.970 70.790 30.000 70.920 ;
        RECT 30.820 70.790 31.070 72.950 ;
        RECT 31.450 72.920 32.900 72.950 ;
        RECT 31.450 72.750 31.700 72.920 ;
        RECT 31.870 72.750 32.060 72.920 ;
        RECT 32.230 72.750 32.500 72.920 ;
        RECT 32.670 72.750 32.900 72.920 ;
        RECT 31.450 71.880 32.900 72.750 ;
        RECT 33.210 72.870 34.160 72.950 ;
        RECT 33.210 72.700 33.240 72.870 ;
        RECT 33.410 72.700 33.600 72.870 ;
        RECT 33.770 72.700 33.960 72.870 ;
        RECT 34.130 72.700 34.160 72.870 ;
        RECT 27.970 70.750 31.070 70.790 ;
      LAYER li1 ;
        RECT 27.620 70.570 27.790 70.740 ;
      LAYER li1 ;
        RECT 29.830 70.620 31.070 70.750 ;
        RECT 24.960 70.040 26.260 70.440 ;
        RECT 24.650 69.560 26.260 70.040 ;
        RECT 26.490 69.560 27.440 70.520 ;
      LAYER li1 ;
        RECT 27.620 70.400 29.430 70.570 ;
        RECT 27.620 69.690 27.870 70.400 ;
      LAYER li1 ;
        RECT 28.050 69.560 29.000 70.220 ;
      LAYER li1 ;
        RECT 29.180 69.690 29.430 70.400 ;
      LAYER li1 ;
        RECT 29.610 69.560 30.560 70.440 ;
        RECT 30.740 69.690 31.070 70.620 ;
        RECT 31.680 70.440 32.010 71.220 ;
        RECT 32.220 70.890 32.550 71.880 ;
        RECT 33.210 71.370 34.160 72.700 ;
      LAYER li1 ;
        RECT 34.340 71.270 34.590 72.950 ;
      LAYER li1 ;
        RECT 34.770 72.870 35.720 72.950 ;
        RECT 34.770 72.700 34.800 72.870 ;
        RECT 34.970 72.700 35.160 72.870 ;
        RECT 35.330 72.700 35.520 72.870 ;
        RECT 35.690 72.700 35.720 72.870 ;
        RECT 34.770 71.450 35.720 72.700 ;
      LAYER li1 ;
        RECT 35.900 71.270 36.230 72.950 ;
      LAYER li1 ;
        RECT 36.410 72.870 37.360 72.950 ;
        RECT 36.410 72.700 36.440 72.870 ;
        RECT 36.610 72.700 36.800 72.870 ;
        RECT 36.970 72.700 37.160 72.870 ;
        RECT 37.330 72.700 37.360 72.870 ;
        RECT 36.410 71.490 37.360 72.700 ;
      LAYER li1 ;
        RECT 34.340 71.100 36.230 71.270 ;
        RECT 34.340 70.970 34.510 71.100 ;
        RECT 37.010 70.970 37.340 71.310 ;
        RECT 33.250 70.740 34.510 70.970 ;
      LAYER li1 ;
        RECT 34.690 70.790 36.720 70.920 ;
        RECT 37.540 70.790 37.790 72.950 ;
        RECT 38.170 72.920 39.620 72.950 ;
        RECT 38.170 72.750 38.420 72.920 ;
        RECT 38.590 72.750 38.780 72.920 ;
        RECT 38.950 72.750 39.220 72.920 ;
        RECT 39.390 72.750 39.620 72.920 ;
        RECT 38.170 71.880 39.620 72.750 ;
        RECT 39.930 72.870 40.880 72.950 ;
        RECT 39.930 72.700 39.960 72.870 ;
        RECT 40.130 72.700 40.320 72.870 ;
        RECT 40.490 72.700 40.680 72.870 ;
        RECT 40.850 72.700 40.880 72.870 ;
        RECT 34.690 70.750 37.790 70.790 ;
      LAYER li1 ;
        RECT 34.340 70.570 34.510 70.740 ;
      LAYER li1 ;
        RECT 36.550 70.620 37.790 70.750 ;
        RECT 31.680 70.040 32.980 70.440 ;
        RECT 31.370 69.560 32.980 70.040 ;
        RECT 33.210 69.560 34.160 70.520 ;
      LAYER li1 ;
        RECT 34.340 70.400 36.150 70.570 ;
        RECT 34.340 69.690 34.590 70.400 ;
      LAYER li1 ;
        RECT 34.770 69.560 35.720 70.220 ;
      LAYER li1 ;
        RECT 35.900 69.690 36.150 70.400 ;
      LAYER li1 ;
        RECT 36.330 69.560 37.280 70.440 ;
        RECT 37.460 69.690 37.790 70.620 ;
        RECT 38.400 70.440 38.730 71.220 ;
        RECT 38.940 70.890 39.270 71.880 ;
        RECT 39.930 71.370 40.880 72.700 ;
      LAYER li1 ;
        RECT 41.060 71.270 41.310 72.950 ;
      LAYER li1 ;
        RECT 41.490 72.870 42.440 72.950 ;
        RECT 41.490 72.700 41.520 72.870 ;
        RECT 41.690 72.700 41.880 72.870 ;
        RECT 42.050 72.700 42.240 72.870 ;
        RECT 42.410 72.700 42.440 72.870 ;
        RECT 41.490 71.450 42.440 72.700 ;
      LAYER li1 ;
        RECT 42.620 71.270 42.950 72.950 ;
      LAYER li1 ;
        RECT 43.130 72.870 44.080 72.950 ;
        RECT 43.130 72.700 43.160 72.870 ;
        RECT 43.330 72.700 43.520 72.870 ;
        RECT 43.690 72.700 43.880 72.870 ;
        RECT 44.050 72.700 44.080 72.870 ;
        RECT 43.130 71.490 44.080 72.700 ;
      LAYER li1 ;
        RECT 41.060 71.100 42.950 71.270 ;
        RECT 41.060 70.970 41.230 71.100 ;
        RECT 43.730 70.970 44.060 71.310 ;
        RECT 39.970 70.740 41.230 70.970 ;
      LAYER li1 ;
        RECT 41.410 70.790 43.440 70.920 ;
        RECT 44.260 70.790 44.510 72.950 ;
        RECT 44.890 72.920 46.340 72.950 ;
        RECT 44.890 72.750 45.140 72.920 ;
        RECT 45.310 72.750 45.500 72.920 ;
        RECT 45.670 72.750 45.940 72.920 ;
        RECT 46.110 72.750 46.340 72.920 ;
        RECT 44.890 71.880 46.340 72.750 ;
        RECT 48.090 72.870 49.040 72.950 ;
        RECT 48.090 72.700 48.120 72.870 ;
        RECT 48.290 72.700 48.480 72.870 ;
        RECT 48.650 72.700 48.840 72.870 ;
        RECT 49.010 72.700 49.040 72.870 ;
        RECT 41.410 70.750 44.510 70.790 ;
      LAYER li1 ;
        RECT 41.060 70.570 41.230 70.740 ;
      LAYER li1 ;
        RECT 43.270 70.620 44.510 70.750 ;
        RECT 38.400 70.040 39.700 70.440 ;
        RECT 38.090 69.560 39.700 70.040 ;
        RECT 39.930 69.560 40.880 70.520 ;
      LAYER li1 ;
        RECT 41.060 70.400 42.870 70.570 ;
        RECT 41.060 69.690 41.310 70.400 ;
      LAYER li1 ;
        RECT 41.490 69.560 42.440 70.220 ;
      LAYER li1 ;
        RECT 42.620 69.690 42.870 70.400 ;
      LAYER li1 ;
        RECT 43.050 69.560 44.000 70.440 ;
        RECT 44.180 69.690 44.510 70.620 ;
        RECT 45.120 70.440 45.450 71.220 ;
        RECT 45.660 70.890 45.990 71.880 ;
        RECT 48.090 71.370 49.040 72.700 ;
      LAYER li1 ;
        RECT 49.220 71.270 49.470 72.950 ;
      LAYER li1 ;
        RECT 49.650 72.870 50.600 72.950 ;
        RECT 49.650 72.700 49.680 72.870 ;
        RECT 49.850 72.700 50.040 72.870 ;
        RECT 50.210 72.700 50.400 72.870 ;
        RECT 50.570 72.700 50.600 72.870 ;
        RECT 49.650 71.450 50.600 72.700 ;
      LAYER li1 ;
        RECT 50.780 71.270 51.110 72.950 ;
      LAYER li1 ;
        RECT 51.290 72.870 52.240 72.950 ;
        RECT 51.290 72.700 51.320 72.870 ;
        RECT 51.490 72.700 51.680 72.870 ;
        RECT 51.850 72.700 52.040 72.870 ;
        RECT 52.210 72.700 52.240 72.870 ;
        RECT 51.290 71.490 52.240 72.700 ;
      LAYER li1 ;
        RECT 49.220 71.100 51.110 71.270 ;
        RECT 49.220 70.970 49.390 71.100 ;
        RECT 51.890 70.970 52.220 71.310 ;
        RECT 48.130 70.740 49.390 70.970 ;
      LAYER li1 ;
        RECT 49.570 70.790 51.600 70.920 ;
        RECT 52.420 70.790 52.670 72.950 ;
        RECT 53.050 72.920 54.500 72.950 ;
        RECT 53.050 72.750 53.300 72.920 ;
        RECT 53.470 72.750 53.660 72.920 ;
        RECT 53.830 72.750 54.100 72.920 ;
        RECT 54.270 72.750 54.500 72.920 ;
        RECT 53.050 71.880 54.500 72.750 ;
        RECT 54.810 72.870 56.480 72.950 ;
        RECT 54.810 72.700 54.840 72.870 ;
        RECT 55.010 72.700 55.200 72.870 ;
        RECT 55.370 72.700 55.560 72.870 ;
        RECT 55.730 72.700 55.920 72.870 ;
        RECT 56.090 72.700 56.280 72.870 ;
        RECT 56.450 72.700 56.480 72.870 ;
        RECT 49.570 70.750 52.670 70.790 ;
      LAYER li1 ;
        RECT 49.220 70.570 49.390 70.740 ;
      LAYER li1 ;
        RECT 51.430 70.620 52.670 70.750 ;
        RECT 45.120 70.040 46.420 70.440 ;
        RECT 44.810 69.560 46.420 70.040 ;
        RECT 48.090 69.560 49.040 70.520 ;
      LAYER li1 ;
        RECT 49.220 70.400 51.030 70.570 ;
        RECT 49.220 69.690 49.470 70.400 ;
      LAYER li1 ;
        RECT 49.650 69.560 50.600 70.220 ;
      LAYER li1 ;
        RECT 50.780 69.690 51.030 70.400 ;
      LAYER li1 ;
        RECT 51.210 69.560 52.160 70.440 ;
        RECT 52.340 69.690 52.670 70.620 ;
        RECT 53.280 70.440 53.610 71.220 ;
        RECT 53.820 70.890 54.150 71.880 ;
        RECT 54.810 71.490 56.480 72.700 ;
      LAYER li1 ;
        RECT 54.850 70.970 56.040 71.310 ;
        RECT 56.220 70.970 56.550 71.310 ;
        RECT 56.740 70.790 57.000 72.950 ;
      LAYER li1 ;
        RECT 57.370 72.920 58.820 72.950 ;
        RECT 57.370 72.750 57.620 72.920 ;
        RECT 57.790 72.750 57.980 72.920 ;
        RECT 58.150 72.750 58.420 72.920 ;
        RECT 58.590 72.750 58.820 72.920 ;
        RECT 57.370 71.880 58.820 72.750 ;
        RECT 59.610 72.870 60.560 72.950 ;
        RECT 59.610 72.700 59.640 72.870 ;
        RECT 59.810 72.700 60.000 72.870 ;
        RECT 60.170 72.700 60.360 72.870 ;
        RECT 60.530 72.700 60.560 72.870 ;
      LAYER li1 ;
        RECT 55.920 70.620 57.000 70.790 ;
      LAYER li1 ;
        RECT 53.280 70.040 54.580 70.440 ;
        RECT 52.970 69.560 54.580 70.040 ;
        RECT 54.810 69.560 55.740 70.520 ;
      LAYER li1 ;
        RECT 55.920 69.690 56.250 70.620 ;
      LAYER li1 ;
        RECT 57.600 70.440 57.930 71.220 ;
        RECT 58.140 70.890 58.470 71.880 ;
        RECT 59.610 71.370 60.560 72.700 ;
      LAYER li1 ;
        RECT 60.740 71.270 60.990 72.950 ;
      LAYER li1 ;
        RECT 61.170 72.870 62.120 72.950 ;
        RECT 61.170 72.700 61.200 72.870 ;
        RECT 61.370 72.700 61.560 72.870 ;
        RECT 61.730 72.700 61.920 72.870 ;
        RECT 62.090 72.700 62.120 72.870 ;
        RECT 61.170 71.450 62.120 72.700 ;
      LAYER li1 ;
        RECT 62.300 71.270 62.630 72.950 ;
      LAYER li1 ;
        RECT 62.810 72.870 63.760 72.950 ;
        RECT 62.810 72.700 62.840 72.870 ;
        RECT 63.010 72.700 63.200 72.870 ;
        RECT 63.370 72.700 63.560 72.870 ;
        RECT 63.730 72.700 63.760 72.870 ;
        RECT 62.810 71.490 63.760 72.700 ;
      LAYER li1 ;
        RECT 60.740 71.100 62.630 71.270 ;
        RECT 60.740 70.970 60.910 71.100 ;
        RECT 63.410 70.970 63.740 71.310 ;
        RECT 59.650 70.740 60.910 70.970 ;
      LAYER li1 ;
        RECT 61.090 70.790 63.120 70.920 ;
        RECT 63.940 70.790 64.190 72.950 ;
        RECT 64.570 72.920 66.020 72.950 ;
        RECT 64.570 72.750 64.820 72.920 ;
        RECT 64.990 72.750 65.180 72.920 ;
        RECT 65.350 72.750 65.620 72.920 ;
        RECT 65.790 72.750 66.020 72.920 ;
        RECT 64.570 71.880 66.020 72.750 ;
        RECT 66.330 72.870 67.280 72.950 ;
        RECT 66.330 72.700 66.360 72.870 ;
        RECT 66.530 72.700 66.720 72.870 ;
        RECT 66.890 72.700 67.080 72.870 ;
        RECT 67.250 72.700 67.280 72.870 ;
        RECT 61.090 70.750 64.190 70.790 ;
      LAYER li1 ;
        RECT 60.740 70.570 60.910 70.740 ;
      LAYER li1 ;
        RECT 62.950 70.620 64.190 70.750 ;
        RECT 56.440 69.560 57.030 70.440 ;
        RECT 57.600 70.040 58.900 70.440 ;
        RECT 57.290 69.560 58.900 70.040 ;
        RECT 59.610 69.560 60.560 70.520 ;
      LAYER li1 ;
        RECT 60.740 70.400 62.550 70.570 ;
        RECT 60.740 69.690 60.990 70.400 ;
      LAYER li1 ;
        RECT 61.170 69.560 62.120 70.220 ;
      LAYER li1 ;
        RECT 62.300 69.690 62.550 70.400 ;
      LAYER li1 ;
        RECT 62.730 69.560 63.680 70.440 ;
        RECT 63.860 69.690 64.190 70.620 ;
        RECT 64.800 70.440 65.130 71.220 ;
        RECT 65.340 70.890 65.670 71.880 ;
        RECT 66.330 71.370 67.280 72.700 ;
      LAYER li1 ;
        RECT 67.460 71.270 67.710 72.950 ;
      LAYER li1 ;
        RECT 67.890 72.870 68.840 72.950 ;
        RECT 67.890 72.700 67.920 72.870 ;
        RECT 68.090 72.700 68.280 72.870 ;
        RECT 68.450 72.700 68.640 72.870 ;
        RECT 68.810 72.700 68.840 72.870 ;
        RECT 67.890 71.450 68.840 72.700 ;
      LAYER li1 ;
        RECT 69.020 71.270 69.350 72.950 ;
      LAYER li1 ;
        RECT 69.530 72.870 70.480 72.950 ;
        RECT 69.530 72.700 69.560 72.870 ;
        RECT 69.730 72.700 69.920 72.870 ;
        RECT 70.090 72.700 70.280 72.870 ;
        RECT 70.450 72.700 70.480 72.870 ;
        RECT 69.530 71.490 70.480 72.700 ;
      LAYER li1 ;
        RECT 67.460 71.100 69.350 71.270 ;
        RECT 67.460 70.970 67.630 71.100 ;
        RECT 70.130 70.970 70.460 71.310 ;
        RECT 66.370 70.740 67.630 70.970 ;
      LAYER li1 ;
        RECT 67.810 70.790 69.840 70.920 ;
        RECT 70.660 70.790 70.910 72.950 ;
        RECT 71.290 72.920 72.740 72.950 ;
        RECT 71.290 72.750 71.540 72.920 ;
        RECT 71.710 72.750 71.900 72.920 ;
        RECT 72.070 72.750 72.340 72.920 ;
        RECT 72.510 72.750 72.740 72.920 ;
        RECT 71.290 71.880 72.740 72.750 ;
        RECT 73.050 72.870 73.640 72.950 ;
        RECT 73.050 72.700 73.080 72.870 ;
        RECT 73.250 72.700 73.440 72.870 ;
        RECT 73.610 72.700 73.640 72.870 ;
        RECT 67.810 70.750 70.910 70.790 ;
      LAYER li1 ;
        RECT 67.460 70.570 67.630 70.740 ;
      LAYER li1 ;
        RECT 69.670 70.620 70.910 70.750 ;
        RECT 64.800 70.040 66.100 70.440 ;
        RECT 64.490 69.560 66.100 70.040 ;
        RECT 66.330 69.560 67.280 70.520 ;
      LAYER li1 ;
        RECT 67.460 70.400 69.270 70.570 ;
        RECT 67.460 69.690 67.710 70.400 ;
      LAYER li1 ;
        RECT 67.890 69.560 68.840 70.220 ;
      LAYER li1 ;
        RECT 69.020 69.690 69.270 70.400 ;
      LAYER li1 ;
        RECT 69.450 69.560 70.400 70.440 ;
        RECT 70.580 69.690 70.910 70.620 ;
        RECT 71.520 70.440 71.850 71.220 ;
        RECT 72.060 70.890 72.390 71.880 ;
        RECT 73.050 71.370 73.640 72.700 ;
      LAYER li1 ;
        RECT 73.920 71.370 74.310 72.950 ;
      LAYER li1 ;
        RECT 74.650 72.920 76.100 72.950 ;
        RECT 74.650 72.750 74.900 72.920 ;
        RECT 75.070 72.750 75.260 72.920 ;
        RECT 75.430 72.750 75.700 72.920 ;
        RECT 75.870 72.750 76.100 72.920 ;
        RECT 74.650 71.880 76.100 72.750 ;
      LAYER li1 ;
        RECT 73.090 70.740 73.800 71.130 ;
      LAYER li1 ;
        RECT 71.520 70.040 72.820 70.440 ;
        RECT 71.210 69.560 72.820 70.040 ;
        RECT 73.050 69.560 73.640 70.520 ;
      LAYER li1 ;
        RECT 73.980 69.690 74.310 71.370 ;
      LAYER li1 ;
        RECT 74.880 70.440 75.210 71.220 ;
        RECT 75.420 70.890 75.750 71.880 ;
        RECT 77.060 71.290 77.310 72.950 ;
        RECT 77.490 72.870 78.740 72.950 ;
        RECT 77.660 72.700 77.850 72.870 ;
        RECT 78.020 72.700 78.210 72.870 ;
        RECT 78.380 72.700 78.570 72.870 ;
        RECT 77.490 71.470 78.740 72.700 ;
        RECT 78.920 71.290 79.090 72.950 ;
        RECT 77.060 71.120 79.090 71.290 ;
      LAYER li1 ;
        RECT 79.270 71.000 79.600 72.450 ;
        RECT 76.930 70.700 78.120 70.940 ;
        RECT 79.780 70.820 80.040 72.950 ;
      LAYER li1 ;
        RECT 80.410 72.920 81.860 72.950 ;
        RECT 80.410 72.750 80.660 72.920 ;
        RECT 80.830 72.750 81.020 72.920 ;
        RECT 81.190 72.750 81.460 72.920 ;
        RECT 81.630 72.750 81.860 72.920 ;
        RECT 80.410 71.880 81.860 72.750 ;
        RECT 82.170 72.870 83.120 72.950 ;
        RECT 82.170 72.700 82.200 72.870 ;
        RECT 82.370 72.700 82.560 72.870 ;
        RECT 82.730 72.700 82.920 72.870 ;
        RECT 83.090 72.700 83.120 72.870 ;
      LAYER li1 ;
        RECT 79.020 70.650 80.040 70.820 ;
      LAYER li1 ;
        RECT 74.880 70.040 76.180 70.440 ;
        RECT 74.570 69.560 76.180 70.040 ;
        RECT 77.130 69.560 78.840 70.520 ;
      LAYER li1 ;
        RECT 79.020 69.690 79.270 70.650 ;
      LAYER li1 ;
        RECT 79.480 69.560 80.070 70.470 ;
        RECT 80.640 70.440 80.970 71.220 ;
        RECT 81.180 70.890 81.510 71.880 ;
        RECT 82.170 71.370 83.120 72.700 ;
      LAYER li1 ;
        RECT 83.300 71.270 83.550 72.950 ;
      LAYER li1 ;
        RECT 83.730 72.870 84.680 72.950 ;
        RECT 83.730 72.700 83.760 72.870 ;
        RECT 83.930 72.700 84.120 72.870 ;
        RECT 84.290 72.700 84.480 72.870 ;
        RECT 84.650 72.700 84.680 72.870 ;
        RECT 83.730 71.450 84.680 72.700 ;
      LAYER li1 ;
        RECT 84.860 71.270 85.190 72.950 ;
      LAYER li1 ;
        RECT 85.370 72.870 86.320 72.950 ;
        RECT 85.370 72.700 85.400 72.870 ;
        RECT 85.570 72.700 85.760 72.870 ;
        RECT 85.930 72.700 86.120 72.870 ;
        RECT 86.290 72.700 86.320 72.870 ;
        RECT 85.370 71.490 86.320 72.700 ;
      LAYER li1 ;
        RECT 83.300 71.100 85.190 71.270 ;
        RECT 83.300 70.970 83.470 71.100 ;
        RECT 85.970 70.970 86.300 71.310 ;
        RECT 82.210 70.740 83.470 70.970 ;
      LAYER li1 ;
        RECT 83.650 70.790 85.680 70.920 ;
        RECT 86.500 70.790 86.750 72.950 ;
        RECT 87.130 72.920 88.580 72.950 ;
        RECT 87.130 72.750 87.380 72.920 ;
        RECT 87.550 72.750 87.740 72.920 ;
        RECT 87.910 72.750 88.180 72.920 ;
        RECT 88.350 72.750 88.580 72.920 ;
        RECT 87.130 71.880 88.580 72.750 ;
        RECT 88.890 72.870 89.840 72.950 ;
        RECT 88.890 72.700 88.920 72.870 ;
        RECT 89.090 72.700 89.280 72.870 ;
        RECT 89.450 72.700 89.640 72.870 ;
        RECT 89.810 72.700 89.840 72.870 ;
        RECT 83.650 70.750 86.750 70.790 ;
      LAYER li1 ;
        RECT 83.300 70.570 83.470 70.740 ;
      LAYER li1 ;
        RECT 85.510 70.620 86.750 70.750 ;
        RECT 80.640 70.040 81.940 70.440 ;
        RECT 80.330 69.560 81.940 70.040 ;
        RECT 82.170 69.560 83.120 70.520 ;
      LAYER li1 ;
        RECT 83.300 70.400 85.110 70.570 ;
        RECT 83.300 69.690 83.550 70.400 ;
      LAYER li1 ;
        RECT 83.730 69.560 84.680 70.220 ;
      LAYER li1 ;
        RECT 84.860 69.690 85.110 70.400 ;
      LAYER li1 ;
        RECT 85.290 69.560 86.240 70.440 ;
        RECT 86.420 69.690 86.750 70.620 ;
        RECT 87.360 70.440 87.690 71.220 ;
        RECT 87.900 70.890 88.230 71.880 ;
        RECT 88.890 71.370 89.840 72.700 ;
      LAYER li1 ;
        RECT 90.020 71.270 90.270 72.950 ;
      LAYER li1 ;
        RECT 90.450 72.870 91.400 72.950 ;
        RECT 90.450 72.700 90.480 72.870 ;
        RECT 90.650 72.700 90.840 72.870 ;
        RECT 91.010 72.700 91.200 72.870 ;
        RECT 91.370 72.700 91.400 72.870 ;
        RECT 90.450 71.450 91.400 72.700 ;
      LAYER li1 ;
        RECT 91.580 71.270 91.910 72.950 ;
      LAYER li1 ;
        RECT 92.090 72.870 93.040 72.950 ;
        RECT 92.090 72.700 92.120 72.870 ;
        RECT 92.290 72.700 92.480 72.870 ;
        RECT 92.650 72.700 92.840 72.870 ;
        RECT 93.010 72.700 93.040 72.870 ;
        RECT 92.090 71.490 93.040 72.700 ;
      LAYER li1 ;
        RECT 90.020 71.100 91.910 71.270 ;
        RECT 90.020 70.970 90.190 71.100 ;
        RECT 92.690 70.970 93.020 71.310 ;
        RECT 88.930 70.740 90.190 70.970 ;
      LAYER li1 ;
        RECT 90.370 70.790 92.400 70.920 ;
        RECT 93.220 70.790 93.470 72.950 ;
        RECT 93.850 72.920 95.300 72.950 ;
        RECT 93.850 72.750 94.100 72.920 ;
        RECT 94.270 72.750 94.460 72.920 ;
        RECT 94.630 72.750 94.900 72.920 ;
        RECT 95.070 72.750 95.300 72.920 ;
        RECT 93.850 71.880 95.300 72.750 ;
        RECT 95.610 72.870 96.200 72.950 ;
        RECT 95.610 72.700 95.640 72.870 ;
        RECT 95.810 72.700 96.000 72.870 ;
        RECT 96.170 72.700 96.200 72.870 ;
        RECT 90.370 70.750 93.470 70.790 ;
      LAYER li1 ;
        RECT 90.020 70.570 90.190 70.740 ;
      LAYER li1 ;
        RECT 92.230 70.620 93.470 70.750 ;
        RECT 87.360 70.040 88.660 70.440 ;
        RECT 87.050 69.560 88.660 70.040 ;
        RECT 88.890 69.560 89.840 70.520 ;
      LAYER li1 ;
        RECT 90.020 70.400 91.830 70.570 ;
        RECT 90.020 69.690 90.270 70.400 ;
      LAYER li1 ;
        RECT 90.450 69.560 91.400 70.220 ;
      LAYER li1 ;
        RECT 91.580 69.690 91.830 70.400 ;
      LAYER li1 ;
        RECT 92.010 69.560 92.960 70.440 ;
        RECT 93.140 69.690 93.470 70.620 ;
        RECT 94.080 70.440 94.410 71.220 ;
        RECT 94.620 70.890 94.950 71.880 ;
        RECT 95.610 71.370 96.200 72.700 ;
      LAYER li1 ;
        RECT 96.480 71.370 96.870 72.950 ;
      LAYER li1 ;
        RECT 97.210 72.920 98.660 72.950 ;
        RECT 97.210 72.750 97.460 72.920 ;
        RECT 97.630 72.750 97.820 72.920 ;
        RECT 97.990 72.750 98.260 72.920 ;
        RECT 98.430 72.750 98.660 72.920 ;
        RECT 97.210 71.880 98.660 72.750 ;
        RECT 94.080 70.040 95.380 70.440 ;
        RECT 93.770 69.560 95.380 70.040 ;
        RECT 95.610 69.560 96.200 70.520 ;
      LAYER li1 ;
        RECT 96.540 69.690 96.870 71.370 ;
      LAYER li1 ;
        RECT 97.440 70.440 97.770 71.220 ;
        RECT 97.980 70.890 98.310 71.880 ;
        RECT 99.140 71.290 99.390 72.950 ;
        RECT 99.570 72.870 100.820 72.950 ;
        RECT 99.740 72.700 99.930 72.870 ;
        RECT 100.100 72.700 100.290 72.870 ;
        RECT 100.460 72.700 100.650 72.870 ;
        RECT 99.570 71.470 100.820 72.700 ;
        RECT 101.000 71.290 101.170 72.950 ;
        RECT 99.140 71.120 101.170 71.290 ;
      LAYER li1 ;
        RECT 101.350 71.000 101.680 72.450 ;
        RECT 99.010 70.700 100.200 70.940 ;
        RECT 100.450 70.700 100.800 70.940 ;
        RECT 101.860 70.820 102.120 72.950 ;
      LAYER li1 ;
        RECT 102.490 72.920 103.940 72.950 ;
        RECT 102.490 72.750 102.740 72.920 ;
        RECT 102.910 72.750 103.100 72.920 ;
        RECT 103.270 72.750 103.540 72.920 ;
        RECT 103.710 72.750 103.940 72.920 ;
        RECT 102.490 71.880 103.940 72.750 ;
        RECT 104.250 72.870 105.200 72.950 ;
        RECT 104.250 72.700 104.280 72.870 ;
        RECT 104.450 72.700 104.640 72.870 ;
        RECT 104.810 72.700 105.000 72.870 ;
        RECT 105.170 72.700 105.200 72.870 ;
      LAYER li1 ;
        RECT 101.100 70.650 102.120 70.820 ;
      LAYER li1 ;
        RECT 97.440 70.040 98.740 70.440 ;
        RECT 97.130 69.560 98.740 70.040 ;
        RECT 99.210 69.560 100.920 70.520 ;
      LAYER li1 ;
        RECT 101.100 69.690 101.350 70.650 ;
      LAYER li1 ;
        RECT 101.560 69.560 102.150 70.470 ;
        RECT 102.720 70.440 103.050 71.220 ;
        RECT 103.260 70.890 103.590 71.880 ;
        RECT 104.250 71.370 105.200 72.700 ;
      LAYER li1 ;
        RECT 104.290 70.740 105.180 71.130 ;
        RECT 105.380 70.890 105.630 72.950 ;
      LAYER li1 ;
        RECT 105.820 72.870 106.410 72.950 ;
        RECT 105.820 72.700 105.850 72.870 ;
        RECT 106.020 72.700 106.210 72.870 ;
        RECT 106.380 72.700 106.410 72.870 ;
        RECT 105.820 71.370 106.410 72.700 ;
        RECT 106.810 72.920 108.260 72.950 ;
        RECT 106.810 72.750 107.060 72.920 ;
        RECT 107.230 72.750 107.420 72.920 ;
        RECT 107.590 72.750 107.860 72.920 ;
        RECT 108.030 72.750 108.260 72.920 ;
        RECT 106.810 71.880 108.260 72.750 ;
        RECT 108.570 72.870 110.240 72.950 ;
        RECT 108.570 72.700 108.600 72.870 ;
        RECT 108.770 72.700 108.960 72.870 ;
        RECT 109.130 72.700 109.320 72.870 ;
        RECT 109.490 72.700 109.680 72.870 ;
        RECT 109.850 72.700 110.040 72.870 ;
        RECT 110.210 72.700 110.240 72.870 ;
      LAYER li1 ;
        RECT 105.380 70.720 105.960 70.890 ;
        RECT 106.140 70.720 106.440 71.050 ;
        RECT 105.740 70.540 105.960 70.720 ;
      LAYER li1 ;
        RECT 102.720 70.040 104.020 70.440 ;
        RECT 102.410 69.560 104.020 70.040 ;
        RECT 104.250 69.560 105.560 70.540 ;
      LAYER li1 ;
        RECT 105.740 70.370 106.340 70.540 ;
        RECT 106.010 70.200 106.340 70.370 ;
      LAYER li1 ;
        RECT 107.040 70.440 107.370 71.220 ;
        RECT 107.580 70.890 107.910 71.880 ;
        RECT 108.570 71.490 110.240 72.700 ;
      LAYER li1 ;
        RECT 108.610 70.970 109.800 71.310 ;
        RECT 109.980 70.970 110.310 71.310 ;
        RECT 110.500 70.790 110.760 72.950 ;
      LAYER li1 ;
        RECT 111.130 72.920 112.580 72.950 ;
        RECT 111.130 72.750 111.380 72.920 ;
        RECT 111.550 72.750 111.740 72.920 ;
        RECT 111.910 72.750 112.180 72.920 ;
        RECT 112.350 72.750 112.580 72.920 ;
        RECT 111.130 71.880 112.580 72.750 ;
        RECT 112.890 72.870 113.480 72.950 ;
        RECT 112.890 72.700 112.920 72.870 ;
        RECT 113.090 72.700 113.280 72.870 ;
        RECT 113.450 72.700 113.480 72.870 ;
      LAYER li1 ;
        RECT 109.680 70.620 110.760 70.790 ;
        RECT 106.010 70.030 106.400 70.200 ;
      LAYER li1 ;
        RECT 107.040 70.040 108.340 70.440 ;
      LAYER li1 ;
        RECT 106.010 69.710 106.340 70.030 ;
      LAYER li1 ;
        RECT 106.730 69.560 108.340 70.040 ;
        RECT 108.570 69.560 109.500 70.520 ;
      LAYER li1 ;
        RECT 109.680 69.690 110.010 70.620 ;
      LAYER li1 ;
        RECT 111.360 70.440 111.690 71.220 ;
        RECT 111.900 70.890 112.230 71.880 ;
        RECT 112.890 71.370 113.480 72.700 ;
      LAYER li1 ;
        RECT 113.760 71.370 114.150 72.950 ;
      LAYER li1 ;
        RECT 114.490 72.920 115.940 72.950 ;
        RECT 114.490 72.750 114.740 72.920 ;
        RECT 114.910 72.750 115.100 72.920 ;
        RECT 115.270 72.750 115.540 72.920 ;
        RECT 115.710 72.750 115.940 72.920 ;
        RECT 114.490 71.880 115.940 72.750 ;
        RECT 116.250 72.870 117.200 72.950 ;
        RECT 116.250 72.700 116.280 72.870 ;
        RECT 116.450 72.700 116.640 72.870 ;
        RECT 116.810 72.700 117.000 72.870 ;
        RECT 117.170 72.700 117.200 72.870 ;
      LAYER li1 ;
        RECT 112.930 70.740 113.640 71.130 ;
      LAYER li1 ;
        RECT 110.200 69.560 110.790 70.440 ;
        RECT 111.360 70.040 112.660 70.440 ;
        RECT 111.050 69.560 112.660 70.040 ;
        RECT 112.890 69.560 113.480 70.520 ;
      LAYER li1 ;
        RECT 113.820 69.690 114.150 71.370 ;
      LAYER li1 ;
        RECT 114.720 70.440 115.050 71.220 ;
        RECT 115.260 70.890 115.590 71.880 ;
        RECT 116.250 71.370 117.200 72.700 ;
      LAYER li1 ;
        RECT 117.380 71.270 117.630 72.950 ;
      LAYER li1 ;
        RECT 117.810 72.870 118.760 72.950 ;
        RECT 117.810 72.700 117.840 72.870 ;
        RECT 118.010 72.700 118.200 72.870 ;
        RECT 118.370 72.700 118.560 72.870 ;
        RECT 118.730 72.700 118.760 72.870 ;
        RECT 117.810 71.450 118.760 72.700 ;
      LAYER li1 ;
        RECT 118.940 71.270 119.270 72.950 ;
      LAYER li1 ;
        RECT 119.450 72.870 120.400 72.950 ;
        RECT 119.450 72.700 119.480 72.870 ;
        RECT 119.650 72.700 119.840 72.870 ;
        RECT 120.010 72.700 120.200 72.870 ;
        RECT 120.370 72.700 120.400 72.870 ;
        RECT 119.450 71.490 120.400 72.700 ;
      LAYER li1 ;
        RECT 117.380 71.100 119.270 71.270 ;
        RECT 117.380 70.970 117.550 71.100 ;
        RECT 120.050 70.970 120.380 71.310 ;
        RECT 116.290 70.740 117.550 70.970 ;
      LAYER li1 ;
        RECT 117.730 70.790 119.760 70.920 ;
        RECT 120.580 70.790 120.830 72.950 ;
        RECT 121.210 72.920 122.660 72.950 ;
        RECT 121.210 72.750 121.460 72.920 ;
        RECT 121.630 72.750 121.820 72.920 ;
        RECT 121.990 72.750 122.260 72.920 ;
        RECT 122.430 72.750 122.660 72.920 ;
        RECT 121.210 71.880 122.660 72.750 ;
        RECT 117.730 70.750 120.830 70.790 ;
      LAYER li1 ;
        RECT 117.380 70.570 117.550 70.740 ;
      LAYER li1 ;
        RECT 119.590 70.620 120.830 70.750 ;
        RECT 114.720 70.040 116.020 70.440 ;
        RECT 114.410 69.560 116.020 70.040 ;
        RECT 116.250 69.560 117.200 70.520 ;
      LAYER li1 ;
        RECT 117.380 70.400 119.190 70.570 ;
        RECT 117.380 69.690 117.630 70.400 ;
      LAYER li1 ;
        RECT 117.810 69.560 118.760 70.220 ;
      LAYER li1 ;
        RECT 118.940 69.690 119.190 70.400 ;
      LAYER li1 ;
        RECT 119.370 69.560 120.320 70.440 ;
        RECT 120.500 69.690 120.830 70.620 ;
        RECT 121.440 70.440 121.770 71.220 ;
        RECT 121.980 70.890 122.310 71.880 ;
      LAYER li1 ;
        RECT 123.000 71.370 123.430 72.950 ;
      LAYER li1 ;
        RECT 123.610 72.870 124.170 72.950 ;
        RECT 123.610 72.700 123.620 72.870 ;
        RECT 123.790 72.700 123.980 72.870 ;
        RECT 124.150 72.700 124.170 72.870 ;
        RECT 123.610 71.370 124.170 72.700 ;
        RECT 125.780 72.920 128.520 72.940 ;
        RECT 125.780 72.750 125.990 72.920 ;
        RECT 126.160 72.750 126.430 72.920 ;
        RECT 126.600 72.750 126.840 72.920 ;
        RECT 127.010 72.750 127.270 72.920 ;
        RECT 127.440 72.750 127.710 72.920 ;
        RECT 127.880 72.750 128.120 72.920 ;
        RECT 128.290 72.750 128.520 72.920 ;
        RECT 121.440 70.040 122.740 70.440 ;
        RECT 121.130 69.560 122.740 70.040 ;
      LAYER li1 ;
        RECT 123.000 69.690 123.250 71.370 ;
      LAYER li1 ;
        RECT 123.560 70.480 123.890 70.940 ;
      LAYER li1 ;
        RECT 124.350 70.660 124.680 72.450 ;
      LAYER li1 ;
        RECT 124.860 70.480 125.110 72.200 ;
        RECT 125.780 71.870 128.520 72.750 ;
        RECT 126.020 70.550 126.350 71.220 ;
        RECT 126.750 70.890 127.080 71.870 ;
        RECT 127.300 70.550 127.630 71.220 ;
        RECT 128.030 70.890 128.360 71.870 ;
      LAYER li1 ;
        RECT 129.240 71.370 129.670 72.950 ;
      LAYER li1 ;
        RECT 129.850 72.870 130.410 72.950 ;
        RECT 129.850 72.700 129.860 72.870 ;
        RECT 130.030 72.700 130.220 72.870 ;
        RECT 130.390 72.700 130.410 72.870 ;
        RECT 129.850 71.370 130.410 72.700 ;
        RECT 132.020 72.920 134.760 72.940 ;
        RECT 132.020 72.750 132.230 72.920 ;
        RECT 132.400 72.750 132.670 72.920 ;
        RECT 132.840 72.750 133.080 72.920 ;
        RECT 133.250 72.750 133.510 72.920 ;
        RECT 133.680 72.750 133.950 72.920 ;
        RECT 134.120 72.750 134.360 72.920 ;
        RECT 134.530 72.750 134.760 72.920 ;
        RECT 123.560 70.310 125.110 70.480 ;
        RECT 123.430 69.560 124.680 70.130 ;
        RECT 124.860 69.690 125.110 70.310 ;
        RECT 125.860 69.550 128.590 70.550 ;
      LAYER li1 ;
        RECT 129.240 69.690 129.490 71.370 ;
      LAYER li1 ;
        RECT 129.800 70.480 130.130 70.940 ;
      LAYER li1 ;
        RECT 130.590 70.660 130.920 72.450 ;
      LAYER li1 ;
        RECT 131.100 70.480 131.350 72.200 ;
        RECT 132.020 71.870 134.760 72.750 ;
        RECT 135.860 72.920 138.600 72.940 ;
        RECT 135.860 72.750 136.070 72.920 ;
        RECT 136.240 72.750 136.510 72.920 ;
        RECT 136.680 72.750 136.920 72.920 ;
        RECT 137.090 72.750 137.350 72.920 ;
        RECT 137.520 72.750 137.790 72.920 ;
        RECT 137.960 72.750 138.200 72.920 ;
        RECT 138.370 72.750 138.600 72.920 ;
        RECT 135.860 71.870 138.600 72.750 ;
        RECT 139.450 72.920 140.900 72.950 ;
        RECT 139.450 72.750 139.700 72.920 ;
        RECT 139.870 72.750 140.060 72.920 ;
        RECT 140.230 72.750 140.500 72.920 ;
        RECT 140.670 72.750 140.900 72.920 ;
        RECT 139.450 71.880 140.900 72.750 ;
        RECT 132.260 70.550 132.590 71.220 ;
        RECT 132.990 70.890 133.320 71.870 ;
        RECT 133.540 70.550 133.870 71.220 ;
        RECT 134.270 70.890 134.600 71.870 ;
        RECT 136.100 70.550 136.430 71.220 ;
        RECT 136.830 70.890 137.160 71.870 ;
        RECT 137.380 70.550 137.710 71.220 ;
        RECT 138.110 70.890 138.440 71.870 ;
        RECT 129.800 70.310 131.350 70.480 ;
        RECT 129.670 69.560 130.920 70.130 ;
        RECT 131.100 69.690 131.350 70.310 ;
        RECT 132.100 69.550 134.830 70.550 ;
        RECT 135.940 69.550 138.670 70.550 ;
        RECT 139.680 70.440 140.010 71.220 ;
        RECT 140.220 70.890 140.550 71.880 ;
        RECT 139.680 70.040 140.980 70.440 ;
        RECT 139.370 69.560 140.980 70.040 ;
        RECT 5.760 69.100 5.920 69.280 ;
        RECT 6.090 69.100 6.400 69.280 ;
        RECT 6.570 69.100 6.880 69.280 ;
        RECT 7.050 69.100 7.360 69.280 ;
        RECT 7.530 69.100 7.840 69.280 ;
        RECT 8.010 69.100 8.320 69.280 ;
        RECT 8.490 69.100 8.800 69.280 ;
        RECT 8.970 69.100 9.280 69.280 ;
        RECT 9.450 69.100 9.760 69.280 ;
        RECT 9.930 69.100 10.240 69.280 ;
        RECT 10.410 69.100 10.720 69.280 ;
        RECT 10.890 69.100 11.200 69.280 ;
        RECT 11.370 69.100 11.680 69.280 ;
        RECT 11.850 69.100 12.160 69.280 ;
        RECT 12.330 69.100 12.640 69.280 ;
        RECT 12.810 69.100 13.120 69.280 ;
        RECT 13.290 69.100 13.600 69.280 ;
        RECT 13.770 69.100 14.080 69.280 ;
        RECT 14.250 69.100 14.560 69.280 ;
        RECT 14.730 69.100 15.040 69.280 ;
        RECT 15.210 69.100 15.520 69.280 ;
        RECT 15.690 69.100 16.000 69.280 ;
        RECT 16.170 69.100 16.480 69.280 ;
        RECT 16.650 69.100 16.960 69.280 ;
        RECT 17.130 69.100 17.440 69.280 ;
        RECT 17.610 69.100 17.920 69.280 ;
        RECT 18.090 69.100 18.400 69.280 ;
        RECT 18.570 69.100 18.880 69.280 ;
        RECT 19.050 69.100 19.360 69.280 ;
        RECT 19.530 69.100 19.840 69.280 ;
        RECT 20.010 69.100 20.320 69.280 ;
        RECT 20.490 69.100 20.800 69.280 ;
        RECT 20.970 69.100 21.280 69.280 ;
        RECT 21.450 69.100 21.760 69.280 ;
        RECT 21.930 69.100 22.240 69.280 ;
        RECT 22.410 69.100 22.720 69.280 ;
        RECT 22.890 69.100 23.200 69.280 ;
        RECT 23.370 69.100 23.680 69.280 ;
        RECT 23.850 69.100 24.160 69.280 ;
        RECT 24.330 69.100 24.640 69.280 ;
        RECT 24.810 69.100 25.120 69.280 ;
        RECT 25.290 69.100 25.600 69.280 ;
        RECT 25.770 69.100 26.080 69.280 ;
        RECT 26.250 69.100 26.560 69.280 ;
        RECT 26.730 69.100 27.040 69.280 ;
        RECT 27.210 69.100 27.520 69.280 ;
        RECT 27.690 69.100 28.000 69.280 ;
        RECT 28.170 69.100 28.480 69.280 ;
        RECT 28.650 69.100 28.960 69.280 ;
        RECT 29.130 69.100 29.440 69.280 ;
        RECT 29.610 69.100 29.920 69.280 ;
        RECT 30.090 69.100 30.400 69.280 ;
        RECT 30.570 69.100 30.880 69.280 ;
        RECT 31.050 69.100 31.360 69.280 ;
        RECT 31.530 69.100 31.840 69.280 ;
        RECT 32.010 69.100 32.320 69.280 ;
        RECT 32.490 69.100 32.800 69.280 ;
        RECT 32.970 69.100 33.280 69.280 ;
        RECT 33.450 69.100 33.760 69.280 ;
        RECT 33.930 69.100 34.240 69.280 ;
        RECT 34.410 69.100 34.720 69.280 ;
        RECT 34.890 69.100 35.200 69.280 ;
        RECT 35.370 69.100 35.680 69.280 ;
        RECT 35.850 69.100 36.160 69.280 ;
        RECT 36.330 69.100 36.640 69.280 ;
        RECT 36.810 69.100 37.120 69.280 ;
        RECT 37.290 69.100 37.600 69.280 ;
        RECT 37.770 69.100 38.080 69.280 ;
        RECT 38.250 69.100 38.560 69.280 ;
        RECT 38.730 69.100 39.040 69.280 ;
        RECT 39.210 69.100 39.520 69.280 ;
        RECT 39.690 69.100 40.000 69.280 ;
        RECT 40.170 69.100 40.480 69.280 ;
        RECT 40.650 69.100 40.960 69.280 ;
        RECT 41.130 69.100 41.440 69.280 ;
        RECT 41.610 69.100 41.920 69.280 ;
        RECT 42.090 69.100 42.400 69.280 ;
        RECT 42.570 69.100 42.880 69.280 ;
        RECT 43.050 69.100 43.360 69.280 ;
        RECT 43.530 69.100 43.840 69.280 ;
        RECT 44.010 69.100 44.320 69.280 ;
        RECT 44.490 69.100 44.800 69.280 ;
        RECT 44.970 69.100 45.280 69.280 ;
        RECT 45.450 69.100 45.760 69.280 ;
        RECT 45.930 69.100 46.240 69.280 ;
        RECT 46.410 69.100 46.720 69.280 ;
        RECT 46.890 69.100 47.200 69.280 ;
        RECT 47.370 69.100 47.520 69.280 ;
        RECT 48.000 69.100 48.160 69.280 ;
        RECT 48.330 69.100 48.640 69.280 ;
        RECT 48.810 69.100 49.120 69.280 ;
        RECT 49.290 69.100 49.600 69.280 ;
        RECT 49.770 69.100 50.080 69.280 ;
        RECT 50.250 69.100 50.560 69.280 ;
        RECT 50.730 69.100 51.040 69.280 ;
        RECT 51.210 69.100 51.520 69.280 ;
        RECT 51.690 69.100 52.000 69.280 ;
        RECT 52.170 69.100 52.480 69.280 ;
        RECT 52.650 69.100 52.960 69.280 ;
        RECT 53.130 69.100 53.440 69.280 ;
        RECT 53.610 69.100 53.920 69.280 ;
        RECT 54.090 69.100 54.400 69.280 ;
        RECT 54.570 69.100 54.880 69.280 ;
        RECT 55.050 69.100 55.360 69.280 ;
        RECT 55.530 69.100 55.840 69.280 ;
        RECT 56.010 69.100 56.320 69.280 ;
        RECT 56.490 69.100 56.800 69.280 ;
        RECT 56.970 69.100 57.280 69.280 ;
        RECT 57.450 69.100 57.760 69.280 ;
        RECT 57.930 69.100 58.240 69.280 ;
        RECT 58.410 69.100 58.720 69.280 ;
        RECT 58.890 69.100 59.040 69.280 ;
        RECT 59.520 69.100 59.680 69.280 ;
        RECT 59.850 69.100 60.160 69.280 ;
        RECT 60.330 69.100 60.640 69.280 ;
        RECT 60.810 69.100 61.120 69.280 ;
        RECT 61.290 69.100 61.600 69.280 ;
        RECT 61.770 69.100 62.080 69.280 ;
        RECT 62.250 69.100 62.560 69.280 ;
        RECT 62.730 69.100 63.040 69.280 ;
        RECT 63.210 69.100 63.520 69.280 ;
        RECT 63.690 69.100 64.000 69.280 ;
        RECT 64.170 69.100 64.480 69.280 ;
        RECT 64.650 69.100 64.960 69.280 ;
        RECT 65.130 69.100 65.440 69.280 ;
        RECT 65.610 69.100 65.920 69.280 ;
        RECT 66.090 69.100 66.400 69.280 ;
        RECT 66.570 69.100 66.880 69.280 ;
        RECT 67.050 69.100 67.360 69.280 ;
        RECT 67.530 69.100 67.840 69.280 ;
        RECT 68.010 69.100 68.320 69.280 ;
        RECT 68.490 69.100 68.800 69.280 ;
        RECT 68.970 69.100 69.280 69.280 ;
        RECT 69.450 69.100 69.760 69.280 ;
        RECT 69.930 69.100 70.240 69.280 ;
        RECT 70.410 69.100 70.720 69.280 ;
        RECT 70.890 69.100 71.200 69.280 ;
        RECT 71.370 69.100 71.680 69.280 ;
        RECT 71.850 69.100 72.160 69.280 ;
        RECT 72.330 69.100 72.640 69.280 ;
        RECT 72.810 69.100 73.120 69.280 ;
        RECT 73.290 69.100 73.600 69.280 ;
        RECT 73.770 69.100 74.080 69.280 ;
        RECT 74.250 69.100 74.560 69.280 ;
        RECT 74.730 69.100 75.040 69.280 ;
        RECT 75.210 69.100 75.520 69.280 ;
        RECT 75.690 69.100 76.000 69.280 ;
        RECT 76.170 69.100 76.320 69.280 ;
        RECT 76.800 69.100 76.960 69.280 ;
        RECT 77.130 69.100 77.440 69.280 ;
        RECT 77.610 69.100 77.920 69.280 ;
        RECT 78.090 69.100 78.400 69.280 ;
        RECT 78.570 69.100 78.880 69.280 ;
        RECT 79.050 69.100 79.360 69.280 ;
        RECT 79.530 69.100 79.840 69.280 ;
        RECT 80.010 69.100 80.320 69.280 ;
        RECT 80.490 69.100 80.800 69.280 ;
        RECT 80.970 69.100 81.280 69.280 ;
        RECT 81.450 69.100 81.760 69.280 ;
        RECT 81.930 69.100 82.240 69.280 ;
        RECT 82.410 69.100 82.720 69.280 ;
        RECT 82.890 69.100 83.200 69.280 ;
        RECT 83.370 69.100 83.680 69.280 ;
        RECT 83.850 69.100 84.160 69.280 ;
        RECT 84.330 69.100 84.640 69.280 ;
        RECT 84.810 69.100 85.120 69.280 ;
        RECT 85.290 69.100 85.600 69.280 ;
        RECT 85.770 69.100 86.080 69.280 ;
        RECT 86.250 69.100 86.560 69.280 ;
        RECT 86.730 69.100 87.040 69.280 ;
        RECT 87.210 69.100 87.520 69.280 ;
        RECT 87.690 69.100 88.000 69.280 ;
        RECT 88.170 69.100 88.480 69.280 ;
        RECT 88.650 69.100 88.960 69.280 ;
        RECT 89.130 69.100 89.440 69.280 ;
        RECT 89.610 69.100 89.920 69.280 ;
        RECT 90.090 69.100 90.400 69.280 ;
        RECT 90.570 69.100 90.880 69.280 ;
        RECT 91.050 69.100 91.360 69.280 ;
        RECT 91.530 69.100 91.840 69.280 ;
        RECT 92.010 69.100 92.320 69.280 ;
        RECT 92.490 69.100 92.800 69.280 ;
        RECT 92.970 69.100 93.280 69.280 ;
        RECT 93.450 69.100 93.760 69.280 ;
        RECT 93.930 69.100 94.240 69.280 ;
        RECT 94.410 69.100 94.720 69.280 ;
        RECT 94.890 69.100 95.200 69.280 ;
        RECT 95.370 69.100 95.680 69.280 ;
        RECT 95.850 69.100 96.160 69.280 ;
        RECT 96.330 69.100 96.640 69.280 ;
        RECT 96.810 69.100 97.120 69.280 ;
        RECT 97.290 69.100 97.600 69.280 ;
        RECT 97.770 69.100 98.080 69.280 ;
        RECT 98.250 69.100 98.560 69.280 ;
        RECT 98.730 69.100 99.040 69.280 ;
        RECT 99.210 69.100 99.520 69.280 ;
        RECT 99.690 69.100 100.000 69.280 ;
        RECT 100.170 69.100 100.480 69.280 ;
        RECT 100.650 69.100 100.960 69.280 ;
        RECT 101.130 69.100 101.440 69.280 ;
        RECT 101.610 69.100 101.920 69.280 ;
        RECT 102.090 69.100 102.400 69.280 ;
        RECT 102.570 69.100 102.880 69.280 ;
        RECT 103.050 69.100 103.360 69.280 ;
        RECT 103.530 69.100 103.840 69.280 ;
        RECT 104.010 69.100 104.320 69.280 ;
        RECT 104.490 69.100 104.800 69.280 ;
        RECT 104.970 69.100 105.280 69.280 ;
        RECT 105.450 69.100 105.760 69.280 ;
        RECT 105.930 69.100 106.240 69.280 ;
        RECT 106.410 69.100 106.720 69.280 ;
        RECT 106.890 69.100 107.200 69.280 ;
        RECT 107.370 69.100 107.680 69.280 ;
        RECT 107.850 69.100 108.160 69.280 ;
        RECT 108.330 69.100 108.640 69.280 ;
        RECT 108.810 69.100 109.120 69.280 ;
        RECT 109.290 69.100 109.600 69.280 ;
        RECT 109.770 69.100 110.080 69.280 ;
        RECT 110.250 69.100 110.560 69.280 ;
        RECT 110.730 69.100 111.040 69.280 ;
        RECT 111.210 69.100 111.520 69.280 ;
        RECT 111.690 69.100 112.000 69.280 ;
        RECT 112.170 69.100 112.480 69.280 ;
        RECT 112.650 69.100 112.960 69.280 ;
        RECT 113.130 69.100 113.440 69.280 ;
        RECT 113.610 69.100 113.920 69.280 ;
        RECT 114.090 69.100 114.400 69.280 ;
        RECT 114.570 69.100 114.880 69.280 ;
        RECT 115.050 69.100 115.360 69.280 ;
        RECT 115.530 69.100 115.840 69.280 ;
        RECT 116.010 69.100 116.320 69.280 ;
        RECT 116.490 69.100 116.800 69.280 ;
        RECT 116.970 69.100 117.280 69.280 ;
        RECT 117.450 69.100 117.760 69.280 ;
        RECT 117.930 69.100 118.240 69.280 ;
        RECT 118.410 69.100 118.720 69.280 ;
        RECT 118.890 69.100 119.200 69.280 ;
        RECT 119.370 69.100 119.680 69.280 ;
        RECT 119.850 69.100 120.160 69.280 ;
        RECT 120.330 69.100 120.640 69.280 ;
        RECT 120.810 69.100 121.120 69.280 ;
        RECT 121.290 69.100 121.600 69.280 ;
        RECT 121.770 69.100 122.080 69.280 ;
        RECT 122.250 69.100 122.560 69.280 ;
        RECT 122.730 69.100 123.040 69.280 ;
        RECT 123.210 69.100 123.520 69.280 ;
        RECT 123.690 69.100 124.000 69.280 ;
        RECT 124.170 69.100 124.480 69.280 ;
        RECT 124.650 69.100 124.960 69.280 ;
        RECT 125.130 69.100 125.440 69.280 ;
        RECT 125.610 69.100 125.920 69.280 ;
        RECT 126.090 69.100 126.400 69.280 ;
        RECT 126.570 69.100 126.880 69.280 ;
        RECT 127.050 69.100 127.360 69.280 ;
        RECT 127.530 69.100 127.840 69.280 ;
        RECT 128.010 69.100 128.320 69.280 ;
        RECT 128.490 69.100 128.800 69.280 ;
        RECT 128.970 69.100 129.280 69.280 ;
        RECT 129.450 69.100 129.760 69.280 ;
        RECT 129.930 69.100 130.240 69.280 ;
        RECT 130.410 69.100 130.720 69.280 ;
        RECT 130.890 69.100 131.200 69.280 ;
        RECT 131.370 69.100 131.680 69.280 ;
        RECT 131.850 69.100 132.160 69.280 ;
        RECT 132.330 69.100 132.640 69.280 ;
        RECT 132.810 69.100 133.120 69.280 ;
        RECT 133.290 69.100 133.600 69.280 ;
        RECT 133.770 69.100 134.080 69.280 ;
        RECT 134.250 69.100 134.560 69.280 ;
        RECT 134.730 69.100 135.040 69.280 ;
        RECT 135.210 69.100 135.520 69.280 ;
        RECT 135.690 69.100 136.000 69.280 ;
        RECT 136.170 69.100 136.480 69.280 ;
        RECT 136.650 69.100 136.960 69.280 ;
        RECT 137.130 69.100 137.440 69.280 ;
        RECT 137.610 69.100 137.920 69.280 ;
        RECT 138.090 69.100 138.400 69.280 ;
        RECT 138.570 69.100 138.880 69.280 ;
        RECT 139.050 69.100 139.360 69.280 ;
        RECT 139.530 69.100 139.840 69.280 ;
        RECT 140.010 69.100 140.320 69.280 ;
        RECT 140.490 69.100 140.800 69.280 ;
        RECT 140.970 69.100 141.280 69.280 ;
        RECT 141.450 69.100 141.760 69.280 ;
        RECT 141.930 69.100 142.080 69.280 ;
        RECT 5.930 68.790 7.540 68.820 ;
        RECT 9.670 68.790 10.920 68.820 ;
        RECT 11.690 68.790 13.300 68.820 ;
        RECT 5.930 68.620 5.980 68.790 ;
        RECT 6.150 68.620 6.420 68.790 ;
        RECT 6.590 68.620 6.860 68.790 ;
        RECT 7.030 68.620 7.270 68.790 ;
        RECT 7.440 68.620 7.540 68.790 ;
        RECT 5.930 68.340 7.540 68.620 ;
        RECT 6.240 67.940 7.540 68.340 ;
        RECT 6.240 67.160 6.570 67.940 ;
        RECT 6.780 66.500 7.110 67.490 ;
      LAYER li1 ;
        RECT 9.240 67.010 9.490 68.690 ;
      LAYER li1 ;
        RECT 9.840 68.620 10.030 68.790 ;
        RECT 10.200 68.620 10.390 68.790 ;
        RECT 10.560 68.620 10.750 68.790 ;
        RECT 9.670 68.250 10.920 68.620 ;
        RECT 11.100 68.070 11.350 68.690 ;
        RECT 11.690 68.620 11.740 68.790 ;
        RECT 11.910 68.620 12.180 68.790 ;
        RECT 12.350 68.620 12.620 68.790 ;
        RECT 12.790 68.620 13.030 68.790 ;
        RECT 13.200 68.620 13.300 68.790 ;
        RECT 11.690 68.340 13.300 68.620 ;
        RECT 9.800 67.900 11.350 68.070 ;
        RECT 9.800 67.440 10.130 67.900 ;
        RECT 6.010 65.630 7.460 66.500 ;
        RECT 6.010 65.460 6.260 65.630 ;
        RECT 6.430 65.460 6.620 65.630 ;
        RECT 6.790 65.460 7.060 65.630 ;
        RECT 7.230 65.460 7.460 65.630 ;
        RECT 6.010 65.430 7.460 65.460 ;
      LAYER li1 ;
        RECT 9.240 65.430 9.670 67.010 ;
      LAYER li1 ;
        RECT 9.850 65.680 10.410 67.010 ;
      LAYER li1 ;
        RECT 10.590 65.930 10.920 67.720 ;
      LAYER li1 ;
        RECT 11.100 66.180 11.350 67.900 ;
        RECT 12.000 67.940 13.300 68.340 ;
        RECT 13.530 68.790 14.460 68.820 ;
        RECT 13.530 68.620 13.550 68.790 ;
        RECT 13.720 68.620 13.910 68.790 ;
        RECT 14.080 68.620 14.270 68.790 ;
        RECT 14.440 68.620 14.460 68.790 ;
        RECT 15.160 68.790 15.750 68.820 ;
        RECT 12.000 67.160 12.330 67.940 ;
        RECT 13.530 67.860 14.460 68.620 ;
      LAYER li1 ;
        RECT 14.640 67.760 14.970 68.690 ;
      LAYER li1 ;
        RECT 15.160 68.620 15.190 68.790 ;
        RECT 15.360 68.620 15.550 68.790 ;
        RECT 15.720 68.620 15.750 68.790 ;
        RECT 15.160 67.940 15.750 68.620 ;
        RECT 16.010 68.790 17.620 68.820 ;
        RECT 16.010 68.620 16.060 68.790 ;
        RECT 16.230 68.620 16.500 68.790 ;
        RECT 16.670 68.620 16.940 68.790 ;
        RECT 17.110 68.620 17.350 68.790 ;
        RECT 17.520 68.620 17.620 68.790 ;
        RECT 16.010 68.340 17.620 68.620 ;
        RECT 16.320 67.940 17.620 68.340 ;
        RECT 17.850 68.790 19.160 68.820 ;
        RECT 17.850 68.620 17.880 68.790 ;
        RECT 18.050 68.620 18.240 68.790 ;
        RECT 18.410 68.620 18.600 68.790 ;
        RECT 18.770 68.620 18.960 68.790 ;
        RECT 19.130 68.620 19.160 68.790 ;
        RECT 20.330 68.790 21.940 68.820 ;
      LAYER li1 ;
        RECT 14.640 67.590 15.720 67.760 ;
      LAYER li1 ;
        RECT 12.540 66.500 12.870 67.490 ;
      LAYER li1 ;
        RECT 13.570 67.070 14.760 67.410 ;
        RECT 14.940 67.070 15.270 67.410 ;
      LAYER li1 ;
        RECT 9.850 65.510 9.860 65.680 ;
        RECT 10.030 65.510 10.220 65.680 ;
        RECT 10.390 65.510 10.410 65.680 ;
        RECT 9.850 65.430 10.410 65.510 ;
        RECT 11.770 65.630 13.220 66.500 ;
        RECT 11.770 65.460 12.020 65.630 ;
        RECT 12.190 65.460 12.380 65.630 ;
        RECT 12.550 65.460 12.820 65.630 ;
        RECT 12.990 65.460 13.220 65.630 ;
        RECT 11.770 65.430 13.220 65.460 ;
        RECT 13.530 65.680 15.200 66.890 ;
        RECT 13.530 65.510 13.560 65.680 ;
        RECT 13.730 65.510 13.920 65.680 ;
        RECT 14.090 65.510 14.280 65.680 ;
        RECT 14.450 65.510 14.640 65.680 ;
        RECT 14.810 65.510 15.000 65.680 ;
        RECT 15.170 65.510 15.200 65.680 ;
        RECT 13.530 65.430 15.200 65.510 ;
      LAYER li1 ;
        RECT 15.460 65.430 15.720 67.590 ;
      LAYER li1 ;
        RECT 16.320 67.160 16.650 67.940 ;
        RECT 17.850 67.840 19.160 68.620 ;
      LAYER li1 ;
        RECT 19.610 68.350 19.940 68.670 ;
      LAYER li1 ;
        RECT 20.330 68.620 20.380 68.790 ;
        RECT 20.550 68.620 20.820 68.790 ;
        RECT 20.990 68.620 21.260 68.790 ;
        RECT 21.430 68.620 21.670 68.790 ;
        RECT 21.840 68.620 21.940 68.790 ;
      LAYER li1 ;
        RECT 19.610 68.180 20.000 68.350 ;
      LAYER li1 ;
        RECT 20.330 68.340 21.940 68.620 ;
      LAYER li1 ;
        RECT 19.610 68.010 19.940 68.180 ;
        RECT 19.340 67.840 19.940 68.010 ;
      LAYER li1 ;
        RECT 20.640 67.940 21.940 68.340 ;
        RECT 22.170 68.790 23.120 68.820 ;
        RECT 22.170 68.620 22.200 68.790 ;
        RECT 22.370 68.620 22.560 68.790 ;
        RECT 22.730 68.620 22.920 68.790 ;
        RECT 23.090 68.620 23.120 68.790 ;
        RECT 23.730 68.790 24.680 68.820 ;
      LAYER li1 ;
        RECT 19.340 67.660 19.560 67.840 ;
      LAYER li1 ;
        RECT 16.860 66.500 17.190 67.490 ;
      LAYER li1 ;
        RECT 17.890 67.250 18.780 67.640 ;
        RECT 18.980 67.490 19.560 67.660 ;
      LAYER li1 ;
        RECT 16.090 65.630 17.540 66.500 ;
        RECT 16.090 65.460 16.340 65.630 ;
        RECT 16.510 65.460 16.700 65.630 ;
        RECT 16.870 65.460 17.140 65.630 ;
        RECT 17.310 65.460 17.540 65.630 ;
        RECT 16.090 65.430 17.540 65.460 ;
        RECT 17.850 65.680 18.800 67.010 ;
        RECT 17.850 65.510 17.880 65.680 ;
        RECT 18.050 65.510 18.240 65.680 ;
        RECT 18.410 65.510 18.600 65.680 ;
        RECT 18.770 65.510 18.800 65.680 ;
        RECT 17.850 65.430 18.800 65.510 ;
      LAYER li1 ;
        RECT 18.980 65.430 19.230 67.490 ;
        RECT 19.740 67.330 20.040 67.660 ;
      LAYER li1 ;
        RECT 20.640 67.160 20.970 67.940 ;
        RECT 22.170 67.860 23.120 68.620 ;
      LAYER li1 ;
        RECT 23.300 67.980 23.550 68.690 ;
      LAYER li1 ;
        RECT 23.730 68.620 23.760 68.790 ;
        RECT 23.930 68.620 24.120 68.790 ;
        RECT 24.290 68.620 24.480 68.790 ;
        RECT 24.650 68.620 24.680 68.790 ;
        RECT 25.290 68.790 26.240 68.820 ;
        RECT 23.730 68.160 24.680 68.620 ;
      LAYER li1 ;
        RECT 24.860 67.980 25.110 68.690 ;
        RECT 23.300 67.810 25.110 67.980 ;
      LAYER li1 ;
        RECT 25.290 68.620 25.320 68.790 ;
        RECT 25.490 68.620 25.680 68.790 ;
        RECT 25.850 68.620 26.040 68.790 ;
        RECT 26.210 68.620 26.240 68.790 ;
        RECT 27.050 68.790 28.660 68.820 ;
        RECT 25.290 67.940 26.240 68.620 ;
      LAYER li1 ;
        RECT 23.300 67.640 23.470 67.810 ;
      LAYER li1 ;
        RECT 26.420 67.760 26.750 68.690 ;
        RECT 27.050 68.620 27.100 68.790 ;
        RECT 27.270 68.620 27.540 68.790 ;
        RECT 27.710 68.620 27.980 68.790 ;
        RECT 28.150 68.620 28.390 68.790 ;
        RECT 28.560 68.620 28.660 68.790 ;
        RECT 27.050 68.340 28.660 68.620 ;
        RECT 19.420 65.680 20.010 67.010 ;
        RECT 21.180 66.500 21.510 67.490 ;
      LAYER li1 ;
        RECT 22.210 67.410 23.470 67.640 ;
      LAYER li1 ;
        RECT 25.510 67.630 26.750 67.760 ;
        RECT 23.650 67.590 26.750 67.630 ;
        RECT 23.650 67.460 25.680 67.590 ;
      LAYER li1 ;
        RECT 23.300 67.280 23.470 67.410 ;
        RECT 23.300 67.110 25.190 67.280 ;
      LAYER li1 ;
        RECT 19.420 65.510 19.450 65.680 ;
        RECT 19.620 65.510 19.810 65.680 ;
        RECT 19.980 65.510 20.010 65.680 ;
        RECT 19.420 65.430 20.010 65.510 ;
        RECT 20.410 65.630 21.860 66.500 ;
        RECT 20.410 65.460 20.660 65.630 ;
        RECT 20.830 65.460 21.020 65.630 ;
        RECT 21.190 65.460 21.460 65.630 ;
        RECT 21.630 65.460 21.860 65.630 ;
        RECT 20.410 65.430 21.860 65.460 ;
        RECT 22.170 65.680 23.120 67.010 ;
        RECT 22.170 65.510 22.200 65.680 ;
        RECT 22.370 65.510 22.560 65.680 ;
        RECT 22.730 65.510 22.920 65.680 ;
        RECT 23.090 65.510 23.120 65.680 ;
        RECT 22.170 65.430 23.120 65.510 ;
      LAYER li1 ;
        RECT 23.300 65.430 23.550 67.110 ;
      LAYER li1 ;
        RECT 23.730 65.680 24.680 66.930 ;
        RECT 23.730 65.510 23.760 65.680 ;
        RECT 23.930 65.510 24.120 65.680 ;
        RECT 24.290 65.510 24.480 65.680 ;
        RECT 24.650 65.510 24.680 65.680 ;
        RECT 23.730 65.430 24.680 65.510 ;
      LAYER li1 ;
        RECT 24.860 65.430 25.190 67.110 ;
        RECT 25.970 67.070 26.300 67.410 ;
      LAYER li1 ;
        RECT 25.370 65.680 26.320 66.890 ;
        RECT 25.370 65.510 25.400 65.680 ;
        RECT 25.570 65.510 25.760 65.680 ;
        RECT 25.930 65.510 26.120 65.680 ;
        RECT 26.290 65.510 26.320 65.680 ;
        RECT 25.370 65.430 26.320 65.510 ;
        RECT 26.500 65.430 26.750 67.590 ;
        RECT 27.360 67.940 28.660 68.340 ;
        RECT 28.890 68.790 29.840 68.820 ;
        RECT 28.890 68.620 28.920 68.790 ;
        RECT 29.090 68.620 29.280 68.790 ;
        RECT 29.450 68.620 29.640 68.790 ;
        RECT 29.810 68.620 29.840 68.790 ;
        RECT 30.450 68.790 31.400 68.820 ;
        RECT 27.360 67.160 27.690 67.940 ;
        RECT 28.890 67.860 29.840 68.620 ;
      LAYER li1 ;
        RECT 30.020 67.980 30.270 68.690 ;
      LAYER li1 ;
        RECT 30.450 68.620 30.480 68.790 ;
        RECT 30.650 68.620 30.840 68.790 ;
        RECT 31.010 68.620 31.200 68.790 ;
        RECT 31.370 68.620 31.400 68.790 ;
        RECT 32.010 68.790 32.960 68.820 ;
        RECT 30.450 68.160 31.400 68.620 ;
      LAYER li1 ;
        RECT 31.580 67.980 31.830 68.690 ;
        RECT 30.020 67.810 31.830 67.980 ;
      LAYER li1 ;
        RECT 32.010 68.620 32.040 68.790 ;
        RECT 32.210 68.620 32.400 68.790 ;
        RECT 32.570 68.620 32.760 68.790 ;
        RECT 32.930 68.620 32.960 68.790 ;
        RECT 33.770 68.790 35.380 68.820 ;
        RECT 32.010 67.940 32.960 68.620 ;
      LAYER li1 ;
        RECT 30.020 67.640 30.190 67.810 ;
      LAYER li1 ;
        RECT 33.140 67.760 33.470 68.690 ;
        RECT 33.770 68.620 33.820 68.790 ;
        RECT 33.990 68.620 34.260 68.790 ;
        RECT 34.430 68.620 34.700 68.790 ;
        RECT 34.870 68.620 35.110 68.790 ;
        RECT 35.280 68.620 35.380 68.790 ;
        RECT 33.770 68.340 35.380 68.620 ;
        RECT 27.900 66.500 28.230 67.490 ;
      LAYER li1 ;
        RECT 28.930 67.410 30.190 67.640 ;
      LAYER li1 ;
        RECT 32.230 67.630 33.470 67.760 ;
        RECT 30.370 67.590 33.470 67.630 ;
        RECT 30.370 67.460 32.400 67.590 ;
      LAYER li1 ;
        RECT 30.020 67.280 30.190 67.410 ;
        RECT 30.020 67.110 31.910 67.280 ;
      LAYER li1 ;
        RECT 27.130 65.630 28.580 66.500 ;
        RECT 27.130 65.460 27.380 65.630 ;
        RECT 27.550 65.460 27.740 65.630 ;
        RECT 27.910 65.460 28.180 65.630 ;
        RECT 28.350 65.460 28.580 65.630 ;
        RECT 27.130 65.430 28.580 65.460 ;
        RECT 28.890 65.680 29.840 67.010 ;
        RECT 28.890 65.510 28.920 65.680 ;
        RECT 29.090 65.510 29.280 65.680 ;
        RECT 29.450 65.510 29.640 65.680 ;
        RECT 29.810 65.510 29.840 65.680 ;
        RECT 28.890 65.430 29.840 65.510 ;
      LAYER li1 ;
        RECT 30.020 65.430 30.270 67.110 ;
      LAYER li1 ;
        RECT 30.450 65.680 31.400 66.930 ;
        RECT 30.450 65.510 30.480 65.680 ;
        RECT 30.650 65.510 30.840 65.680 ;
        RECT 31.010 65.510 31.200 65.680 ;
        RECT 31.370 65.510 31.400 65.680 ;
        RECT 30.450 65.430 31.400 65.510 ;
      LAYER li1 ;
        RECT 31.580 65.430 31.910 67.110 ;
        RECT 32.690 67.070 33.020 67.410 ;
      LAYER li1 ;
        RECT 32.090 65.680 33.040 66.890 ;
        RECT 32.090 65.510 32.120 65.680 ;
        RECT 32.290 65.510 32.480 65.680 ;
        RECT 32.650 65.510 32.840 65.680 ;
        RECT 33.010 65.510 33.040 65.680 ;
        RECT 32.090 65.430 33.040 65.510 ;
        RECT 33.220 65.430 33.470 67.590 ;
        RECT 34.080 67.940 35.380 68.340 ;
        RECT 35.610 68.790 36.200 68.820 ;
        RECT 35.610 68.620 35.640 68.790 ;
        RECT 35.810 68.620 36.000 68.790 ;
        RECT 36.170 68.620 36.200 68.790 ;
        RECT 37.130 68.790 38.740 68.820 ;
        RECT 34.080 67.160 34.410 67.940 ;
        RECT 35.610 67.860 36.200 68.620 ;
        RECT 34.620 66.500 34.950 67.490 ;
      LAYER li1 ;
        RECT 35.650 67.250 36.360 67.640 ;
        RECT 36.540 67.010 36.870 68.690 ;
      LAYER li1 ;
        RECT 37.130 68.620 37.180 68.790 ;
        RECT 37.350 68.620 37.620 68.790 ;
        RECT 37.790 68.620 38.060 68.790 ;
        RECT 38.230 68.620 38.470 68.790 ;
        RECT 38.640 68.620 38.740 68.790 ;
        RECT 37.130 68.340 38.740 68.620 ;
        RECT 37.440 67.940 38.740 68.340 ;
        RECT 38.970 68.790 39.920 68.820 ;
        RECT 38.970 68.620 39.000 68.790 ;
        RECT 39.170 68.620 39.360 68.790 ;
        RECT 39.530 68.620 39.720 68.790 ;
        RECT 39.890 68.620 39.920 68.790 ;
        RECT 40.530 68.790 41.480 68.820 ;
        RECT 37.440 67.160 37.770 67.940 ;
        RECT 38.970 67.860 39.920 68.620 ;
      LAYER li1 ;
        RECT 40.100 67.980 40.350 68.690 ;
      LAYER li1 ;
        RECT 40.530 68.620 40.560 68.790 ;
        RECT 40.730 68.620 40.920 68.790 ;
        RECT 41.090 68.620 41.280 68.790 ;
        RECT 41.450 68.620 41.480 68.790 ;
        RECT 42.090 68.790 43.040 68.820 ;
        RECT 40.530 68.160 41.480 68.620 ;
      LAYER li1 ;
        RECT 41.660 67.980 41.910 68.690 ;
        RECT 40.100 67.810 41.910 67.980 ;
      LAYER li1 ;
        RECT 42.090 68.620 42.120 68.790 ;
        RECT 42.290 68.620 42.480 68.790 ;
        RECT 42.650 68.620 42.840 68.790 ;
        RECT 43.010 68.620 43.040 68.790 ;
        RECT 44.260 68.800 46.990 68.830 ;
        RECT 42.090 67.940 43.040 68.620 ;
      LAYER li1 ;
        RECT 40.100 67.640 40.270 67.810 ;
      LAYER li1 ;
        RECT 43.220 67.760 43.550 68.690 ;
        RECT 44.260 68.630 44.430 68.800 ;
        RECT 44.600 68.630 44.870 68.800 ;
        RECT 45.040 68.630 45.280 68.800 ;
        RECT 45.450 68.630 45.710 68.800 ;
        RECT 45.880 68.630 46.150 68.800 ;
        RECT 46.320 68.630 46.560 68.800 ;
        RECT 46.730 68.630 46.990 68.800 ;
        RECT 44.260 67.830 46.990 68.630 ;
        RECT 48.090 68.790 49.040 68.820 ;
        RECT 48.090 68.620 48.120 68.790 ;
        RECT 48.290 68.620 48.480 68.790 ;
        RECT 48.650 68.620 48.840 68.790 ;
        RECT 49.010 68.620 49.040 68.790 ;
        RECT 49.650 68.790 50.600 68.820 ;
        RECT 48.090 67.860 49.040 68.620 ;
      LAYER li1 ;
        RECT 49.220 67.980 49.470 68.690 ;
      LAYER li1 ;
        RECT 49.650 68.620 49.680 68.790 ;
        RECT 49.850 68.620 50.040 68.790 ;
        RECT 50.210 68.620 50.400 68.790 ;
        RECT 50.570 68.620 50.600 68.790 ;
        RECT 51.210 68.790 52.160 68.820 ;
        RECT 49.650 68.160 50.600 68.620 ;
      LAYER li1 ;
        RECT 50.780 67.980 51.030 68.690 ;
      LAYER li1 ;
        RECT 33.850 65.630 35.300 66.500 ;
        RECT 33.850 65.460 34.100 65.630 ;
        RECT 34.270 65.460 34.460 65.630 ;
        RECT 34.630 65.460 34.900 65.630 ;
        RECT 35.070 65.460 35.300 65.630 ;
        RECT 33.850 65.430 35.300 65.460 ;
        RECT 35.610 65.680 36.200 67.010 ;
        RECT 35.610 65.510 35.640 65.680 ;
        RECT 35.810 65.510 36.000 65.680 ;
        RECT 36.170 65.510 36.200 65.680 ;
        RECT 35.610 65.430 36.200 65.510 ;
      LAYER li1 ;
        RECT 36.480 65.430 36.870 67.010 ;
      LAYER li1 ;
        RECT 37.980 66.500 38.310 67.490 ;
      LAYER li1 ;
        RECT 39.010 67.410 40.270 67.640 ;
      LAYER li1 ;
        RECT 42.310 67.630 43.550 67.760 ;
        RECT 40.450 67.590 43.550 67.630 ;
        RECT 40.450 67.460 42.480 67.590 ;
      LAYER li1 ;
        RECT 40.100 67.280 40.270 67.410 ;
        RECT 40.100 67.110 41.990 67.280 ;
      LAYER li1 ;
        RECT 37.210 65.630 38.660 66.500 ;
        RECT 37.210 65.460 37.460 65.630 ;
        RECT 37.630 65.460 37.820 65.630 ;
        RECT 37.990 65.460 38.260 65.630 ;
        RECT 38.430 65.460 38.660 65.630 ;
        RECT 37.210 65.430 38.660 65.460 ;
        RECT 38.970 65.680 39.920 67.010 ;
        RECT 38.970 65.510 39.000 65.680 ;
        RECT 39.170 65.510 39.360 65.680 ;
        RECT 39.530 65.510 39.720 65.680 ;
        RECT 39.890 65.510 39.920 65.680 ;
        RECT 38.970 65.430 39.920 65.510 ;
      LAYER li1 ;
        RECT 40.100 65.430 40.350 67.110 ;
      LAYER li1 ;
        RECT 40.530 65.680 41.480 66.930 ;
        RECT 40.530 65.510 40.560 65.680 ;
        RECT 40.730 65.510 40.920 65.680 ;
        RECT 41.090 65.510 41.280 65.680 ;
        RECT 41.450 65.510 41.480 65.680 ;
        RECT 40.530 65.430 41.480 65.510 ;
      LAYER li1 ;
        RECT 41.660 65.430 41.990 67.110 ;
        RECT 42.770 67.070 43.100 67.410 ;
      LAYER li1 ;
        RECT 42.170 65.680 43.120 66.890 ;
        RECT 42.170 65.510 42.200 65.680 ;
        RECT 42.370 65.510 42.560 65.680 ;
        RECT 42.730 65.510 42.920 65.680 ;
        RECT 43.090 65.510 43.120 65.680 ;
        RECT 42.170 65.430 43.120 65.510 ;
        RECT 43.300 65.430 43.550 67.590 ;
        RECT 44.420 67.160 44.750 67.830 ;
        RECT 45.150 66.510 45.480 67.490 ;
        RECT 45.700 67.160 46.030 67.830 ;
      LAYER li1 ;
        RECT 49.220 67.810 51.030 67.980 ;
      LAYER li1 ;
        RECT 51.210 68.620 51.240 68.790 ;
        RECT 51.410 68.620 51.600 68.790 ;
        RECT 51.770 68.620 51.960 68.790 ;
        RECT 52.130 68.620 52.160 68.790 ;
        RECT 53.380 68.800 56.110 68.830 ;
        RECT 51.210 67.940 52.160 68.620 ;
      LAYER li1 ;
        RECT 49.220 67.640 49.390 67.810 ;
      LAYER li1 ;
        RECT 52.340 67.760 52.670 68.690 ;
        RECT 53.380 68.630 53.550 68.800 ;
        RECT 53.720 68.630 53.990 68.800 ;
        RECT 54.160 68.630 54.400 68.800 ;
        RECT 54.570 68.630 54.830 68.800 ;
        RECT 55.000 68.630 55.270 68.800 ;
        RECT 55.440 68.630 55.680 68.800 ;
        RECT 55.850 68.630 56.110 68.800 ;
        RECT 53.380 67.830 56.110 68.630 ;
        RECT 57.690 68.790 58.640 68.820 ;
        RECT 57.690 68.620 57.720 68.790 ;
        RECT 57.890 68.620 58.080 68.790 ;
        RECT 58.250 68.620 58.440 68.790 ;
        RECT 58.610 68.620 58.640 68.790 ;
        RECT 59.250 68.790 60.200 68.820 ;
        RECT 57.690 67.860 58.640 68.620 ;
      LAYER li1 ;
        RECT 58.820 67.980 59.070 68.690 ;
      LAYER li1 ;
        RECT 59.250 68.620 59.280 68.790 ;
        RECT 59.450 68.620 59.640 68.790 ;
        RECT 59.810 68.620 60.000 68.790 ;
        RECT 60.170 68.620 60.200 68.790 ;
        RECT 60.810 68.790 61.760 68.820 ;
        RECT 59.250 68.160 60.200 68.620 ;
      LAYER li1 ;
        RECT 60.380 67.980 60.630 68.690 ;
      LAYER li1 ;
        RECT 46.430 66.510 46.760 67.490 ;
      LAYER li1 ;
        RECT 48.130 67.410 49.390 67.640 ;
      LAYER li1 ;
        RECT 51.430 67.630 52.670 67.760 ;
        RECT 49.570 67.590 52.670 67.630 ;
        RECT 49.570 67.460 51.600 67.590 ;
      LAYER li1 ;
        RECT 49.220 67.280 49.390 67.410 ;
        RECT 49.220 67.110 51.110 67.280 ;
      LAYER li1 ;
        RECT 44.180 65.630 46.920 66.510 ;
        RECT 44.180 65.460 44.390 65.630 ;
        RECT 44.560 65.460 44.830 65.630 ;
        RECT 45.000 65.460 45.240 65.630 ;
        RECT 45.410 65.460 45.670 65.630 ;
        RECT 45.840 65.460 46.110 65.630 ;
        RECT 46.280 65.460 46.520 65.630 ;
        RECT 46.690 65.460 46.920 65.630 ;
        RECT 44.180 65.440 46.920 65.460 ;
        RECT 48.090 65.680 49.040 67.010 ;
        RECT 48.090 65.510 48.120 65.680 ;
        RECT 48.290 65.510 48.480 65.680 ;
        RECT 48.650 65.510 48.840 65.680 ;
        RECT 49.010 65.510 49.040 65.680 ;
        RECT 48.090 65.430 49.040 65.510 ;
      LAYER li1 ;
        RECT 49.220 65.430 49.470 67.110 ;
      LAYER li1 ;
        RECT 49.650 65.680 50.600 66.930 ;
        RECT 49.650 65.510 49.680 65.680 ;
        RECT 49.850 65.510 50.040 65.680 ;
        RECT 50.210 65.510 50.400 65.680 ;
        RECT 50.570 65.510 50.600 65.680 ;
        RECT 49.650 65.430 50.600 65.510 ;
      LAYER li1 ;
        RECT 50.780 65.430 51.110 67.110 ;
        RECT 51.890 67.070 52.220 67.410 ;
      LAYER li1 ;
        RECT 51.290 65.680 52.240 66.890 ;
        RECT 51.290 65.510 51.320 65.680 ;
        RECT 51.490 65.510 51.680 65.680 ;
        RECT 51.850 65.510 52.040 65.680 ;
        RECT 52.210 65.510 52.240 65.680 ;
        RECT 51.290 65.430 52.240 65.510 ;
        RECT 52.420 65.430 52.670 67.590 ;
        RECT 53.540 67.160 53.870 67.830 ;
        RECT 54.270 66.510 54.600 67.490 ;
        RECT 54.820 67.160 55.150 67.830 ;
      LAYER li1 ;
        RECT 58.820 67.810 60.630 67.980 ;
      LAYER li1 ;
        RECT 60.810 68.620 60.840 68.790 ;
        RECT 61.010 68.620 61.200 68.790 ;
        RECT 61.370 68.620 61.560 68.790 ;
        RECT 61.730 68.620 61.760 68.790 ;
        RECT 62.570 68.790 64.180 68.820 ;
        RECT 60.810 67.940 61.760 68.620 ;
      LAYER li1 ;
        RECT 58.820 67.640 58.990 67.810 ;
      LAYER li1 ;
        RECT 61.940 67.760 62.270 68.690 ;
        RECT 62.570 68.620 62.620 68.790 ;
        RECT 62.790 68.620 63.060 68.790 ;
        RECT 63.230 68.620 63.500 68.790 ;
        RECT 63.670 68.620 63.910 68.790 ;
        RECT 64.080 68.620 64.180 68.790 ;
        RECT 62.570 68.340 64.180 68.620 ;
        RECT 55.550 66.510 55.880 67.490 ;
      LAYER li1 ;
        RECT 57.730 67.410 58.990 67.640 ;
      LAYER li1 ;
        RECT 61.030 67.630 62.270 67.760 ;
        RECT 59.170 67.590 62.270 67.630 ;
        RECT 59.170 67.460 61.200 67.590 ;
      LAYER li1 ;
        RECT 58.820 67.280 58.990 67.410 ;
        RECT 58.820 67.110 60.710 67.280 ;
      LAYER li1 ;
        RECT 53.300 65.630 56.040 66.510 ;
        RECT 53.300 65.460 53.510 65.630 ;
        RECT 53.680 65.460 53.950 65.630 ;
        RECT 54.120 65.460 54.360 65.630 ;
        RECT 54.530 65.460 54.790 65.630 ;
        RECT 54.960 65.460 55.230 65.630 ;
        RECT 55.400 65.460 55.640 65.630 ;
        RECT 55.810 65.460 56.040 65.630 ;
        RECT 53.300 65.440 56.040 65.460 ;
        RECT 57.690 65.680 58.640 67.010 ;
        RECT 57.690 65.510 57.720 65.680 ;
        RECT 57.890 65.510 58.080 65.680 ;
        RECT 58.250 65.510 58.440 65.680 ;
        RECT 58.610 65.510 58.640 65.680 ;
        RECT 57.690 65.430 58.640 65.510 ;
      LAYER li1 ;
        RECT 58.820 65.430 59.070 67.110 ;
      LAYER li1 ;
        RECT 59.250 65.680 60.200 66.930 ;
        RECT 59.250 65.510 59.280 65.680 ;
        RECT 59.450 65.510 59.640 65.680 ;
        RECT 59.810 65.510 60.000 65.680 ;
        RECT 60.170 65.510 60.200 65.680 ;
        RECT 59.250 65.430 60.200 65.510 ;
      LAYER li1 ;
        RECT 60.380 65.430 60.710 67.110 ;
        RECT 61.490 67.070 61.820 67.410 ;
      LAYER li1 ;
        RECT 60.890 65.680 61.840 66.890 ;
        RECT 60.890 65.510 60.920 65.680 ;
        RECT 61.090 65.510 61.280 65.680 ;
        RECT 61.450 65.510 61.640 65.680 ;
        RECT 61.810 65.510 61.840 65.680 ;
        RECT 60.890 65.430 61.840 65.510 ;
        RECT 62.020 65.430 62.270 67.590 ;
        RECT 62.880 67.940 64.180 68.340 ;
        RECT 64.410 68.790 65.360 68.820 ;
        RECT 64.410 68.620 64.440 68.790 ;
        RECT 64.610 68.620 64.800 68.790 ;
        RECT 64.970 68.620 65.160 68.790 ;
        RECT 65.330 68.620 65.360 68.790 ;
        RECT 65.970 68.790 66.920 68.820 ;
        RECT 62.880 67.160 63.210 67.940 ;
        RECT 64.410 67.860 65.360 68.620 ;
      LAYER li1 ;
        RECT 65.540 67.980 65.790 68.690 ;
      LAYER li1 ;
        RECT 65.970 68.620 66.000 68.790 ;
        RECT 66.170 68.620 66.360 68.790 ;
        RECT 66.530 68.620 66.720 68.790 ;
        RECT 66.890 68.620 66.920 68.790 ;
        RECT 67.530 68.790 68.480 68.820 ;
        RECT 65.970 68.160 66.920 68.620 ;
      LAYER li1 ;
        RECT 67.100 67.980 67.350 68.690 ;
        RECT 65.540 67.810 67.350 67.980 ;
      LAYER li1 ;
        RECT 67.530 68.620 67.560 68.790 ;
        RECT 67.730 68.620 67.920 68.790 ;
        RECT 68.090 68.620 68.280 68.790 ;
        RECT 68.450 68.620 68.480 68.790 ;
        RECT 69.290 68.790 70.900 68.820 ;
        RECT 67.530 67.940 68.480 68.620 ;
      LAYER li1 ;
        RECT 65.540 67.640 65.710 67.810 ;
      LAYER li1 ;
        RECT 68.660 67.760 68.990 68.690 ;
        RECT 69.290 68.620 69.340 68.790 ;
        RECT 69.510 68.620 69.780 68.790 ;
        RECT 69.950 68.620 70.220 68.790 ;
        RECT 70.390 68.620 70.630 68.790 ;
        RECT 70.800 68.620 70.900 68.790 ;
        RECT 69.290 68.340 70.900 68.620 ;
        RECT 63.420 66.500 63.750 67.490 ;
      LAYER li1 ;
        RECT 64.450 67.410 65.710 67.640 ;
      LAYER li1 ;
        RECT 67.750 67.630 68.990 67.760 ;
        RECT 65.890 67.590 68.990 67.630 ;
        RECT 65.890 67.460 67.920 67.590 ;
      LAYER li1 ;
        RECT 65.540 67.280 65.710 67.410 ;
        RECT 65.540 67.110 67.430 67.280 ;
      LAYER li1 ;
        RECT 62.650 65.630 64.100 66.500 ;
        RECT 62.650 65.460 62.900 65.630 ;
        RECT 63.070 65.460 63.260 65.630 ;
        RECT 63.430 65.460 63.700 65.630 ;
        RECT 63.870 65.460 64.100 65.630 ;
        RECT 62.650 65.430 64.100 65.460 ;
        RECT 64.410 65.680 65.360 67.010 ;
        RECT 64.410 65.510 64.440 65.680 ;
        RECT 64.610 65.510 64.800 65.680 ;
        RECT 64.970 65.510 65.160 65.680 ;
        RECT 65.330 65.510 65.360 65.680 ;
        RECT 64.410 65.430 65.360 65.510 ;
      LAYER li1 ;
        RECT 65.540 65.430 65.790 67.110 ;
      LAYER li1 ;
        RECT 65.970 65.680 66.920 66.930 ;
        RECT 65.970 65.510 66.000 65.680 ;
        RECT 66.170 65.510 66.360 65.680 ;
        RECT 66.530 65.510 66.720 65.680 ;
        RECT 66.890 65.510 66.920 65.680 ;
        RECT 65.970 65.430 66.920 65.510 ;
      LAYER li1 ;
        RECT 67.100 65.430 67.430 67.110 ;
        RECT 68.210 67.070 68.540 67.410 ;
      LAYER li1 ;
        RECT 67.610 65.680 68.560 66.890 ;
        RECT 67.610 65.510 67.640 65.680 ;
        RECT 67.810 65.510 68.000 65.680 ;
        RECT 68.170 65.510 68.360 65.680 ;
        RECT 68.530 65.510 68.560 65.680 ;
        RECT 67.610 65.430 68.560 65.510 ;
        RECT 68.740 65.430 68.990 67.590 ;
        RECT 69.600 67.940 70.900 68.340 ;
        RECT 71.130 68.790 72.080 68.820 ;
        RECT 71.130 68.620 71.160 68.790 ;
        RECT 71.330 68.620 71.520 68.790 ;
        RECT 71.690 68.620 71.880 68.790 ;
        RECT 72.050 68.620 72.080 68.790 ;
        RECT 72.690 68.790 73.640 68.820 ;
        RECT 69.600 67.160 69.930 67.940 ;
        RECT 71.130 67.860 72.080 68.620 ;
      LAYER li1 ;
        RECT 72.260 67.980 72.510 68.690 ;
      LAYER li1 ;
        RECT 72.690 68.620 72.720 68.790 ;
        RECT 72.890 68.620 73.080 68.790 ;
        RECT 73.250 68.620 73.440 68.790 ;
        RECT 73.610 68.620 73.640 68.790 ;
        RECT 74.250 68.790 75.200 68.820 ;
        RECT 72.690 68.160 73.640 68.620 ;
      LAYER li1 ;
        RECT 73.820 67.980 74.070 68.690 ;
        RECT 72.260 67.810 74.070 67.980 ;
      LAYER li1 ;
        RECT 74.250 68.620 74.280 68.790 ;
        RECT 74.450 68.620 74.640 68.790 ;
        RECT 74.810 68.620 75.000 68.790 ;
        RECT 75.170 68.620 75.200 68.790 ;
        RECT 76.010 68.790 77.620 68.820 ;
        RECT 74.250 67.940 75.200 68.620 ;
      LAYER li1 ;
        RECT 72.260 67.640 72.430 67.810 ;
      LAYER li1 ;
        RECT 75.380 67.760 75.710 68.690 ;
        RECT 76.010 68.620 76.060 68.790 ;
        RECT 76.230 68.620 76.500 68.790 ;
        RECT 76.670 68.620 76.940 68.790 ;
        RECT 77.110 68.620 77.350 68.790 ;
        RECT 77.520 68.620 77.620 68.790 ;
        RECT 76.010 68.340 77.620 68.620 ;
        RECT 70.140 66.500 70.470 67.490 ;
      LAYER li1 ;
        RECT 71.170 67.410 72.430 67.640 ;
      LAYER li1 ;
        RECT 74.470 67.630 75.710 67.760 ;
        RECT 72.610 67.590 75.710 67.630 ;
        RECT 72.610 67.460 74.640 67.590 ;
      LAYER li1 ;
        RECT 72.260 67.280 72.430 67.410 ;
        RECT 72.260 67.110 74.150 67.280 ;
      LAYER li1 ;
        RECT 69.370 65.630 70.820 66.500 ;
        RECT 69.370 65.460 69.620 65.630 ;
        RECT 69.790 65.460 69.980 65.630 ;
        RECT 70.150 65.460 70.420 65.630 ;
        RECT 70.590 65.460 70.820 65.630 ;
        RECT 69.370 65.430 70.820 65.460 ;
        RECT 71.130 65.680 72.080 67.010 ;
        RECT 71.130 65.510 71.160 65.680 ;
        RECT 71.330 65.510 71.520 65.680 ;
        RECT 71.690 65.510 71.880 65.680 ;
        RECT 72.050 65.510 72.080 65.680 ;
        RECT 71.130 65.430 72.080 65.510 ;
      LAYER li1 ;
        RECT 72.260 65.430 72.510 67.110 ;
      LAYER li1 ;
        RECT 72.690 65.680 73.640 66.930 ;
        RECT 72.690 65.510 72.720 65.680 ;
        RECT 72.890 65.510 73.080 65.680 ;
        RECT 73.250 65.510 73.440 65.680 ;
        RECT 73.610 65.510 73.640 65.680 ;
        RECT 72.690 65.430 73.640 65.510 ;
      LAYER li1 ;
        RECT 73.820 65.430 74.150 67.110 ;
        RECT 74.930 67.070 75.260 67.410 ;
      LAYER li1 ;
        RECT 74.330 65.680 75.280 66.890 ;
        RECT 74.330 65.510 74.360 65.680 ;
        RECT 74.530 65.510 74.720 65.680 ;
        RECT 74.890 65.510 75.080 65.680 ;
        RECT 75.250 65.510 75.280 65.680 ;
        RECT 74.330 65.430 75.280 65.510 ;
        RECT 75.460 65.430 75.710 67.590 ;
        RECT 76.320 67.940 77.620 68.340 ;
        RECT 77.850 68.790 79.470 68.820 ;
        RECT 81.290 68.790 82.900 68.820 ;
        RECT 83.680 68.790 85.290 68.820 ;
        RECT 85.900 68.790 87.210 68.820 ;
        RECT 77.850 68.620 77.860 68.790 ;
        RECT 78.030 68.620 78.220 68.790 ;
        RECT 78.390 68.620 78.580 68.790 ;
        RECT 78.750 68.620 78.940 68.790 ;
        RECT 79.110 68.620 79.300 68.790 ;
        RECT 76.320 67.160 76.650 67.940 ;
        RECT 77.850 67.860 79.470 68.620 ;
        RECT 76.860 66.500 77.190 67.490 ;
      LAYER li1 ;
        RECT 77.890 67.350 78.760 67.680 ;
        RECT 79.650 67.460 80.040 68.380 ;
        RECT 80.220 67.460 80.490 68.380 ;
        RECT 80.670 67.860 81.000 68.690 ;
      LAYER li1 ;
        RECT 81.290 68.620 81.340 68.790 ;
        RECT 81.510 68.620 81.780 68.790 ;
        RECT 81.950 68.620 82.220 68.790 ;
        RECT 82.390 68.620 82.630 68.790 ;
        RECT 82.800 68.620 82.900 68.790 ;
        RECT 81.290 68.340 82.900 68.620 ;
      LAYER li1 ;
        RECT 80.740 67.280 81.000 67.860 ;
        RECT 78.960 67.110 81.000 67.280 ;
      LAYER li1 ;
        RECT 81.600 67.940 82.900 68.340 ;
        RECT 81.600 67.160 81.930 67.940 ;
      LAYER li1 ;
        RECT 83.150 67.860 83.500 68.690 ;
      LAYER li1 ;
        RECT 83.850 68.620 84.040 68.790 ;
        RECT 84.210 68.620 84.400 68.790 ;
        RECT 84.570 68.620 84.760 68.790 ;
        RECT 84.930 68.620 85.120 68.790 ;
        RECT 83.680 67.860 85.290 68.620 ;
        RECT 85.470 67.860 85.720 68.690 ;
        RECT 85.900 68.620 85.930 68.790 ;
        RECT 86.100 68.620 86.290 68.790 ;
        RECT 86.460 68.620 86.650 68.790 ;
        RECT 86.820 68.620 87.010 68.790 ;
        RECT 87.180 68.620 87.210 68.790 ;
        RECT 85.900 67.860 87.210 68.620 ;
        RECT 87.940 68.800 90.670 68.830 ;
        RECT 87.940 68.630 88.110 68.800 ;
        RECT 88.280 68.630 88.550 68.800 ;
        RECT 88.720 68.630 88.960 68.800 ;
        RECT 89.130 68.630 89.390 68.800 ;
        RECT 89.560 68.630 89.830 68.800 ;
        RECT 90.000 68.630 90.240 68.800 ;
        RECT 90.410 68.630 90.670 68.800 ;
        RECT 92.240 68.790 93.190 68.820 ;
        RECT 76.090 65.630 77.540 66.500 ;
        RECT 76.090 65.460 76.340 65.630 ;
        RECT 76.510 65.460 76.700 65.630 ;
        RECT 76.870 65.460 77.140 65.630 ;
        RECT 77.310 65.460 77.540 65.630 ;
        RECT 76.090 65.430 77.540 65.460 ;
        RECT 77.850 65.680 78.780 67.010 ;
        RECT 77.850 65.510 77.870 65.680 ;
        RECT 78.040 65.510 78.230 65.680 ;
        RECT 78.400 65.510 78.590 65.680 ;
        RECT 78.760 65.510 78.780 65.680 ;
        RECT 77.850 65.430 78.780 65.510 ;
      LAYER li1 ;
        RECT 78.960 65.430 79.130 67.110 ;
      LAYER li1 ;
        RECT 79.310 65.680 80.560 66.930 ;
        RECT 79.480 65.510 79.670 65.680 ;
        RECT 79.840 65.510 80.030 65.680 ;
        RECT 80.200 65.510 80.390 65.680 ;
        RECT 79.310 65.430 80.560 65.510 ;
      LAYER li1 ;
        RECT 80.740 65.430 81.000 67.110 ;
      LAYER li1 ;
        RECT 82.140 66.500 82.470 67.490 ;
        RECT 81.370 65.630 82.820 66.500 ;
        RECT 81.370 65.460 81.620 65.630 ;
        RECT 81.790 65.460 81.980 65.630 ;
        RECT 82.150 65.460 82.420 65.630 ;
        RECT 82.590 65.460 82.820 65.630 ;
        RECT 81.370 65.430 82.820 65.460 ;
      LAYER li1 ;
        RECT 83.150 65.450 83.400 67.860 ;
      LAYER li1 ;
        RECT 83.610 67.260 83.940 67.460 ;
      LAYER li1 ;
        RECT 84.130 67.440 85.320 67.680 ;
      LAYER li1 ;
        RECT 85.500 67.260 85.670 67.860 ;
        RECT 87.940 67.830 90.670 68.630 ;
      LAYER li1 ;
        RECT 85.850 67.350 86.760 67.680 ;
        RECT 86.940 67.350 87.240 67.680 ;
      LAYER li1 ;
        RECT 83.610 67.090 85.670 67.260 ;
        RECT 88.100 67.160 88.430 67.830 ;
        RECT 83.580 65.680 84.480 66.910 ;
        RECT 83.580 65.510 83.590 65.680 ;
        RECT 83.760 65.510 83.950 65.680 ;
        RECT 84.120 65.510 84.310 65.680 ;
        RECT 83.580 65.430 84.480 65.510 ;
        RECT 84.660 65.430 84.910 67.090 ;
        RECT 87.000 66.910 87.250 66.990 ;
        RECT 85.360 66.740 87.250 66.910 ;
        RECT 85.360 65.430 85.690 66.740 ;
        RECT 85.870 65.680 86.820 66.560 ;
        RECT 85.870 65.510 85.900 65.680 ;
        RECT 86.070 65.510 86.260 65.680 ;
        RECT 86.430 65.510 86.620 65.680 ;
        RECT 86.790 65.510 86.820 65.680 ;
        RECT 85.870 65.430 86.820 65.510 ;
        RECT 87.000 65.450 87.250 66.740 ;
        RECT 88.830 66.510 89.160 67.490 ;
        RECT 89.380 67.160 89.710 67.830 ;
        RECT 90.110 66.510 90.440 67.490 ;
        RECT 91.790 66.830 92.060 68.690 ;
        RECT 92.240 68.620 92.270 68.790 ;
        RECT 92.440 68.620 92.630 68.790 ;
        RECT 92.800 68.620 92.990 68.790 ;
        RECT 93.160 68.620 93.190 68.790 ;
        RECT 93.880 68.790 94.470 68.820 ;
        RECT 92.240 68.190 93.190 68.620 ;
        RECT 93.370 68.190 93.700 68.690 ;
        RECT 92.920 66.830 93.250 67.330 ;
        RECT 91.790 66.660 93.250 66.830 ;
        RECT 87.860 65.630 90.600 66.510 ;
        RECT 91.790 65.730 92.120 66.660 ;
        RECT 87.860 65.460 88.070 65.630 ;
        RECT 88.240 65.460 88.510 65.630 ;
        RECT 88.680 65.460 88.920 65.630 ;
        RECT 89.090 65.460 89.350 65.630 ;
        RECT 89.520 65.460 89.790 65.630 ;
        RECT 89.960 65.460 90.200 65.630 ;
        RECT 90.370 65.460 90.600 65.630 ;
        RECT 92.310 65.680 92.900 66.460 ;
        RECT 92.310 65.510 92.340 65.680 ;
        RECT 92.510 65.510 92.700 65.680 ;
        RECT 92.870 65.510 92.900 65.680 ;
        RECT 92.310 65.480 92.900 65.510 ;
        RECT 93.080 65.550 93.250 66.660 ;
        RECT 93.430 67.270 93.700 68.190 ;
        RECT 93.880 68.620 93.910 68.790 ;
        RECT 94.080 68.620 94.270 68.790 ;
        RECT 94.440 68.620 94.470 68.790 ;
        RECT 98.840 68.790 99.790 68.820 ;
        RECT 93.880 67.940 94.470 68.620 ;
      LAYER li1 ;
        RECT 94.750 68.560 97.690 68.730 ;
        RECT 94.750 67.570 94.920 68.560 ;
      LAYER li1 ;
        RECT 93.430 67.040 93.960 67.270 ;
        RECT 93.430 65.730 93.680 67.040 ;
      LAYER li1 ;
        RECT 94.380 66.700 94.920 67.570 ;
        RECT 95.100 67.080 95.430 68.380 ;
      LAYER li1 ;
        RECT 95.610 67.860 95.880 68.360 ;
        RECT 96.330 68.110 96.660 68.360 ;
        RECT 96.330 67.940 97.340 68.110 ;
        RECT 95.610 66.870 95.780 67.860 ;
        RECT 96.660 67.270 96.990 67.760 ;
        RECT 95.560 66.700 95.780 66.870 ;
        RECT 95.960 67.040 96.990 67.270 ;
        RECT 97.170 67.710 97.340 67.940 ;
      LAYER li1 ;
        RECT 97.520 68.060 97.690 68.560 ;
      LAYER li1 ;
        RECT 98.840 68.620 98.870 68.790 ;
        RECT 99.040 68.620 99.230 68.790 ;
        RECT 99.400 68.620 99.590 68.790 ;
        RECT 99.760 68.620 99.790 68.790 ;
        RECT 98.840 68.240 99.790 68.620 ;
      LAYER li1 ;
        RECT 99.970 68.750 102.630 68.920 ;
        RECT 99.970 68.060 100.140 68.750 ;
        RECT 97.520 67.890 100.140 68.060 ;
      LAYER li1 ;
        RECT 97.170 67.540 99.790 67.710 ;
        RECT 95.560 66.520 95.730 66.700 ;
        RECT 95.960 66.520 96.130 67.040 ;
        RECT 97.170 66.860 97.340 67.540 ;
      LAYER li1 ;
        RECT 99.970 67.360 100.140 67.890 ;
      LAYER li1 ;
        RECT 93.920 66.350 95.730 66.520 ;
        RECT 93.920 65.730 94.170 66.350 ;
        RECT 94.350 66.000 95.380 66.170 ;
        RECT 94.350 65.550 94.520 66.000 ;
        RECT 87.860 65.440 90.600 65.460 ;
        RECT 93.080 65.380 94.520 65.550 ;
        RECT 94.700 65.680 95.030 65.820 ;
        RECT 94.700 65.510 94.730 65.680 ;
        RECT 94.900 65.510 95.030 65.680 ;
        RECT 94.700 65.480 95.030 65.510 ;
        RECT 95.210 65.550 95.380 66.000 ;
        RECT 95.560 65.730 95.730 66.350 ;
        RECT 95.910 66.190 96.130 66.520 ;
        RECT 96.310 66.690 97.340 66.860 ;
        RECT 97.520 67.010 97.850 67.360 ;
      LAYER li1 ;
        RECT 98.290 67.190 100.140 67.360 ;
      LAYER li1 ;
        RECT 100.320 67.860 100.650 68.570 ;
        RECT 101.110 68.400 102.280 68.570 ;
        RECT 101.110 67.860 101.440 68.400 ;
        RECT 100.320 67.010 100.580 67.860 ;
        RECT 101.650 67.600 101.930 68.100 ;
        RECT 97.520 66.840 100.580 67.010 ;
        RECT 96.310 65.990 96.480 66.690 ;
        RECT 97.170 66.660 97.340 66.690 ;
        RECT 96.660 66.310 96.990 66.510 ;
        RECT 97.170 66.490 98.940 66.660 ;
        RECT 96.660 66.190 98.430 66.310 ;
        RECT 96.780 66.140 98.430 66.190 ;
        RECT 96.260 65.730 96.590 65.990 ;
        RECT 96.780 65.550 96.950 66.140 ;
        RECT 95.210 65.380 96.950 65.550 ;
        RECT 97.130 65.680 98.080 65.960 ;
        RECT 97.130 65.510 97.160 65.680 ;
        RECT 97.330 65.510 97.520 65.680 ;
        RECT 97.690 65.510 97.880 65.680 ;
        RECT 98.050 65.510 98.080 65.680 ;
        RECT 97.130 65.480 98.080 65.510 ;
        RECT 98.260 65.550 98.430 66.140 ;
        RECT 98.610 65.730 98.940 66.490 ;
        RECT 100.250 66.260 100.580 66.840 ;
        RECT 100.760 67.430 101.930 67.600 ;
        RECT 100.760 66.080 100.930 67.430 ;
        RECT 101.310 66.750 101.640 67.250 ;
        RECT 102.110 67.000 102.280 68.400 ;
      LAYER li1 ;
        RECT 102.460 68.090 102.630 68.750 ;
      LAYER li1 ;
        RECT 102.810 68.790 103.760 68.820 ;
        RECT 102.810 68.620 102.840 68.790 ;
        RECT 103.010 68.620 103.200 68.790 ;
        RECT 103.370 68.620 103.560 68.790 ;
        RECT 103.730 68.620 103.760 68.790 ;
        RECT 105.420 68.790 106.370 68.820 ;
        RECT 102.810 68.270 103.760 68.620 ;
        RECT 104.300 68.190 104.630 68.690 ;
        RECT 105.420 68.620 105.450 68.790 ;
        RECT 105.620 68.620 105.810 68.790 ;
        RECT 105.980 68.620 106.170 68.790 ;
        RECT 106.340 68.620 106.370 68.790 ;
      LAYER li1 ;
        RECT 102.460 67.980 103.470 68.090 ;
        RECT 102.460 67.920 103.520 67.980 ;
        RECT 103.140 67.810 103.520 67.920 ;
      LAYER li1 ;
        RECT 102.490 67.350 102.820 67.740 ;
      LAYER li1 ;
        RECT 103.140 67.530 103.470 67.810 ;
      LAYER li1 ;
        RECT 104.300 67.350 104.530 68.190 ;
        RECT 104.910 67.690 105.240 68.190 ;
        RECT 105.420 67.690 106.370 68.620 ;
        RECT 107.620 68.800 110.350 68.830 ;
        RECT 107.620 68.630 107.790 68.800 ;
        RECT 107.960 68.630 108.230 68.800 ;
        RECT 108.400 68.630 108.640 68.800 ;
        RECT 108.810 68.630 109.070 68.800 ;
        RECT 109.240 68.630 109.510 68.800 ;
        RECT 109.680 68.630 109.920 68.800 ;
        RECT 110.090 68.630 110.350 68.800 ;
        RECT 111.520 68.790 112.410 68.820 ;
        RECT 114.410 68.790 116.020 68.820 ;
        RECT 102.490 67.180 104.530 67.350 ;
        RECT 101.820 66.830 104.180 67.000 ;
        RECT 101.820 66.510 101.990 66.830 ;
        RECT 104.360 66.650 104.530 67.180 ;
        RECT 99.120 65.910 100.930 66.080 ;
        RECT 101.110 66.340 101.990 66.510 ;
        RECT 99.120 65.550 99.290 65.910 ;
        RECT 98.260 65.380 99.290 65.550 ;
        RECT 99.470 65.680 100.420 65.730 ;
        RECT 99.470 65.510 99.500 65.680 ;
        RECT 99.670 65.510 99.860 65.680 ;
        RECT 100.030 65.510 100.220 65.680 ;
        RECT 100.390 65.510 100.420 65.680 ;
        RECT 99.470 65.430 100.420 65.510 ;
        RECT 101.110 65.430 101.360 66.340 ;
        RECT 102.170 65.680 103.120 66.510 ;
        RECT 103.520 66.480 104.530 66.650 ;
        RECT 105.030 67.510 105.240 67.690 ;
        RECT 105.030 67.180 106.400 67.510 ;
        RECT 103.520 66.010 103.770 66.480 ;
        RECT 103.950 65.680 104.850 66.300 ;
        RECT 105.030 66.180 105.280 67.180 ;
        RECT 102.170 65.510 102.200 65.680 ;
        RECT 102.370 65.510 102.560 65.680 ;
        RECT 102.730 65.510 102.920 65.680 ;
        RECT 103.090 65.510 103.120 65.680 ;
        RECT 104.120 65.510 104.310 65.680 ;
        RECT 104.480 65.510 104.670 65.680 ;
        RECT 104.840 65.510 104.850 65.680 ;
        RECT 102.170 65.480 103.120 65.510 ;
        RECT 103.950 65.480 104.850 65.510 ;
        RECT 105.460 65.680 106.400 66.990 ;
        RECT 105.460 65.510 105.480 65.680 ;
        RECT 105.650 65.510 105.840 65.680 ;
        RECT 106.010 65.510 106.200 65.680 ;
        RECT 106.370 65.510 106.400 65.680 ;
        RECT 105.460 65.450 106.400 65.510 ;
      LAYER li1 ;
        RECT 106.580 65.450 106.920 68.520 ;
      LAYER li1 ;
        RECT 107.620 67.830 110.350 68.630 ;
        RECT 111.010 68.080 111.340 68.690 ;
        RECT 111.690 68.620 111.880 68.790 ;
        RECT 112.050 68.620 112.240 68.790 ;
        RECT 111.520 68.260 112.410 68.620 ;
        RECT 112.590 68.080 112.920 68.690 ;
        RECT 111.010 67.910 112.920 68.080 ;
        RECT 111.010 67.860 111.340 67.910 ;
        RECT 107.780 67.160 108.110 67.830 ;
        RECT 108.510 66.510 108.840 67.490 ;
        RECT 109.060 67.160 109.390 67.830 ;
      LAYER li1 ;
        RECT 113.370 67.730 113.700 68.690 ;
      LAYER li1 ;
        RECT 114.410 68.620 114.460 68.790 ;
        RECT 114.630 68.620 114.900 68.790 ;
        RECT 115.070 68.620 115.340 68.790 ;
        RECT 115.510 68.620 115.750 68.790 ;
        RECT 115.920 68.620 116.020 68.790 ;
        RECT 114.410 68.340 116.020 68.620 ;
        RECT 109.790 66.510 110.120 67.490 ;
      LAYER li1 ;
        RECT 111.010 67.350 111.740 67.680 ;
        RECT 111.950 67.430 112.680 67.680 ;
        RECT 112.860 67.560 113.700 67.730 ;
      LAYER li1 ;
        RECT 114.720 67.940 116.020 68.340 ;
        RECT 116.250 68.790 117.200 68.820 ;
        RECT 116.250 68.620 116.280 68.790 ;
        RECT 116.450 68.620 116.640 68.790 ;
        RECT 116.810 68.620 117.000 68.790 ;
        RECT 117.170 68.620 117.200 68.790 ;
        RECT 117.810 68.790 118.760 68.820 ;
      LAYER li1 ;
        RECT 112.860 67.250 113.030 67.560 ;
        RECT 112.450 67.080 113.030 67.250 ;
      LAYER li1 ;
        RECT 107.540 65.630 110.280 66.510 ;
        RECT 107.540 65.460 107.750 65.630 ;
        RECT 107.920 65.460 108.190 65.630 ;
        RECT 108.360 65.460 108.600 65.630 ;
        RECT 108.770 65.460 109.030 65.630 ;
        RECT 109.200 65.460 109.470 65.630 ;
        RECT 109.640 65.460 109.880 65.630 ;
        RECT 110.050 65.460 110.280 65.630 ;
        RECT 107.540 65.440 110.280 65.460 ;
        RECT 110.970 65.680 111.920 67.010 ;
        RECT 110.970 65.510 111.000 65.680 ;
        RECT 111.170 65.510 111.360 65.680 ;
        RECT 111.530 65.510 111.720 65.680 ;
        RECT 111.890 65.510 111.920 65.680 ;
        RECT 110.970 65.430 111.920 65.510 ;
      LAYER li1 ;
        RECT 112.450 65.430 112.920 67.080 ;
        RECT 113.210 67.070 114.120 67.380 ;
      LAYER li1 ;
        RECT 114.720 67.160 115.050 67.940 ;
        RECT 116.250 67.860 117.200 68.620 ;
      LAYER li1 ;
        RECT 117.380 67.980 117.630 68.690 ;
      LAYER li1 ;
        RECT 117.810 68.620 117.840 68.790 ;
        RECT 118.010 68.620 118.200 68.790 ;
        RECT 118.370 68.620 118.560 68.790 ;
        RECT 118.730 68.620 118.760 68.790 ;
        RECT 119.370 68.790 120.320 68.820 ;
        RECT 117.810 68.160 118.760 68.620 ;
      LAYER li1 ;
        RECT 118.940 67.980 119.190 68.690 ;
        RECT 117.380 67.810 119.190 67.980 ;
      LAYER li1 ;
        RECT 119.370 68.620 119.400 68.790 ;
        RECT 119.570 68.620 119.760 68.790 ;
        RECT 119.930 68.620 120.120 68.790 ;
        RECT 120.290 68.620 120.320 68.790 ;
        RECT 121.130 68.790 122.740 68.820 ;
        RECT 119.370 67.940 120.320 68.620 ;
      LAYER li1 ;
        RECT 117.380 67.640 117.550 67.810 ;
      LAYER li1 ;
        RECT 120.500 67.760 120.830 68.690 ;
        RECT 121.130 68.620 121.180 68.790 ;
        RECT 121.350 68.620 121.620 68.790 ;
        RECT 121.790 68.620 122.060 68.790 ;
        RECT 122.230 68.620 122.470 68.790 ;
        RECT 122.640 68.620 122.740 68.790 ;
        RECT 121.130 68.340 122.740 68.620 ;
        RECT 113.100 65.680 114.050 66.890 ;
        RECT 115.260 66.500 115.590 67.490 ;
      LAYER li1 ;
        RECT 116.290 67.410 117.550 67.640 ;
      LAYER li1 ;
        RECT 119.590 67.630 120.830 67.760 ;
        RECT 117.730 67.590 120.830 67.630 ;
        RECT 117.730 67.460 119.760 67.590 ;
      LAYER li1 ;
        RECT 117.380 67.280 117.550 67.410 ;
        RECT 117.380 67.110 119.270 67.280 ;
      LAYER li1 ;
        RECT 113.100 65.510 113.130 65.680 ;
        RECT 113.300 65.510 113.490 65.680 ;
        RECT 113.660 65.510 113.850 65.680 ;
        RECT 114.020 65.510 114.050 65.680 ;
        RECT 113.100 65.430 114.050 65.510 ;
        RECT 114.490 65.630 115.940 66.500 ;
        RECT 114.490 65.460 114.740 65.630 ;
        RECT 114.910 65.460 115.100 65.630 ;
        RECT 115.270 65.460 115.540 65.630 ;
        RECT 115.710 65.460 115.940 65.630 ;
        RECT 114.490 65.430 115.940 65.460 ;
        RECT 116.250 65.680 117.200 67.010 ;
        RECT 116.250 65.510 116.280 65.680 ;
        RECT 116.450 65.510 116.640 65.680 ;
        RECT 116.810 65.510 117.000 65.680 ;
        RECT 117.170 65.510 117.200 65.680 ;
        RECT 116.250 65.430 117.200 65.510 ;
      LAYER li1 ;
        RECT 117.380 65.430 117.630 67.110 ;
      LAYER li1 ;
        RECT 117.810 65.680 118.760 66.930 ;
        RECT 117.810 65.510 117.840 65.680 ;
        RECT 118.010 65.510 118.200 65.680 ;
        RECT 118.370 65.510 118.560 65.680 ;
        RECT 118.730 65.510 118.760 65.680 ;
        RECT 117.810 65.430 118.760 65.510 ;
      LAYER li1 ;
        RECT 118.940 65.430 119.270 67.110 ;
        RECT 120.050 67.070 120.380 67.410 ;
      LAYER li1 ;
        RECT 119.450 65.680 120.400 66.890 ;
        RECT 119.450 65.510 119.480 65.680 ;
        RECT 119.650 65.510 119.840 65.680 ;
        RECT 120.010 65.510 120.200 65.680 ;
        RECT 120.370 65.510 120.400 65.680 ;
        RECT 119.450 65.430 120.400 65.510 ;
        RECT 120.580 65.430 120.830 67.590 ;
        RECT 121.440 67.940 122.740 68.340 ;
        RECT 122.970 68.790 123.560 68.820 ;
        RECT 122.970 68.620 123.000 68.790 ;
        RECT 123.170 68.620 123.360 68.790 ;
        RECT 123.530 68.620 123.560 68.790 ;
        RECT 124.240 68.790 125.190 68.820 ;
        RECT 121.440 67.160 121.770 67.940 ;
        RECT 122.970 67.860 123.560 68.620 ;
      LAYER li1 ;
        RECT 123.810 67.760 124.060 68.690 ;
      LAYER li1 ;
        RECT 124.240 68.620 124.270 68.790 ;
        RECT 124.440 68.620 124.630 68.790 ;
        RECT 124.800 68.620 124.990 68.790 ;
        RECT 125.160 68.620 125.190 68.790 ;
        RECT 126.820 68.800 129.550 68.830 ;
        RECT 124.240 67.940 125.190 68.620 ;
      LAYER li1 ;
        RECT 125.370 67.760 125.640 68.690 ;
      LAYER li1 ;
        RECT 126.820 68.630 126.990 68.800 ;
        RECT 127.160 68.630 127.430 68.800 ;
        RECT 127.600 68.630 127.840 68.800 ;
        RECT 128.010 68.630 128.270 68.800 ;
        RECT 128.440 68.630 128.710 68.800 ;
        RECT 128.880 68.630 129.120 68.800 ;
        RECT 129.290 68.630 129.550 68.800 ;
        RECT 131.110 68.790 132.360 68.820 ;
        RECT 133.130 68.790 134.740 68.820 ;
        RECT 126.820 67.830 129.550 68.630 ;
        RECT 121.980 66.500 122.310 67.490 ;
      LAYER li1 ;
        RECT 123.010 67.070 123.310 67.660 ;
        RECT 123.810 67.590 125.640 67.760 ;
        RECT 123.490 67.070 124.680 67.410 ;
      LAYER li1 ;
        RECT 121.210 65.630 122.660 66.500 ;
        RECT 121.210 65.460 121.460 65.630 ;
        RECT 121.630 65.460 121.820 65.630 ;
        RECT 121.990 65.460 122.260 65.630 ;
        RECT 122.430 65.460 122.660 65.630 ;
        RECT 121.210 65.430 122.660 65.460 ;
        RECT 122.970 65.680 124.640 66.890 ;
      LAYER li1 ;
        RECT 124.860 65.930 125.190 67.410 ;
      LAYER li1 ;
        RECT 122.970 65.510 123.000 65.680 ;
        RECT 123.170 65.510 123.360 65.680 ;
        RECT 123.530 65.510 123.720 65.680 ;
        RECT 123.890 65.510 124.080 65.680 ;
        RECT 124.250 65.510 124.440 65.680 ;
        RECT 124.610 65.510 124.640 65.680 ;
        RECT 122.970 65.430 124.640 65.510 ;
      LAYER li1 ;
        RECT 125.370 65.430 125.640 67.590 ;
      LAYER li1 ;
        RECT 126.980 67.160 127.310 67.830 ;
        RECT 127.710 66.510 128.040 67.490 ;
        RECT 128.260 67.160 128.590 67.830 ;
        RECT 128.990 66.510 129.320 67.490 ;
      LAYER li1 ;
        RECT 130.680 67.010 130.930 68.690 ;
      LAYER li1 ;
        RECT 131.280 68.620 131.470 68.790 ;
        RECT 131.640 68.620 131.830 68.790 ;
        RECT 132.000 68.620 132.190 68.790 ;
        RECT 131.110 68.250 132.360 68.620 ;
        RECT 132.540 68.070 132.790 68.690 ;
        RECT 133.130 68.620 133.180 68.790 ;
        RECT 133.350 68.620 133.620 68.790 ;
        RECT 133.790 68.620 134.060 68.790 ;
        RECT 134.230 68.620 134.470 68.790 ;
        RECT 134.640 68.620 134.740 68.790 ;
        RECT 133.130 68.340 134.740 68.620 ;
        RECT 131.240 67.900 132.790 68.070 ;
        RECT 131.240 67.440 131.570 67.900 ;
        RECT 126.740 65.630 129.480 66.510 ;
        RECT 126.740 65.460 126.950 65.630 ;
        RECT 127.120 65.460 127.390 65.630 ;
        RECT 127.560 65.460 127.800 65.630 ;
        RECT 127.970 65.460 128.230 65.630 ;
        RECT 128.400 65.460 128.670 65.630 ;
        RECT 128.840 65.460 129.080 65.630 ;
        RECT 129.250 65.460 129.480 65.630 ;
        RECT 126.740 65.440 129.480 65.460 ;
      LAYER li1 ;
        RECT 130.680 65.430 131.110 67.010 ;
      LAYER li1 ;
        RECT 131.290 65.680 131.850 67.010 ;
      LAYER li1 ;
        RECT 132.030 65.930 132.360 67.720 ;
      LAYER li1 ;
        RECT 132.540 66.180 132.790 67.900 ;
        RECT 133.440 67.940 134.740 68.340 ;
        RECT 134.970 68.790 135.560 68.820 ;
        RECT 134.970 68.620 135.000 68.790 ;
        RECT 135.170 68.620 135.360 68.790 ;
        RECT 135.530 68.620 135.560 68.790 ;
        RECT 136.900 68.800 139.630 68.830 ;
        RECT 133.440 67.160 133.770 67.940 ;
        RECT 134.970 67.860 135.560 68.620 ;
        RECT 133.980 66.500 134.310 67.490 ;
      LAYER li1 ;
        RECT 135.010 67.250 135.720 67.640 ;
        RECT 135.900 67.010 136.230 68.690 ;
      LAYER li1 ;
        RECT 136.900 68.630 137.070 68.800 ;
        RECT 137.240 68.630 137.510 68.800 ;
        RECT 137.680 68.630 137.920 68.800 ;
        RECT 138.090 68.630 138.350 68.800 ;
        RECT 138.520 68.630 138.790 68.800 ;
        RECT 138.960 68.630 139.200 68.800 ;
        RECT 139.370 68.630 139.630 68.800 ;
        RECT 136.900 67.830 139.630 68.630 ;
        RECT 140.330 68.790 141.940 68.820 ;
        RECT 140.330 68.620 140.380 68.790 ;
        RECT 140.550 68.620 140.820 68.790 ;
        RECT 140.990 68.620 141.260 68.790 ;
        RECT 141.430 68.620 141.670 68.790 ;
        RECT 141.840 68.620 141.940 68.790 ;
        RECT 140.330 68.340 141.940 68.620 ;
        RECT 140.640 67.940 141.940 68.340 ;
        RECT 137.060 67.160 137.390 67.830 ;
        RECT 131.290 65.510 131.300 65.680 ;
        RECT 131.470 65.510 131.660 65.680 ;
        RECT 131.830 65.510 131.850 65.680 ;
        RECT 131.290 65.430 131.850 65.510 ;
        RECT 133.210 65.630 134.660 66.500 ;
        RECT 133.210 65.460 133.460 65.630 ;
        RECT 133.630 65.460 133.820 65.630 ;
        RECT 133.990 65.460 134.260 65.630 ;
        RECT 134.430 65.460 134.660 65.630 ;
        RECT 133.210 65.430 134.660 65.460 ;
        RECT 134.970 65.680 135.560 67.010 ;
        RECT 134.970 65.510 135.000 65.680 ;
        RECT 135.170 65.510 135.360 65.680 ;
        RECT 135.530 65.510 135.560 65.680 ;
        RECT 134.970 65.430 135.560 65.510 ;
      LAYER li1 ;
        RECT 135.840 65.430 136.230 67.010 ;
      LAYER li1 ;
        RECT 137.790 66.510 138.120 67.490 ;
        RECT 138.340 67.160 138.670 67.830 ;
        RECT 139.070 66.510 139.400 67.490 ;
        RECT 140.640 67.160 140.970 67.940 ;
        RECT 136.820 65.630 139.560 66.510 ;
        RECT 141.180 66.500 141.510 67.490 ;
        RECT 136.820 65.460 137.030 65.630 ;
        RECT 137.200 65.460 137.470 65.630 ;
        RECT 137.640 65.460 137.880 65.630 ;
        RECT 138.050 65.460 138.310 65.630 ;
        RECT 138.480 65.460 138.750 65.630 ;
        RECT 138.920 65.460 139.160 65.630 ;
        RECT 139.330 65.460 139.560 65.630 ;
        RECT 136.820 65.440 139.560 65.460 ;
        RECT 140.410 65.630 141.860 66.500 ;
        RECT 140.410 65.460 140.660 65.630 ;
        RECT 140.830 65.460 141.020 65.630 ;
        RECT 141.190 65.460 141.460 65.630 ;
        RECT 141.630 65.460 141.860 65.630 ;
        RECT 140.410 65.430 141.860 65.460 ;
        RECT 5.760 65.030 5.920 65.210 ;
        RECT 6.090 65.030 6.400 65.210 ;
        RECT 6.570 65.030 6.880 65.210 ;
        RECT 7.050 65.030 7.360 65.210 ;
        RECT 7.530 65.030 7.840 65.210 ;
        RECT 8.010 65.030 8.320 65.210 ;
        RECT 8.490 65.200 8.800 65.210 ;
        RECT 8.970 65.200 9.280 65.210 ;
        RECT 8.490 65.030 8.640 65.200 ;
        RECT 9.120 65.030 9.280 65.200 ;
        RECT 9.450 65.030 9.760 65.210 ;
        RECT 9.930 65.030 10.240 65.210 ;
        RECT 10.410 65.030 10.720 65.210 ;
        RECT 10.890 65.030 11.200 65.210 ;
        RECT 11.370 65.030 11.680 65.210 ;
        RECT 11.850 65.030 12.160 65.210 ;
        RECT 12.330 65.030 12.640 65.210 ;
        RECT 12.810 65.030 13.120 65.210 ;
        RECT 13.290 65.030 13.600 65.210 ;
        RECT 13.770 65.030 14.080 65.210 ;
        RECT 14.250 65.030 14.560 65.210 ;
        RECT 14.730 65.030 15.040 65.210 ;
        RECT 15.210 65.030 15.520 65.210 ;
        RECT 15.690 65.030 16.000 65.210 ;
        RECT 16.170 65.030 16.480 65.210 ;
        RECT 16.650 65.030 16.960 65.210 ;
        RECT 17.130 65.030 17.440 65.210 ;
        RECT 17.610 65.030 17.920 65.210 ;
        RECT 18.090 65.030 18.400 65.210 ;
        RECT 18.570 65.030 18.880 65.210 ;
        RECT 19.050 65.030 19.360 65.210 ;
        RECT 19.530 65.030 19.840 65.210 ;
        RECT 20.010 65.030 20.320 65.210 ;
        RECT 20.490 65.030 20.800 65.210 ;
        RECT 20.970 65.030 21.280 65.210 ;
        RECT 21.450 65.030 21.760 65.210 ;
        RECT 21.930 65.030 22.240 65.210 ;
        RECT 22.410 65.030 22.720 65.210 ;
        RECT 22.890 65.030 23.200 65.210 ;
        RECT 23.370 65.030 23.680 65.210 ;
        RECT 23.850 65.030 24.160 65.210 ;
        RECT 24.330 65.030 24.640 65.210 ;
        RECT 24.810 65.030 25.120 65.210 ;
        RECT 25.290 65.030 25.600 65.210 ;
        RECT 25.770 65.030 26.080 65.210 ;
        RECT 26.250 65.030 26.560 65.210 ;
        RECT 26.730 65.030 27.040 65.210 ;
        RECT 27.210 65.030 27.520 65.210 ;
        RECT 27.690 65.030 28.000 65.210 ;
        RECT 28.170 65.030 28.480 65.210 ;
        RECT 28.650 65.030 28.960 65.210 ;
        RECT 29.130 65.030 29.440 65.210 ;
        RECT 29.610 65.030 29.920 65.210 ;
        RECT 30.090 65.030 30.400 65.210 ;
        RECT 30.570 65.030 30.880 65.210 ;
        RECT 31.050 65.030 31.360 65.210 ;
        RECT 31.530 65.030 31.840 65.210 ;
        RECT 32.010 65.030 32.320 65.210 ;
        RECT 32.490 65.030 32.800 65.210 ;
        RECT 32.970 65.030 33.280 65.210 ;
        RECT 33.450 65.030 33.760 65.210 ;
        RECT 33.930 65.030 34.240 65.210 ;
        RECT 34.410 65.030 34.720 65.210 ;
        RECT 34.890 65.030 35.200 65.210 ;
        RECT 35.370 65.030 35.680 65.210 ;
        RECT 35.850 65.030 36.160 65.210 ;
        RECT 36.330 65.030 36.640 65.210 ;
        RECT 36.810 65.030 37.120 65.210 ;
        RECT 37.290 65.030 37.600 65.210 ;
        RECT 37.770 65.030 38.080 65.210 ;
        RECT 38.250 65.030 38.560 65.210 ;
        RECT 38.730 65.030 39.040 65.210 ;
        RECT 39.210 65.030 39.520 65.210 ;
        RECT 39.690 65.030 40.000 65.210 ;
        RECT 40.170 65.030 40.480 65.210 ;
        RECT 40.650 65.030 40.960 65.210 ;
        RECT 41.130 65.030 41.440 65.210 ;
        RECT 41.610 65.030 41.920 65.210 ;
        RECT 42.090 65.030 42.400 65.210 ;
        RECT 42.570 65.030 42.880 65.210 ;
        RECT 43.050 65.030 43.360 65.210 ;
        RECT 43.530 65.030 43.840 65.210 ;
        RECT 44.010 65.030 44.320 65.210 ;
        RECT 44.490 65.030 44.800 65.210 ;
        RECT 44.970 65.030 45.280 65.210 ;
        RECT 45.450 65.030 45.760 65.210 ;
        RECT 45.930 65.030 46.240 65.210 ;
        RECT 46.410 65.030 46.720 65.210 ;
        RECT 46.890 65.030 47.200 65.210 ;
        RECT 47.370 65.200 47.680 65.210 ;
        RECT 47.850 65.200 48.160 65.210 ;
        RECT 47.370 65.030 47.520 65.200 ;
        RECT 48.000 65.030 48.160 65.200 ;
        RECT 48.330 65.030 48.640 65.210 ;
        RECT 48.810 65.030 49.120 65.210 ;
        RECT 49.290 65.030 49.600 65.210 ;
        RECT 49.770 65.030 50.080 65.210 ;
        RECT 50.250 65.030 50.560 65.210 ;
        RECT 50.730 65.030 51.040 65.210 ;
        RECT 51.210 65.030 51.520 65.210 ;
        RECT 51.690 65.030 52.000 65.210 ;
        RECT 52.170 65.030 52.480 65.210 ;
        RECT 52.650 65.030 52.960 65.210 ;
        RECT 53.130 65.030 53.440 65.210 ;
        RECT 53.610 65.030 53.920 65.210 ;
        RECT 54.090 65.030 54.400 65.210 ;
        RECT 54.570 65.030 54.880 65.210 ;
        RECT 55.050 65.030 55.360 65.210 ;
        RECT 55.530 65.030 55.840 65.210 ;
        RECT 56.010 65.030 56.320 65.210 ;
        RECT 56.490 65.030 56.800 65.210 ;
        RECT 56.970 65.030 57.280 65.210 ;
        RECT 57.450 65.030 57.760 65.210 ;
        RECT 57.930 65.030 58.240 65.210 ;
        RECT 58.410 65.030 58.720 65.210 ;
        RECT 58.890 65.030 59.200 65.210 ;
        RECT 59.370 65.030 59.680 65.210 ;
        RECT 59.850 65.030 60.160 65.210 ;
        RECT 60.330 65.030 60.640 65.210 ;
        RECT 60.810 65.030 61.120 65.210 ;
        RECT 61.290 65.030 61.600 65.210 ;
        RECT 61.770 65.030 62.080 65.210 ;
        RECT 62.250 65.030 62.560 65.210 ;
        RECT 62.730 65.030 63.040 65.210 ;
        RECT 63.210 65.030 63.520 65.210 ;
        RECT 63.690 65.030 64.000 65.210 ;
        RECT 64.170 65.030 64.480 65.210 ;
        RECT 64.650 65.030 64.960 65.210 ;
        RECT 65.130 65.030 65.440 65.210 ;
        RECT 65.610 65.030 65.920 65.210 ;
        RECT 66.090 65.030 66.400 65.210 ;
        RECT 66.570 65.030 66.880 65.210 ;
        RECT 67.050 65.030 67.360 65.210 ;
        RECT 67.530 65.030 67.840 65.210 ;
        RECT 68.010 65.030 68.320 65.210 ;
        RECT 68.490 65.030 68.800 65.210 ;
        RECT 68.970 65.030 69.280 65.210 ;
        RECT 69.450 65.030 69.760 65.210 ;
        RECT 69.930 65.030 70.240 65.210 ;
        RECT 70.410 65.030 70.720 65.210 ;
        RECT 70.890 65.030 71.200 65.210 ;
        RECT 71.370 65.030 71.680 65.210 ;
        RECT 71.850 65.030 72.160 65.210 ;
        RECT 72.330 65.030 72.640 65.210 ;
        RECT 72.810 65.030 73.120 65.210 ;
        RECT 73.290 65.030 73.600 65.210 ;
        RECT 73.770 65.030 74.080 65.210 ;
        RECT 74.250 65.030 74.560 65.210 ;
        RECT 74.730 65.030 75.040 65.210 ;
        RECT 75.210 65.030 75.520 65.210 ;
        RECT 75.690 65.030 76.000 65.210 ;
        RECT 76.170 65.030 76.480 65.210 ;
        RECT 76.650 65.030 76.960 65.210 ;
        RECT 77.130 65.030 77.440 65.210 ;
        RECT 77.610 65.030 77.920 65.210 ;
        RECT 78.090 65.030 78.400 65.210 ;
        RECT 78.570 65.030 78.880 65.210 ;
        RECT 79.050 65.030 79.360 65.210 ;
        RECT 79.530 65.030 79.840 65.210 ;
        RECT 80.010 65.030 80.320 65.210 ;
        RECT 80.490 65.030 80.800 65.210 ;
        RECT 80.970 65.030 81.280 65.210 ;
        RECT 81.450 65.030 81.760 65.210 ;
        RECT 81.930 65.030 82.240 65.210 ;
        RECT 82.410 65.030 82.720 65.210 ;
        RECT 82.890 65.030 83.200 65.210 ;
        RECT 83.370 65.030 83.680 65.210 ;
        RECT 83.850 65.030 84.160 65.210 ;
        RECT 84.330 65.030 84.640 65.210 ;
        RECT 84.810 65.030 85.120 65.210 ;
        RECT 85.290 65.030 85.600 65.210 ;
        RECT 85.770 65.030 86.080 65.210 ;
        RECT 86.250 65.030 86.560 65.210 ;
        RECT 86.730 65.030 87.040 65.210 ;
        RECT 87.210 65.030 87.520 65.210 ;
        RECT 87.690 65.030 88.000 65.210 ;
        RECT 88.170 65.030 88.480 65.210 ;
        RECT 88.650 65.030 88.960 65.210 ;
        RECT 89.130 65.030 89.440 65.210 ;
        RECT 89.610 65.030 89.920 65.210 ;
        RECT 90.090 65.030 90.400 65.210 ;
        RECT 90.570 65.030 90.880 65.210 ;
        RECT 91.050 65.030 91.200 65.210 ;
        RECT 91.680 65.030 91.840 65.210 ;
        RECT 92.010 65.030 92.320 65.210 ;
        RECT 92.490 65.030 92.800 65.210 ;
        RECT 92.970 65.030 93.280 65.210 ;
        RECT 93.450 65.030 93.760 65.210 ;
        RECT 93.930 65.030 94.240 65.210 ;
        RECT 94.410 65.030 94.720 65.210 ;
        RECT 94.890 65.030 95.200 65.210 ;
        RECT 95.370 65.030 95.680 65.210 ;
        RECT 95.850 65.030 96.160 65.210 ;
        RECT 96.330 65.030 96.640 65.210 ;
        RECT 96.810 65.030 97.120 65.210 ;
        RECT 97.290 65.030 97.600 65.210 ;
        RECT 97.770 65.030 98.080 65.210 ;
        RECT 98.250 65.030 98.560 65.210 ;
        RECT 98.730 65.030 99.040 65.210 ;
        RECT 99.210 65.030 99.520 65.210 ;
        RECT 99.690 65.030 100.000 65.210 ;
        RECT 100.170 65.030 100.480 65.210 ;
        RECT 100.650 65.030 100.960 65.210 ;
        RECT 101.130 65.030 101.440 65.210 ;
        RECT 101.610 65.030 101.920 65.210 ;
        RECT 102.090 65.030 102.400 65.210 ;
        RECT 102.570 65.030 102.880 65.210 ;
        RECT 103.050 65.030 103.360 65.210 ;
        RECT 103.530 65.030 103.840 65.210 ;
        RECT 104.010 65.030 104.320 65.210 ;
        RECT 104.490 65.030 104.800 65.210 ;
        RECT 104.970 65.030 105.280 65.210 ;
        RECT 105.450 65.200 105.600 65.210 ;
        RECT 106.080 65.200 106.240 65.210 ;
        RECT 105.450 65.030 105.760 65.200 ;
        RECT 105.930 65.030 106.240 65.200 ;
        RECT 106.410 65.030 106.720 65.210 ;
        RECT 106.890 65.030 107.200 65.210 ;
        RECT 107.370 65.030 107.680 65.210 ;
        RECT 107.850 65.030 108.160 65.210 ;
        RECT 108.330 65.030 108.640 65.210 ;
        RECT 108.810 65.030 109.120 65.210 ;
        RECT 109.290 65.030 109.600 65.210 ;
        RECT 109.770 65.030 110.080 65.210 ;
        RECT 110.250 65.030 110.560 65.210 ;
        RECT 110.730 65.030 111.040 65.210 ;
        RECT 111.210 65.030 111.520 65.210 ;
        RECT 111.690 65.030 112.000 65.210 ;
        RECT 112.170 65.030 112.480 65.210 ;
        RECT 112.650 65.030 112.960 65.210 ;
        RECT 113.130 65.030 113.440 65.210 ;
        RECT 113.610 65.030 113.920 65.210 ;
        RECT 114.090 65.030 114.400 65.210 ;
        RECT 114.570 65.030 114.880 65.210 ;
        RECT 115.050 65.030 115.360 65.210 ;
        RECT 115.530 65.030 115.840 65.210 ;
        RECT 116.010 65.030 116.320 65.210 ;
        RECT 116.490 65.030 116.800 65.210 ;
        RECT 116.970 65.030 117.280 65.210 ;
        RECT 117.450 65.030 117.760 65.210 ;
        RECT 117.930 65.030 118.240 65.210 ;
        RECT 118.410 65.030 118.720 65.210 ;
        RECT 118.890 65.030 119.200 65.210 ;
        RECT 119.370 65.030 119.680 65.210 ;
        RECT 119.850 65.030 120.160 65.210 ;
        RECT 120.330 65.030 120.640 65.210 ;
        RECT 120.810 65.030 121.120 65.210 ;
        RECT 121.290 65.030 121.600 65.210 ;
        RECT 121.770 65.030 122.080 65.210 ;
        RECT 122.250 65.030 122.560 65.210 ;
        RECT 122.730 65.030 123.040 65.210 ;
        RECT 123.210 65.030 123.520 65.210 ;
        RECT 123.690 65.030 124.000 65.210 ;
        RECT 124.170 65.030 124.480 65.210 ;
        RECT 124.650 65.030 124.960 65.210 ;
        RECT 125.130 65.030 125.440 65.210 ;
        RECT 125.610 65.030 125.920 65.210 ;
        RECT 126.090 65.030 126.400 65.210 ;
        RECT 126.570 65.030 126.880 65.210 ;
        RECT 127.050 65.030 127.360 65.210 ;
        RECT 127.530 65.030 127.840 65.210 ;
        RECT 128.010 65.030 128.320 65.210 ;
        RECT 128.490 65.030 128.800 65.210 ;
        RECT 128.970 65.030 129.280 65.210 ;
        RECT 129.450 65.030 129.760 65.210 ;
        RECT 129.930 65.200 130.240 65.210 ;
        RECT 130.410 65.200 130.720 65.210 ;
        RECT 129.930 65.030 130.080 65.200 ;
        RECT 130.560 65.030 130.720 65.200 ;
        RECT 130.890 65.030 131.200 65.210 ;
        RECT 131.370 65.030 131.680 65.210 ;
        RECT 131.850 65.030 132.160 65.210 ;
        RECT 132.330 65.030 132.640 65.210 ;
        RECT 132.810 65.030 133.120 65.210 ;
        RECT 133.290 65.030 133.600 65.210 ;
        RECT 133.770 65.030 134.080 65.210 ;
        RECT 134.250 65.030 134.560 65.210 ;
        RECT 134.730 65.030 135.040 65.210 ;
        RECT 135.210 65.030 135.520 65.210 ;
        RECT 135.690 65.030 136.000 65.210 ;
        RECT 136.170 65.030 136.480 65.210 ;
        RECT 136.650 65.030 136.960 65.210 ;
        RECT 137.130 65.030 137.440 65.210 ;
        RECT 137.610 65.030 137.920 65.210 ;
        RECT 138.090 65.030 138.400 65.210 ;
        RECT 138.570 65.030 138.880 65.210 ;
        RECT 139.050 65.030 139.360 65.210 ;
        RECT 139.530 65.030 139.840 65.210 ;
        RECT 140.010 65.030 140.320 65.210 ;
        RECT 140.490 65.030 140.800 65.210 ;
        RECT 140.970 65.030 141.280 65.210 ;
        RECT 141.450 65.200 141.600 65.210 ;
        RECT 141.450 65.030 141.760 65.200 ;
        RECT 141.930 65.030 142.080 65.200 ;
        RECT 6.010 64.780 7.460 64.810 ;
        RECT 6.010 64.610 6.260 64.780 ;
        RECT 6.430 64.610 6.620 64.780 ;
        RECT 6.790 64.610 7.060 64.780 ;
        RECT 7.230 64.610 7.460 64.780 ;
        RECT 6.010 63.740 7.460 64.610 ;
        RECT 7.770 64.730 9.440 64.810 ;
        RECT 7.770 64.560 7.800 64.730 ;
        RECT 7.970 64.560 8.160 64.730 ;
        RECT 8.330 64.560 8.520 64.730 ;
        RECT 8.690 64.560 8.880 64.730 ;
        RECT 9.050 64.560 9.240 64.730 ;
        RECT 9.410 64.560 9.440 64.730 ;
        RECT 6.240 62.300 6.570 63.080 ;
        RECT 6.780 62.750 7.110 63.740 ;
        RECT 7.770 63.350 9.440 64.560 ;
      LAYER li1 ;
        RECT 7.810 62.830 9.000 63.170 ;
        RECT 9.180 62.830 9.510 63.170 ;
        RECT 9.700 62.650 9.960 64.810 ;
      LAYER li1 ;
        RECT 10.330 64.780 11.780 64.810 ;
        RECT 10.330 64.610 10.580 64.780 ;
        RECT 10.750 64.610 10.940 64.780 ;
        RECT 11.110 64.610 11.380 64.780 ;
        RECT 11.550 64.610 11.780 64.780 ;
        RECT 10.330 63.740 11.780 64.610 ;
        RECT 12.090 64.730 13.040 64.810 ;
        RECT 12.090 64.560 12.120 64.730 ;
        RECT 12.290 64.560 12.480 64.730 ;
        RECT 12.650 64.560 12.840 64.730 ;
        RECT 13.010 64.560 13.040 64.730 ;
      LAYER li1 ;
        RECT 8.880 62.480 9.960 62.650 ;
      LAYER li1 ;
        RECT 6.240 61.900 7.540 62.300 ;
        RECT 5.930 61.420 7.540 61.900 ;
        RECT 7.770 61.420 8.700 62.380 ;
      LAYER li1 ;
        RECT 8.880 61.550 9.210 62.480 ;
      LAYER li1 ;
        RECT 10.560 62.300 10.890 63.080 ;
        RECT 11.100 62.750 11.430 63.740 ;
        RECT 12.090 63.230 13.040 64.560 ;
      LAYER li1 ;
        RECT 12.130 62.600 13.020 62.990 ;
        RECT 13.220 62.750 13.470 64.810 ;
      LAYER li1 ;
        RECT 13.660 64.730 14.250 64.810 ;
        RECT 13.660 64.560 13.690 64.730 ;
        RECT 13.860 64.560 14.050 64.730 ;
        RECT 14.220 64.560 14.250 64.730 ;
        RECT 13.660 63.230 14.250 64.560 ;
        RECT 14.650 64.780 16.100 64.810 ;
        RECT 14.650 64.610 14.900 64.780 ;
        RECT 15.070 64.610 15.260 64.780 ;
        RECT 15.430 64.610 15.700 64.780 ;
        RECT 15.870 64.610 16.100 64.780 ;
        RECT 14.650 63.740 16.100 64.610 ;
      LAYER li1 ;
        RECT 13.220 62.580 13.800 62.750 ;
        RECT 13.980 62.580 14.280 62.910 ;
        RECT 13.580 62.400 13.800 62.580 ;
      LAYER li1 ;
        RECT 9.400 61.420 9.990 62.300 ;
        RECT 10.560 61.900 11.860 62.300 ;
        RECT 10.250 61.420 11.860 61.900 ;
        RECT 12.090 61.420 13.400 62.400 ;
      LAYER li1 ;
        RECT 13.580 62.230 14.180 62.400 ;
        RECT 13.850 61.570 14.180 62.230 ;
      LAYER li1 ;
        RECT 14.880 62.300 15.210 63.080 ;
        RECT 15.420 62.750 15.750 63.740 ;
        RECT 16.580 63.150 16.830 64.810 ;
        RECT 17.010 64.730 18.260 64.810 ;
        RECT 17.180 64.560 17.370 64.730 ;
        RECT 17.540 64.560 17.730 64.730 ;
        RECT 17.900 64.560 18.090 64.730 ;
        RECT 17.010 63.330 18.260 64.560 ;
        RECT 18.440 63.150 18.610 64.810 ;
        RECT 16.580 62.980 18.610 63.150 ;
      LAYER li1 ;
        RECT 18.790 62.860 19.120 64.310 ;
        RECT 16.450 62.560 17.640 62.800 ;
        RECT 17.890 62.560 18.240 62.800 ;
        RECT 19.300 62.680 19.560 64.810 ;
      LAYER li1 ;
        RECT 19.930 64.780 21.380 64.810 ;
        RECT 19.930 64.610 20.180 64.780 ;
        RECT 20.350 64.610 20.540 64.780 ;
        RECT 20.710 64.610 20.980 64.780 ;
        RECT 21.150 64.610 21.380 64.780 ;
        RECT 19.930 63.740 21.380 64.610 ;
        RECT 22.230 64.730 22.820 64.760 ;
        RECT 22.230 64.560 22.260 64.730 ;
        RECT 22.430 64.560 22.620 64.730 ;
        RECT 22.790 64.560 22.820 64.730 ;
      LAYER li1 ;
        RECT 18.540 62.510 19.560 62.680 ;
      LAYER li1 ;
        RECT 14.880 61.900 16.180 62.300 ;
        RECT 14.570 61.420 16.180 61.900 ;
        RECT 16.650 61.420 18.360 62.380 ;
      LAYER li1 ;
        RECT 18.540 61.550 18.790 62.510 ;
      LAYER li1 ;
        RECT 19.000 61.420 19.590 62.330 ;
        RECT 20.160 62.300 20.490 63.080 ;
        RECT 20.700 62.750 21.030 63.740 ;
        RECT 21.710 63.580 22.040 64.510 ;
        RECT 22.230 63.780 22.820 64.560 ;
        RECT 23.000 64.690 24.440 64.860 ;
        RECT 23.000 63.580 23.170 64.690 ;
        RECT 21.710 63.410 23.170 63.580 ;
        RECT 20.160 61.900 21.460 62.300 ;
        RECT 19.850 61.420 21.460 61.900 ;
        RECT 21.710 61.550 21.980 63.410 ;
        RECT 22.840 62.910 23.170 63.410 ;
        RECT 23.350 63.200 23.600 64.510 ;
        RECT 23.840 63.890 24.090 64.510 ;
        RECT 24.270 64.240 24.440 64.690 ;
        RECT 24.620 64.730 24.950 64.760 ;
        RECT 24.620 64.560 24.650 64.730 ;
        RECT 24.820 64.560 24.950 64.730 ;
        RECT 24.620 64.420 24.950 64.560 ;
        RECT 25.130 64.690 26.870 64.860 ;
        RECT 25.130 64.240 25.300 64.690 ;
        RECT 24.270 64.070 25.300 64.240 ;
        RECT 25.480 63.890 25.650 64.510 ;
        RECT 26.180 64.250 26.510 64.510 ;
        RECT 23.840 63.720 25.650 63.890 ;
        RECT 25.830 63.720 26.050 64.050 ;
        RECT 25.480 63.540 25.650 63.720 ;
        RECT 23.350 62.970 23.880 63.200 ;
        RECT 23.350 62.050 23.620 62.970 ;
      LAYER li1 ;
        RECT 24.300 62.670 24.840 63.540 ;
      LAYER li1 ;
        RECT 25.480 63.370 25.700 63.540 ;
        RECT 22.160 61.420 23.110 62.050 ;
        RECT 23.290 61.550 23.620 62.050 ;
        RECT 23.800 61.420 24.390 62.300 ;
      LAYER li1 ;
        RECT 24.670 61.680 24.840 62.670 ;
        RECT 25.020 61.860 25.350 63.160 ;
      LAYER li1 ;
        RECT 25.530 62.380 25.700 63.370 ;
        RECT 25.880 63.200 26.050 63.720 ;
        RECT 26.230 63.550 26.400 64.250 ;
        RECT 26.700 64.100 26.870 64.690 ;
        RECT 27.050 64.730 28.000 64.760 ;
        RECT 27.050 64.560 27.080 64.730 ;
        RECT 27.250 64.560 27.440 64.730 ;
        RECT 27.610 64.560 27.800 64.730 ;
        RECT 27.970 64.560 28.000 64.730 ;
        RECT 27.050 64.280 28.000 64.560 ;
        RECT 28.180 64.690 29.210 64.860 ;
        RECT 28.180 64.100 28.350 64.690 ;
        RECT 26.700 64.050 28.350 64.100 ;
        RECT 26.580 63.930 28.350 64.050 ;
        RECT 26.580 63.730 26.910 63.930 ;
        RECT 28.530 63.750 28.860 64.510 ;
        RECT 29.040 64.330 29.210 64.690 ;
        RECT 29.390 64.730 30.340 64.810 ;
        RECT 29.390 64.560 29.420 64.730 ;
        RECT 29.590 64.560 29.780 64.730 ;
        RECT 29.950 64.560 30.140 64.730 ;
        RECT 30.310 64.560 30.340 64.730 ;
        RECT 29.390 64.510 30.340 64.560 ;
        RECT 29.040 64.160 30.850 64.330 ;
        RECT 27.090 63.580 28.860 63.750 ;
        RECT 27.090 63.550 27.260 63.580 ;
        RECT 26.230 63.380 27.260 63.550 ;
        RECT 30.170 63.400 30.500 63.980 ;
        RECT 25.880 62.970 26.910 63.200 ;
        RECT 26.580 62.480 26.910 62.970 ;
        RECT 27.090 62.700 27.260 63.380 ;
        RECT 27.440 63.230 30.500 63.400 ;
        RECT 27.440 62.880 27.770 63.230 ;
      LAYER li1 ;
        RECT 28.210 62.880 30.060 63.050 ;
      LAYER li1 ;
        RECT 27.090 62.530 29.710 62.700 ;
        RECT 25.530 61.880 25.800 62.380 ;
        RECT 27.090 62.300 27.260 62.530 ;
      LAYER li1 ;
        RECT 29.890 62.350 30.060 62.880 ;
      LAYER li1 ;
        RECT 26.250 62.130 27.260 62.300 ;
      LAYER li1 ;
        RECT 27.440 62.180 30.060 62.350 ;
      LAYER li1 ;
        RECT 26.250 61.880 26.580 62.130 ;
      LAYER li1 ;
        RECT 27.440 61.680 27.610 62.180 ;
        RECT 24.670 61.510 27.610 61.680 ;
      LAYER li1 ;
        RECT 28.760 61.420 29.710 62.000 ;
      LAYER li1 ;
        RECT 29.890 61.490 30.060 62.180 ;
      LAYER li1 ;
        RECT 30.240 62.380 30.500 63.230 ;
        RECT 30.680 62.810 30.850 64.160 ;
        RECT 31.030 63.900 31.280 64.810 ;
        RECT 32.090 64.730 33.040 64.760 ;
        RECT 33.870 64.730 34.770 64.760 ;
        RECT 32.090 64.560 32.120 64.730 ;
        RECT 32.290 64.560 32.480 64.730 ;
        RECT 32.650 64.560 32.840 64.730 ;
        RECT 33.010 64.560 33.040 64.730 ;
        RECT 34.040 64.560 34.230 64.730 ;
        RECT 34.400 64.560 34.590 64.730 ;
        RECT 34.760 64.560 34.770 64.730 ;
        RECT 31.030 63.730 31.910 63.900 ;
        RECT 32.090 63.730 33.040 64.560 ;
        RECT 33.440 63.760 33.690 64.230 ;
        RECT 33.870 63.940 34.770 64.560 ;
        RECT 35.380 64.730 36.320 64.790 ;
        RECT 35.380 64.560 35.400 64.730 ;
        RECT 35.570 64.560 35.760 64.730 ;
        RECT 35.930 64.560 36.120 64.730 ;
        RECT 36.290 64.560 36.320 64.730 ;
        RECT 31.230 62.990 31.560 63.490 ;
        RECT 31.740 63.410 31.910 63.730 ;
        RECT 33.440 63.590 34.450 63.760 ;
        RECT 31.740 63.240 34.100 63.410 ;
        RECT 30.680 62.640 31.850 62.810 ;
        RECT 30.240 61.670 30.570 62.380 ;
        RECT 31.030 61.840 31.360 62.380 ;
        RECT 31.570 62.140 31.850 62.640 ;
        RECT 32.030 61.840 32.200 63.240 ;
        RECT 34.280 63.060 34.450 63.590 ;
        RECT 32.410 62.890 34.450 63.060 ;
        RECT 32.410 62.500 32.740 62.890 ;
      LAYER li1 ;
        RECT 33.060 62.320 33.390 62.710 ;
      LAYER li1 ;
        RECT 31.030 61.670 32.200 61.840 ;
      LAYER li1 ;
        RECT 32.380 62.150 33.390 62.320 ;
        RECT 32.380 61.490 32.550 62.150 ;
      LAYER li1 ;
        RECT 34.220 62.050 34.450 62.890 ;
        RECT 34.950 63.060 35.200 64.060 ;
        RECT 35.380 63.250 36.320 64.560 ;
        RECT 34.950 62.730 36.320 63.060 ;
        RECT 34.950 62.550 35.160 62.730 ;
        RECT 34.830 62.050 35.160 62.550 ;
      LAYER li1 ;
        RECT 29.890 61.320 32.550 61.490 ;
      LAYER li1 ;
        RECT 32.730 61.420 33.680 61.970 ;
        RECT 34.220 61.550 34.550 62.050 ;
        RECT 35.340 61.420 36.290 62.550 ;
      LAYER li1 ;
        RECT 36.500 61.720 36.840 64.790 ;
      LAYER li1 ;
        RECT 37.210 64.780 38.660 64.810 ;
        RECT 37.210 64.610 37.460 64.780 ;
        RECT 37.630 64.610 37.820 64.780 ;
        RECT 37.990 64.610 38.260 64.780 ;
        RECT 38.430 64.610 38.660 64.780 ;
        RECT 37.210 63.740 38.660 64.610 ;
        RECT 38.970 64.730 39.920 64.810 ;
        RECT 38.970 64.560 39.000 64.730 ;
        RECT 39.170 64.560 39.360 64.730 ;
        RECT 39.530 64.560 39.720 64.730 ;
        RECT 39.890 64.560 39.920 64.730 ;
        RECT 37.440 62.300 37.770 63.080 ;
        RECT 37.980 62.750 38.310 63.740 ;
        RECT 38.970 63.230 39.920 64.560 ;
      LAYER li1 ;
        RECT 40.100 63.130 40.350 64.810 ;
      LAYER li1 ;
        RECT 40.530 64.730 41.480 64.810 ;
        RECT 40.530 64.560 40.560 64.730 ;
        RECT 40.730 64.560 40.920 64.730 ;
        RECT 41.090 64.560 41.280 64.730 ;
        RECT 41.450 64.560 41.480 64.730 ;
        RECT 40.530 63.310 41.480 64.560 ;
      LAYER li1 ;
        RECT 41.660 63.130 41.990 64.810 ;
      LAYER li1 ;
        RECT 42.170 64.730 43.120 64.810 ;
        RECT 42.170 64.560 42.200 64.730 ;
        RECT 42.370 64.560 42.560 64.730 ;
        RECT 42.730 64.560 42.920 64.730 ;
        RECT 43.090 64.560 43.120 64.730 ;
        RECT 42.170 63.350 43.120 64.560 ;
      LAYER li1 ;
        RECT 40.100 62.960 41.990 63.130 ;
        RECT 40.100 62.830 40.270 62.960 ;
        RECT 42.770 62.830 43.100 63.170 ;
        RECT 39.010 62.600 40.270 62.830 ;
      LAYER li1 ;
        RECT 40.450 62.650 42.480 62.780 ;
        RECT 43.300 62.650 43.550 64.810 ;
        RECT 43.930 64.780 45.380 64.810 ;
        RECT 43.930 64.610 44.180 64.780 ;
        RECT 44.350 64.610 44.540 64.780 ;
        RECT 44.710 64.610 44.980 64.780 ;
        RECT 45.150 64.610 45.380 64.780 ;
        RECT 43.930 63.740 45.380 64.610 ;
        RECT 47.190 64.730 47.780 64.760 ;
        RECT 47.190 64.560 47.220 64.730 ;
        RECT 47.390 64.560 47.580 64.730 ;
        RECT 47.750 64.560 47.780 64.730 ;
        RECT 40.450 62.610 43.550 62.650 ;
      LAYER li1 ;
        RECT 40.100 62.430 40.270 62.600 ;
      LAYER li1 ;
        RECT 42.310 62.480 43.550 62.610 ;
        RECT 37.440 61.900 38.740 62.300 ;
        RECT 37.130 61.420 38.740 61.900 ;
        RECT 38.970 61.420 39.920 62.380 ;
      LAYER li1 ;
        RECT 40.100 62.260 41.910 62.430 ;
        RECT 40.100 61.550 40.350 62.260 ;
      LAYER li1 ;
        RECT 40.530 61.420 41.480 62.080 ;
      LAYER li1 ;
        RECT 41.660 61.550 41.910 62.260 ;
      LAYER li1 ;
        RECT 42.090 61.420 43.040 62.300 ;
        RECT 43.220 61.550 43.550 62.480 ;
        RECT 44.160 62.300 44.490 63.080 ;
        RECT 44.700 62.750 45.030 63.740 ;
        RECT 46.670 63.580 47.000 64.510 ;
        RECT 47.190 63.780 47.780 64.560 ;
        RECT 47.960 64.690 49.400 64.860 ;
        RECT 47.960 63.580 48.130 64.690 ;
        RECT 46.670 63.410 48.130 63.580 ;
        RECT 44.160 61.900 45.460 62.300 ;
        RECT 43.850 61.420 45.460 61.900 ;
        RECT 46.670 61.550 46.940 63.410 ;
        RECT 47.800 62.910 48.130 63.410 ;
        RECT 48.310 63.200 48.560 64.510 ;
        RECT 48.800 63.890 49.050 64.510 ;
        RECT 49.230 64.240 49.400 64.690 ;
        RECT 49.580 64.730 49.910 64.760 ;
        RECT 49.580 64.560 49.610 64.730 ;
        RECT 49.780 64.560 49.910 64.730 ;
        RECT 49.580 64.420 49.910 64.560 ;
        RECT 50.090 64.690 51.830 64.860 ;
        RECT 50.090 64.240 50.260 64.690 ;
        RECT 49.230 64.070 50.260 64.240 ;
        RECT 50.440 63.890 50.610 64.510 ;
        RECT 51.140 64.250 51.470 64.510 ;
        RECT 48.800 63.720 50.610 63.890 ;
        RECT 50.790 63.720 51.010 64.050 ;
        RECT 50.440 63.540 50.610 63.720 ;
        RECT 48.310 62.970 48.840 63.200 ;
        RECT 48.310 62.050 48.580 62.970 ;
      LAYER li1 ;
        RECT 49.260 62.670 49.800 63.540 ;
      LAYER li1 ;
        RECT 50.440 63.370 50.660 63.540 ;
        RECT 47.120 61.420 48.070 62.050 ;
        RECT 48.250 61.550 48.580 62.050 ;
        RECT 48.760 61.420 49.350 62.300 ;
      LAYER li1 ;
        RECT 49.630 61.680 49.800 62.670 ;
        RECT 49.980 61.860 50.310 63.160 ;
      LAYER li1 ;
        RECT 50.490 62.380 50.660 63.370 ;
        RECT 50.840 63.200 51.010 63.720 ;
        RECT 51.190 63.550 51.360 64.250 ;
        RECT 51.660 64.100 51.830 64.690 ;
        RECT 52.010 64.730 52.960 64.760 ;
        RECT 52.010 64.560 52.040 64.730 ;
        RECT 52.210 64.560 52.400 64.730 ;
        RECT 52.570 64.560 52.760 64.730 ;
        RECT 52.930 64.560 52.960 64.730 ;
        RECT 52.010 64.280 52.960 64.560 ;
        RECT 53.140 64.690 54.170 64.860 ;
        RECT 53.140 64.100 53.310 64.690 ;
        RECT 51.660 64.050 53.310 64.100 ;
        RECT 51.540 63.930 53.310 64.050 ;
        RECT 51.540 63.730 51.870 63.930 ;
        RECT 53.490 63.750 53.820 64.510 ;
        RECT 54.000 64.330 54.170 64.690 ;
        RECT 54.350 64.730 55.300 64.810 ;
        RECT 54.350 64.560 54.380 64.730 ;
        RECT 54.550 64.560 54.740 64.730 ;
        RECT 54.910 64.560 55.100 64.730 ;
        RECT 55.270 64.560 55.300 64.730 ;
        RECT 54.350 64.510 55.300 64.560 ;
        RECT 54.000 64.160 55.810 64.330 ;
        RECT 52.050 63.580 53.820 63.750 ;
        RECT 52.050 63.550 52.220 63.580 ;
        RECT 51.190 63.380 52.220 63.550 ;
        RECT 55.130 63.400 55.460 63.980 ;
        RECT 50.840 62.970 51.870 63.200 ;
        RECT 51.540 62.480 51.870 62.970 ;
        RECT 52.050 62.700 52.220 63.380 ;
        RECT 52.400 63.230 55.460 63.400 ;
        RECT 52.400 62.880 52.730 63.230 ;
      LAYER li1 ;
        RECT 53.170 62.880 55.020 63.050 ;
      LAYER li1 ;
        RECT 52.050 62.530 54.670 62.700 ;
        RECT 50.490 61.880 50.760 62.380 ;
        RECT 52.050 62.300 52.220 62.530 ;
      LAYER li1 ;
        RECT 54.850 62.350 55.020 62.880 ;
      LAYER li1 ;
        RECT 51.210 62.130 52.220 62.300 ;
      LAYER li1 ;
        RECT 52.400 62.180 55.020 62.350 ;
      LAYER li1 ;
        RECT 51.210 61.880 51.540 62.130 ;
      LAYER li1 ;
        RECT 52.400 61.680 52.570 62.180 ;
        RECT 49.630 61.510 52.570 61.680 ;
      LAYER li1 ;
        RECT 53.720 61.420 54.670 62.000 ;
      LAYER li1 ;
        RECT 54.850 61.490 55.020 62.180 ;
      LAYER li1 ;
        RECT 55.200 62.380 55.460 63.230 ;
        RECT 55.640 62.810 55.810 64.160 ;
        RECT 55.990 63.900 56.240 64.810 ;
        RECT 57.050 64.730 58.000 64.760 ;
        RECT 58.830 64.730 59.730 64.760 ;
        RECT 57.050 64.560 57.080 64.730 ;
        RECT 57.250 64.560 57.440 64.730 ;
        RECT 57.610 64.560 57.800 64.730 ;
        RECT 57.970 64.560 58.000 64.730 ;
        RECT 59.000 64.560 59.190 64.730 ;
        RECT 59.360 64.560 59.550 64.730 ;
        RECT 59.720 64.560 59.730 64.730 ;
        RECT 55.990 63.730 56.870 63.900 ;
        RECT 57.050 63.730 58.000 64.560 ;
        RECT 58.400 63.760 58.650 64.230 ;
        RECT 58.830 63.940 59.730 64.560 ;
        RECT 60.340 64.730 61.280 64.790 ;
        RECT 60.340 64.560 60.360 64.730 ;
        RECT 60.530 64.560 60.720 64.730 ;
        RECT 60.890 64.560 61.080 64.730 ;
        RECT 61.250 64.560 61.280 64.730 ;
        RECT 56.190 62.990 56.520 63.490 ;
        RECT 56.700 63.410 56.870 63.730 ;
        RECT 58.400 63.590 59.410 63.760 ;
        RECT 56.700 63.240 59.060 63.410 ;
        RECT 55.640 62.640 56.810 62.810 ;
        RECT 55.200 61.670 55.530 62.380 ;
        RECT 55.990 61.840 56.320 62.380 ;
        RECT 56.530 62.140 56.810 62.640 ;
        RECT 56.990 61.840 57.160 63.240 ;
        RECT 59.240 63.060 59.410 63.590 ;
        RECT 57.370 62.890 59.410 63.060 ;
        RECT 57.370 62.500 57.700 62.890 ;
      LAYER li1 ;
        RECT 58.020 62.320 58.350 62.710 ;
      LAYER li1 ;
        RECT 55.990 61.670 57.160 61.840 ;
      LAYER li1 ;
        RECT 57.340 62.150 58.350 62.320 ;
        RECT 57.340 61.490 57.510 62.150 ;
      LAYER li1 ;
        RECT 59.180 62.050 59.410 62.890 ;
        RECT 59.910 63.060 60.160 64.060 ;
        RECT 60.340 63.250 61.280 64.560 ;
        RECT 59.910 62.730 61.280 63.060 ;
        RECT 59.910 62.550 60.120 62.730 ;
        RECT 59.790 62.050 60.120 62.550 ;
      LAYER li1 ;
        RECT 54.850 61.320 57.510 61.490 ;
      LAYER li1 ;
        RECT 57.690 61.420 58.640 61.970 ;
        RECT 59.180 61.550 59.510 62.050 ;
        RECT 60.300 61.420 61.250 62.550 ;
      LAYER li1 ;
        RECT 61.460 61.720 61.800 64.790 ;
      LAYER li1 ;
        RECT 62.170 64.780 63.620 64.810 ;
        RECT 62.170 64.610 62.420 64.780 ;
        RECT 62.590 64.610 62.780 64.780 ;
        RECT 62.950 64.610 63.220 64.780 ;
        RECT 63.390 64.610 63.620 64.780 ;
        RECT 62.170 63.740 63.620 64.610 ;
        RECT 63.930 64.730 64.880 64.810 ;
        RECT 63.930 64.560 63.960 64.730 ;
        RECT 64.130 64.560 64.320 64.730 ;
        RECT 64.490 64.560 64.680 64.730 ;
        RECT 64.850 64.560 64.880 64.730 ;
        RECT 62.400 62.300 62.730 63.080 ;
        RECT 62.940 62.750 63.270 63.740 ;
        RECT 63.930 63.230 64.880 64.560 ;
      LAYER li1 ;
        RECT 63.970 62.600 64.860 62.990 ;
        RECT 65.060 62.750 65.310 64.810 ;
      LAYER li1 ;
        RECT 65.500 64.730 66.090 64.810 ;
        RECT 65.500 64.560 65.530 64.730 ;
        RECT 65.700 64.560 65.890 64.730 ;
        RECT 66.060 64.560 66.090 64.730 ;
        RECT 65.500 63.230 66.090 64.560 ;
        RECT 66.490 64.780 67.940 64.810 ;
        RECT 66.490 64.610 66.740 64.780 ;
        RECT 66.910 64.610 67.100 64.780 ;
        RECT 67.270 64.610 67.540 64.780 ;
        RECT 67.710 64.610 67.940 64.780 ;
        RECT 66.490 63.740 67.940 64.610 ;
      LAYER li1 ;
        RECT 65.060 62.580 65.640 62.750 ;
        RECT 65.820 62.580 66.120 62.910 ;
        RECT 65.420 62.400 65.640 62.580 ;
      LAYER li1 ;
        RECT 62.400 61.900 63.700 62.300 ;
        RECT 62.090 61.420 63.700 61.900 ;
        RECT 63.930 61.420 65.240 62.400 ;
      LAYER li1 ;
        RECT 65.420 62.230 66.020 62.400 ;
        RECT 65.690 62.060 66.020 62.230 ;
      LAYER li1 ;
        RECT 66.720 62.300 67.050 63.080 ;
        RECT 67.260 62.750 67.590 63.740 ;
      LAYER li1 ;
        RECT 68.290 62.980 68.660 64.810 ;
      LAYER li1 ;
        RECT 68.840 64.730 69.420 64.810 ;
        RECT 73.690 64.780 75.140 64.810 ;
        RECT 68.840 64.560 68.860 64.730 ;
        RECT 69.030 64.560 69.220 64.730 ;
        RECT 69.390 64.560 69.420 64.730 ;
        RECT 68.840 63.230 69.420 64.560 ;
        RECT 71.570 64.730 72.880 64.760 ;
        RECT 71.570 64.560 71.600 64.730 ;
        RECT 71.770 64.560 71.960 64.730 ;
        RECT 72.130 64.560 72.320 64.730 ;
        RECT 72.490 64.560 72.680 64.730 ;
        RECT 72.850 64.560 72.880 64.730 ;
      LAYER li1 ;
        RECT 69.600 64.150 71.390 64.320 ;
        RECT 65.690 61.890 66.080 62.060 ;
      LAYER li1 ;
        RECT 66.720 61.900 68.020 62.300 ;
      LAYER li1 ;
        RECT 65.690 61.570 66.020 61.890 ;
      LAYER li1 ;
        RECT 66.410 61.420 68.020 61.900 ;
      LAYER li1 ;
        RECT 68.290 61.550 68.580 62.980 ;
      LAYER li1 ;
        RECT 68.780 62.580 69.110 62.800 ;
      LAYER li1 ;
        RECT 69.600 62.760 69.930 64.150 ;
      LAYER li1 ;
        RECT 70.710 63.640 71.040 63.970 ;
        RECT 70.110 63.470 71.040 63.640 ;
        RECT 70.110 62.580 70.280 63.470 ;
      LAYER li1 ;
        RECT 71.220 63.360 71.390 64.150 ;
      LAYER li1 ;
        RECT 71.570 63.550 72.880 64.560 ;
        RECT 73.690 64.610 73.940 64.780 ;
        RECT 74.110 64.610 74.300 64.780 ;
        RECT 74.470 64.610 74.740 64.780 ;
        RECT 74.910 64.610 75.140 64.780 ;
      LAYER li1 ;
        RECT 70.460 63.010 70.790 63.290 ;
        RECT 71.220 63.190 72.840 63.360 ;
        RECT 70.460 62.840 71.070 63.010 ;
      LAYER li1 ;
        RECT 68.780 62.410 70.720 62.580 ;
        RECT 68.760 61.420 70.370 62.230 ;
        RECT 70.550 61.970 70.720 62.410 ;
      LAYER li1 ;
        RECT 70.900 62.440 71.070 62.840 ;
        RECT 71.250 62.620 71.850 63.010 ;
        RECT 70.900 62.150 71.850 62.440 ;
      LAYER li1 ;
        RECT 72.030 62.330 72.280 62.830 ;
      LAYER li1 ;
        RECT 72.530 62.600 72.840 63.190 ;
      LAYER li1 ;
        RECT 73.060 62.330 73.310 63.970 ;
        RECT 73.690 63.740 75.140 64.610 ;
        RECT 75.450 64.730 76.400 64.810 ;
        RECT 75.450 64.560 75.480 64.730 ;
        RECT 75.650 64.560 75.840 64.730 ;
        RECT 76.010 64.560 76.200 64.730 ;
        RECT 76.370 64.560 76.400 64.730 ;
        RECT 72.030 62.160 73.310 62.330 ;
        RECT 70.550 61.550 71.040 61.970 ;
        RECT 71.220 61.420 72.880 61.970 ;
        RECT 73.060 61.550 73.310 62.160 ;
        RECT 73.920 62.300 74.250 63.080 ;
        RECT 74.460 62.750 74.790 63.740 ;
        RECT 75.450 63.230 76.400 64.560 ;
      LAYER li1 ;
        RECT 76.580 63.130 76.830 64.810 ;
      LAYER li1 ;
        RECT 77.010 64.730 77.960 64.810 ;
        RECT 77.010 64.560 77.040 64.730 ;
        RECT 77.210 64.560 77.400 64.730 ;
        RECT 77.570 64.560 77.760 64.730 ;
        RECT 77.930 64.560 77.960 64.730 ;
        RECT 77.010 63.310 77.960 64.560 ;
      LAYER li1 ;
        RECT 78.140 63.130 78.470 64.810 ;
      LAYER li1 ;
        RECT 78.650 64.730 79.600 64.810 ;
        RECT 78.650 64.560 78.680 64.730 ;
        RECT 78.850 64.560 79.040 64.730 ;
        RECT 79.210 64.560 79.400 64.730 ;
        RECT 79.570 64.560 79.600 64.730 ;
        RECT 78.650 63.350 79.600 64.560 ;
      LAYER li1 ;
        RECT 76.580 62.960 78.470 63.130 ;
        RECT 76.580 62.830 76.750 62.960 ;
        RECT 79.250 62.830 79.580 63.170 ;
        RECT 75.490 62.600 76.750 62.830 ;
      LAYER li1 ;
        RECT 76.930 62.650 78.960 62.780 ;
        RECT 79.780 62.650 80.030 64.810 ;
        RECT 80.410 64.780 81.860 64.810 ;
        RECT 80.410 64.610 80.660 64.780 ;
        RECT 80.830 64.610 81.020 64.780 ;
        RECT 81.190 64.610 81.460 64.780 ;
        RECT 81.630 64.610 81.860 64.780 ;
        RECT 80.410 63.740 81.860 64.610 ;
        RECT 82.170 64.730 82.760 64.810 ;
        RECT 82.170 64.560 82.200 64.730 ;
        RECT 82.370 64.560 82.560 64.730 ;
        RECT 82.730 64.560 82.760 64.730 ;
        RECT 76.930 62.610 80.030 62.650 ;
      LAYER li1 ;
        RECT 76.580 62.430 76.750 62.600 ;
      LAYER li1 ;
        RECT 78.790 62.480 80.030 62.610 ;
        RECT 73.920 61.900 75.220 62.300 ;
        RECT 73.610 61.420 75.220 61.900 ;
        RECT 75.450 61.420 76.400 62.380 ;
      LAYER li1 ;
        RECT 76.580 62.260 78.390 62.430 ;
        RECT 76.580 61.550 76.830 62.260 ;
      LAYER li1 ;
        RECT 77.010 61.420 77.960 62.080 ;
      LAYER li1 ;
        RECT 78.140 61.550 78.390 62.260 ;
      LAYER li1 ;
        RECT 78.570 61.420 79.520 62.300 ;
        RECT 79.700 61.550 80.030 62.480 ;
        RECT 80.640 62.300 80.970 63.080 ;
        RECT 81.180 62.750 81.510 63.740 ;
        RECT 82.170 63.230 82.760 64.560 ;
      LAYER li1 ;
        RECT 83.040 63.230 83.430 64.810 ;
      LAYER li1 ;
        RECT 83.770 64.780 85.220 64.810 ;
        RECT 83.770 64.610 84.020 64.780 ;
        RECT 84.190 64.610 84.380 64.780 ;
        RECT 84.550 64.610 84.820 64.780 ;
        RECT 84.990 64.610 85.220 64.780 ;
        RECT 83.770 63.740 85.220 64.610 ;
        RECT 85.530 64.730 86.790 64.810 ;
        RECT 85.530 64.560 85.540 64.730 ;
        RECT 85.710 64.560 85.900 64.730 ;
        RECT 86.070 64.560 86.260 64.730 ;
        RECT 86.430 64.560 86.620 64.730 ;
      LAYER li1 ;
        RECT 82.210 62.600 82.920 62.990 ;
      LAYER li1 ;
        RECT 80.640 61.900 81.940 62.300 ;
        RECT 80.330 61.420 81.940 61.900 ;
        RECT 82.170 61.420 82.760 62.380 ;
      LAYER li1 ;
        RECT 83.100 61.550 83.430 63.230 ;
      LAYER li1 ;
        RECT 84.000 62.300 84.330 63.080 ;
        RECT 84.540 62.750 84.870 63.740 ;
        RECT 85.530 63.330 86.790 64.560 ;
      LAYER li1 ;
        RECT 87.320 64.310 87.490 64.810 ;
        RECT 86.970 63.230 87.490 64.310 ;
      LAYER li1 ;
        RECT 87.750 64.730 89.060 64.810 ;
        RECT 87.750 64.560 87.780 64.730 ;
        RECT 87.950 64.560 88.140 64.730 ;
        RECT 88.310 64.560 88.500 64.730 ;
        RECT 88.670 64.560 88.860 64.730 ;
        RECT 89.030 64.560 89.060 64.730 ;
        RECT 87.750 63.350 89.060 64.560 ;
        RECT 89.530 64.780 90.980 64.810 ;
        RECT 89.530 64.610 89.780 64.780 ;
        RECT 89.950 64.610 90.140 64.780 ;
        RECT 90.310 64.610 90.580 64.780 ;
        RECT 90.750 64.610 90.980 64.780 ;
        RECT 89.530 63.740 90.980 64.610 ;
        RECT 91.770 64.730 92.720 64.810 ;
        RECT 91.770 64.560 91.800 64.730 ;
        RECT 91.970 64.560 92.160 64.730 ;
        RECT 92.330 64.560 92.520 64.730 ;
        RECT 92.690 64.560 92.720 64.730 ;
      LAYER li1 ;
        RECT 86.970 63.150 87.240 63.230 ;
        RECT 86.180 62.980 87.240 63.150 ;
        RECT 85.570 62.590 85.990 62.920 ;
        RECT 86.180 62.410 86.350 62.980 ;
        RECT 87.690 62.860 88.200 63.170 ;
        RECT 88.450 62.860 89.160 63.170 ;
        RECT 86.530 62.590 87.040 62.800 ;
      LAYER li1 ;
        RECT 87.240 62.510 89.110 62.680 ;
        RECT 84.000 61.900 85.300 62.300 ;
        RECT 83.690 61.420 85.300 61.900 ;
        RECT 85.600 61.490 85.930 62.410 ;
      LAYER li1 ;
        RECT 86.180 61.670 86.710 62.410 ;
      LAYER li1 ;
        RECT 87.240 61.490 87.410 62.510 ;
        RECT 85.600 61.320 87.410 61.490 ;
        RECT 87.590 61.420 88.690 62.330 ;
        RECT 88.860 61.580 89.110 62.510 ;
        RECT 89.760 62.300 90.090 63.080 ;
        RECT 90.300 62.750 90.630 63.740 ;
        RECT 91.770 63.230 92.720 64.560 ;
      LAYER li1 ;
        RECT 92.900 63.130 93.150 64.810 ;
      LAYER li1 ;
        RECT 93.330 64.730 94.280 64.810 ;
        RECT 93.330 64.560 93.360 64.730 ;
        RECT 93.530 64.560 93.720 64.730 ;
        RECT 93.890 64.560 94.080 64.730 ;
        RECT 94.250 64.560 94.280 64.730 ;
        RECT 93.330 63.310 94.280 64.560 ;
      LAYER li1 ;
        RECT 94.460 63.130 94.790 64.810 ;
      LAYER li1 ;
        RECT 94.970 64.730 95.920 64.810 ;
        RECT 94.970 64.560 95.000 64.730 ;
        RECT 95.170 64.560 95.360 64.730 ;
        RECT 95.530 64.560 95.720 64.730 ;
        RECT 95.890 64.560 95.920 64.730 ;
        RECT 94.970 63.350 95.920 64.560 ;
      LAYER li1 ;
        RECT 92.900 62.960 94.790 63.130 ;
        RECT 92.900 62.830 93.070 62.960 ;
        RECT 95.570 62.830 95.900 63.170 ;
        RECT 91.810 62.600 93.070 62.830 ;
      LAYER li1 ;
        RECT 93.250 62.650 95.280 62.780 ;
        RECT 96.100 62.650 96.350 64.810 ;
        RECT 96.730 64.780 98.180 64.810 ;
        RECT 96.730 64.610 96.980 64.780 ;
        RECT 97.150 64.610 97.340 64.780 ;
        RECT 97.510 64.610 97.780 64.780 ;
        RECT 97.950 64.610 98.180 64.780 ;
        RECT 96.730 63.740 98.180 64.610 ;
        RECT 93.250 62.610 96.350 62.650 ;
      LAYER li1 ;
        RECT 92.900 62.430 93.070 62.600 ;
      LAYER li1 ;
        RECT 95.110 62.480 96.350 62.610 ;
        RECT 89.760 61.900 91.060 62.300 ;
        RECT 89.450 61.420 91.060 61.900 ;
        RECT 91.770 61.420 92.720 62.380 ;
      LAYER li1 ;
        RECT 92.900 62.260 94.710 62.430 ;
        RECT 92.900 61.550 93.150 62.260 ;
      LAYER li1 ;
        RECT 93.330 61.420 94.280 62.080 ;
      LAYER li1 ;
        RECT 94.460 61.550 94.710 62.260 ;
      LAYER li1 ;
        RECT 94.890 61.420 95.840 62.300 ;
        RECT 96.020 61.550 96.350 62.480 ;
        RECT 96.960 62.300 97.290 63.080 ;
        RECT 97.500 62.750 97.830 63.740 ;
        RECT 98.660 63.150 98.910 64.810 ;
        RECT 99.090 64.730 100.340 64.810 ;
        RECT 99.260 64.560 99.450 64.730 ;
        RECT 99.620 64.560 99.810 64.730 ;
        RECT 99.980 64.560 100.170 64.730 ;
        RECT 99.090 63.330 100.340 64.560 ;
        RECT 100.520 63.150 100.690 64.810 ;
        RECT 98.660 62.980 100.690 63.150 ;
      LAYER li1 ;
        RECT 100.870 62.860 101.200 64.310 ;
        RECT 98.530 62.560 99.720 62.800 ;
        RECT 99.970 62.560 100.320 62.800 ;
        RECT 101.380 62.680 101.640 64.810 ;
      LAYER li1 ;
        RECT 102.260 64.780 105.000 64.800 ;
        RECT 102.260 64.610 102.470 64.780 ;
        RECT 102.640 64.610 102.910 64.780 ;
        RECT 103.080 64.610 103.320 64.780 ;
        RECT 103.490 64.610 103.750 64.780 ;
        RECT 103.920 64.610 104.190 64.780 ;
        RECT 104.360 64.610 104.600 64.780 ;
        RECT 104.770 64.610 105.000 64.780 ;
        RECT 102.260 63.730 105.000 64.610 ;
        RECT 106.710 64.730 107.300 64.760 ;
        RECT 106.710 64.560 106.740 64.730 ;
        RECT 106.910 64.560 107.100 64.730 ;
        RECT 107.270 64.560 107.300 64.730 ;
      LAYER li1 ;
        RECT 100.620 62.510 101.640 62.680 ;
      LAYER li1 ;
        RECT 96.960 61.900 98.260 62.300 ;
        RECT 96.650 61.420 98.260 61.900 ;
        RECT 98.730 61.420 100.440 62.380 ;
      LAYER li1 ;
        RECT 100.620 61.550 100.870 62.510 ;
      LAYER li1 ;
        RECT 102.500 62.410 102.830 63.080 ;
        RECT 103.230 62.750 103.560 63.730 ;
        RECT 103.780 62.410 104.110 63.080 ;
        RECT 104.510 62.750 104.840 63.730 ;
        RECT 106.190 63.580 106.520 64.510 ;
        RECT 106.710 63.780 107.300 64.560 ;
        RECT 107.480 64.690 108.920 64.860 ;
        RECT 107.480 63.580 107.650 64.690 ;
        RECT 106.190 63.410 107.650 63.580 ;
        RECT 101.080 61.420 101.670 62.330 ;
        RECT 102.340 61.410 105.070 62.410 ;
        RECT 106.190 61.550 106.460 63.410 ;
        RECT 107.320 62.910 107.650 63.410 ;
        RECT 107.830 63.200 108.080 64.510 ;
        RECT 108.320 63.890 108.570 64.510 ;
        RECT 108.750 64.240 108.920 64.690 ;
        RECT 109.100 64.730 109.430 64.760 ;
        RECT 109.100 64.560 109.130 64.730 ;
        RECT 109.300 64.560 109.430 64.730 ;
        RECT 109.100 64.420 109.430 64.560 ;
        RECT 109.610 64.690 111.350 64.860 ;
        RECT 109.610 64.240 109.780 64.690 ;
        RECT 108.750 64.070 109.780 64.240 ;
        RECT 109.960 63.890 110.130 64.510 ;
        RECT 110.660 64.250 110.990 64.510 ;
        RECT 108.320 63.720 110.130 63.890 ;
        RECT 110.310 63.720 110.530 64.050 ;
        RECT 109.960 63.540 110.130 63.720 ;
        RECT 107.830 62.970 108.360 63.200 ;
        RECT 107.830 62.050 108.100 62.970 ;
      LAYER li1 ;
        RECT 108.780 62.670 109.320 63.540 ;
      LAYER li1 ;
        RECT 109.960 63.370 110.180 63.540 ;
        RECT 106.640 61.420 107.590 62.050 ;
        RECT 107.770 61.550 108.100 62.050 ;
        RECT 108.280 61.420 108.870 62.300 ;
      LAYER li1 ;
        RECT 109.150 61.680 109.320 62.670 ;
        RECT 109.500 61.860 109.830 63.160 ;
      LAYER li1 ;
        RECT 110.010 62.380 110.180 63.370 ;
        RECT 110.360 63.200 110.530 63.720 ;
        RECT 110.710 63.550 110.880 64.250 ;
        RECT 111.180 64.100 111.350 64.690 ;
        RECT 111.530 64.730 112.480 64.760 ;
        RECT 111.530 64.560 111.560 64.730 ;
        RECT 111.730 64.560 111.920 64.730 ;
        RECT 112.090 64.560 112.280 64.730 ;
        RECT 112.450 64.560 112.480 64.730 ;
        RECT 111.530 64.280 112.480 64.560 ;
        RECT 112.660 64.690 113.690 64.860 ;
        RECT 112.660 64.100 112.830 64.690 ;
        RECT 111.180 64.050 112.830 64.100 ;
        RECT 111.060 63.930 112.830 64.050 ;
        RECT 111.060 63.730 111.390 63.930 ;
        RECT 113.010 63.750 113.340 64.510 ;
        RECT 113.520 64.330 113.690 64.690 ;
        RECT 113.870 64.730 114.820 64.810 ;
        RECT 113.870 64.560 113.900 64.730 ;
        RECT 114.070 64.560 114.260 64.730 ;
        RECT 114.430 64.560 114.620 64.730 ;
        RECT 114.790 64.560 114.820 64.730 ;
        RECT 113.870 64.510 114.820 64.560 ;
        RECT 113.520 64.160 115.330 64.330 ;
        RECT 111.570 63.580 113.340 63.750 ;
        RECT 111.570 63.550 111.740 63.580 ;
        RECT 110.710 63.380 111.740 63.550 ;
        RECT 114.650 63.400 114.980 63.980 ;
        RECT 110.360 62.970 111.390 63.200 ;
        RECT 111.060 62.480 111.390 62.970 ;
        RECT 111.570 62.700 111.740 63.380 ;
        RECT 111.920 63.230 114.980 63.400 ;
        RECT 111.920 62.880 112.250 63.230 ;
      LAYER li1 ;
        RECT 112.690 62.880 114.540 63.050 ;
      LAYER li1 ;
        RECT 111.570 62.530 114.190 62.700 ;
        RECT 110.010 61.880 110.280 62.380 ;
        RECT 111.570 62.300 111.740 62.530 ;
      LAYER li1 ;
        RECT 114.370 62.350 114.540 62.880 ;
      LAYER li1 ;
        RECT 110.730 62.130 111.740 62.300 ;
      LAYER li1 ;
        RECT 111.920 62.180 114.540 62.350 ;
      LAYER li1 ;
        RECT 110.730 61.880 111.060 62.130 ;
      LAYER li1 ;
        RECT 111.920 61.680 112.090 62.180 ;
        RECT 109.150 61.510 112.090 61.680 ;
      LAYER li1 ;
        RECT 113.240 61.420 114.190 62.000 ;
      LAYER li1 ;
        RECT 114.370 61.490 114.540 62.180 ;
      LAYER li1 ;
        RECT 114.720 62.380 114.980 63.230 ;
        RECT 115.160 62.810 115.330 64.160 ;
        RECT 115.510 63.900 115.760 64.810 ;
        RECT 116.570 64.730 117.520 64.760 ;
        RECT 118.350 64.730 119.250 64.760 ;
        RECT 116.570 64.560 116.600 64.730 ;
        RECT 116.770 64.560 116.960 64.730 ;
        RECT 117.130 64.560 117.320 64.730 ;
        RECT 117.490 64.560 117.520 64.730 ;
        RECT 118.520 64.560 118.710 64.730 ;
        RECT 118.880 64.560 119.070 64.730 ;
        RECT 119.240 64.560 119.250 64.730 ;
        RECT 115.510 63.730 116.390 63.900 ;
        RECT 116.570 63.730 117.520 64.560 ;
        RECT 117.920 63.760 118.170 64.230 ;
        RECT 118.350 63.940 119.250 64.560 ;
        RECT 119.860 64.730 120.800 64.790 ;
        RECT 119.860 64.560 119.880 64.730 ;
        RECT 120.050 64.560 120.240 64.730 ;
        RECT 120.410 64.560 120.600 64.730 ;
        RECT 120.770 64.560 120.800 64.730 ;
        RECT 115.710 62.990 116.040 63.490 ;
        RECT 116.220 63.410 116.390 63.730 ;
        RECT 117.920 63.590 118.930 63.760 ;
        RECT 116.220 63.240 118.580 63.410 ;
        RECT 115.160 62.640 116.330 62.810 ;
        RECT 114.720 61.670 115.050 62.380 ;
        RECT 115.510 61.840 115.840 62.380 ;
        RECT 116.050 62.140 116.330 62.640 ;
        RECT 116.510 61.840 116.680 63.240 ;
        RECT 118.760 63.060 118.930 63.590 ;
        RECT 116.890 62.890 118.930 63.060 ;
        RECT 116.890 62.500 117.220 62.890 ;
      LAYER li1 ;
        RECT 117.540 62.430 117.870 62.710 ;
        RECT 117.540 62.320 117.920 62.430 ;
      LAYER li1 ;
        RECT 115.510 61.670 116.680 61.840 ;
      LAYER li1 ;
        RECT 116.860 62.260 117.920 62.320 ;
        RECT 116.860 62.150 117.870 62.260 ;
        RECT 116.860 61.490 117.030 62.150 ;
      LAYER li1 ;
        RECT 118.700 62.050 118.930 62.890 ;
        RECT 119.430 63.060 119.680 64.060 ;
        RECT 119.860 63.250 120.800 64.560 ;
        RECT 119.430 62.730 120.800 63.060 ;
        RECT 119.430 62.550 119.640 62.730 ;
        RECT 119.310 62.050 119.640 62.550 ;
      LAYER li1 ;
        RECT 114.370 61.320 117.030 61.490 ;
      LAYER li1 ;
        RECT 117.210 61.420 118.160 61.970 ;
        RECT 118.700 61.550 119.030 62.050 ;
        RECT 119.820 61.420 120.770 62.550 ;
      LAYER li1 ;
        RECT 120.980 61.720 121.320 64.790 ;
      LAYER li1 ;
        RECT 121.690 64.780 123.140 64.810 ;
        RECT 121.690 64.610 121.940 64.780 ;
        RECT 122.110 64.610 122.300 64.780 ;
        RECT 122.470 64.610 122.740 64.780 ;
        RECT 122.910 64.610 123.140 64.780 ;
        RECT 121.690 63.740 123.140 64.610 ;
        RECT 123.990 64.730 124.580 64.760 ;
        RECT 123.990 64.560 124.020 64.730 ;
        RECT 124.190 64.560 124.380 64.730 ;
        RECT 124.550 64.560 124.580 64.730 ;
        RECT 121.920 62.300 122.250 63.080 ;
        RECT 122.460 62.750 122.790 63.740 ;
        RECT 123.470 63.580 123.800 64.510 ;
        RECT 123.990 63.780 124.580 64.560 ;
        RECT 124.760 64.690 126.200 64.860 ;
        RECT 124.760 63.580 124.930 64.690 ;
        RECT 123.470 63.410 124.930 63.580 ;
        RECT 121.920 61.900 123.220 62.300 ;
        RECT 121.610 61.420 123.220 61.900 ;
        RECT 123.470 61.550 123.740 63.410 ;
        RECT 124.600 62.910 124.930 63.410 ;
        RECT 125.110 63.200 125.360 64.510 ;
        RECT 125.600 63.890 125.850 64.510 ;
        RECT 126.030 64.240 126.200 64.690 ;
        RECT 126.380 64.730 126.710 64.760 ;
        RECT 126.380 64.560 126.410 64.730 ;
        RECT 126.580 64.560 126.710 64.730 ;
        RECT 126.380 64.420 126.710 64.560 ;
        RECT 126.890 64.690 128.630 64.860 ;
        RECT 126.890 64.240 127.060 64.690 ;
        RECT 126.030 64.070 127.060 64.240 ;
        RECT 127.240 63.890 127.410 64.510 ;
        RECT 127.940 64.250 128.270 64.510 ;
        RECT 125.600 63.720 127.410 63.890 ;
        RECT 127.590 63.720 127.810 64.050 ;
        RECT 127.240 63.540 127.410 63.720 ;
        RECT 125.110 62.970 125.640 63.200 ;
        RECT 125.110 62.050 125.380 62.970 ;
      LAYER li1 ;
        RECT 126.060 62.670 126.600 63.540 ;
      LAYER li1 ;
        RECT 127.240 63.370 127.460 63.540 ;
        RECT 123.920 61.420 124.870 62.050 ;
        RECT 125.050 61.550 125.380 62.050 ;
        RECT 125.560 61.420 126.150 62.300 ;
      LAYER li1 ;
        RECT 126.430 61.680 126.600 62.670 ;
        RECT 126.780 61.860 127.110 63.160 ;
      LAYER li1 ;
        RECT 127.290 62.380 127.460 63.370 ;
        RECT 127.640 63.200 127.810 63.720 ;
        RECT 127.990 63.550 128.160 64.250 ;
        RECT 128.460 64.100 128.630 64.690 ;
        RECT 128.810 64.730 129.760 64.760 ;
        RECT 128.810 64.560 128.840 64.730 ;
        RECT 129.010 64.560 129.200 64.730 ;
        RECT 129.370 64.560 129.560 64.730 ;
        RECT 129.730 64.560 129.760 64.730 ;
        RECT 128.810 64.280 129.760 64.560 ;
        RECT 129.940 64.690 130.970 64.860 ;
        RECT 129.940 64.100 130.110 64.690 ;
        RECT 128.460 64.050 130.110 64.100 ;
        RECT 128.340 63.930 130.110 64.050 ;
        RECT 128.340 63.730 128.670 63.930 ;
        RECT 130.290 63.750 130.620 64.510 ;
        RECT 130.800 64.330 130.970 64.690 ;
        RECT 131.150 64.730 132.100 64.810 ;
        RECT 131.150 64.560 131.180 64.730 ;
        RECT 131.350 64.560 131.540 64.730 ;
        RECT 131.710 64.560 131.900 64.730 ;
        RECT 132.070 64.560 132.100 64.730 ;
        RECT 131.150 64.510 132.100 64.560 ;
        RECT 130.800 64.160 132.610 64.330 ;
        RECT 128.850 63.580 130.620 63.750 ;
        RECT 128.850 63.550 129.020 63.580 ;
        RECT 127.990 63.380 129.020 63.550 ;
        RECT 131.930 63.400 132.260 63.980 ;
        RECT 127.640 62.970 128.670 63.200 ;
        RECT 128.340 62.480 128.670 62.970 ;
        RECT 128.850 62.700 129.020 63.380 ;
        RECT 129.200 63.230 132.260 63.400 ;
        RECT 129.200 62.880 129.530 63.230 ;
      LAYER li1 ;
        RECT 129.970 62.880 131.820 63.050 ;
      LAYER li1 ;
        RECT 128.850 62.530 131.470 62.700 ;
        RECT 127.290 61.880 127.560 62.380 ;
        RECT 128.850 62.300 129.020 62.530 ;
      LAYER li1 ;
        RECT 131.650 62.350 131.820 62.880 ;
      LAYER li1 ;
        RECT 128.010 62.130 129.020 62.300 ;
      LAYER li1 ;
        RECT 129.200 62.180 131.820 62.350 ;
      LAYER li1 ;
        RECT 128.010 61.880 128.340 62.130 ;
      LAYER li1 ;
        RECT 129.200 61.680 129.370 62.180 ;
        RECT 126.430 61.510 129.370 61.680 ;
      LAYER li1 ;
        RECT 130.520 61.420 131.470 62.000 ;
      LAYER li1 ;
        RECT 131.650 61.490 131.820 62.180 ;
      LAYER li1 ;
        RECT 132.000 62.380 132.260 63.230 ;
        RECT 132.440 62.810 132.610 64.160 ;
        RECT 132.790 63.900 133.040 64.810 ;
        RECT 133.850 64.730 134.800 64.760 ;
        RECT 135.630 64.730 136.530 64.760 ;
        RECT 133.850 64.560 133.880 64.730 ;
        RECT 134.050 64.560 134.240 64.730 ;
        RECT 134.410 64.560 134.600 64.730 ;
        RECT 134.770 64.560 134.800 64.730 ;
        RECT 135.800 64.560 135.990 64.730 ;
        RECT 136.160 64.560 136.350 64.730 ;
        RECT 136.520 64.560 136.530 64.730 ;
        RECT 132.790 63.730 133.670 63.900 ;
        RECT 133.850 63.730 134.800 64.560 ;
        RECT 135.200 63.760 135.450 64.230 ;
        RECT 135.630 63.940 136.530 64.560 ;
        RECT 137.140 64.730 138.080 64.790 ;
        RECT 137.140 64.560 137.160 64.730 ;
        RECT 137.330 64.560 137.520 64.730 ;
        RECT 137.690 64.560 137.880 64.730 ;
        RECT 138.050 64.560 138.080 64.730 ;
        RECT 132.990 62.990 133.320 63.490 ;
        RECT 133.500 63.410 133.670 63.730 ;
        RECT 135.200 63.590 136.210 63.760 ;
        RECT 133.500 63.240 135.860 63.410 ;
        RECT 132.440 62.640 133.610 62.810 ;
        RECT 132.000 61.670 132.330 62.380 ;
        RECT 132.790 61.840 133.120 62.380 ;
        RECT 133.330 62.140 133.610 62.640 ;
        RECT 133.790 61.840 133.960 63.240 ;
        RECT 136.040 63.060 136.210 63.590 ;
        RECT 134.170 62.890 136.210 63.060 ;
        RECT 134.170 62.500 134.500 62.890 ;
      LAYER li1 ;
        RECT 134.820 62.430 135.150 62.710 ;
        RECT 134.820 62.320 135.200 62.430 ;
      LAYER li1 ;
        RECT 132.790 61.670 133.960 61.840 ;
      LAYER li1 ;
        RECT 134.140 62.260 135.200 62.320 ;
        RECT 134.140 62.150 135.150 62.260 ;
        RECT 134.140 61.490 134.310 62.150 ;
      LAYER li1 ;
        RECT 135.980 62.050 136.210 62.890 ;
        RECT 136.710 63.060 136.960 64.060 ;
        RECT 137.140 63.250 138.080 64.560 ;
        RECT 136.710 62.730 138.080 63.060 ;
        RECT 136.710 62.550 136.920 62.730 ;
        RECT 136.590 62.050 136.920 62.550 ;
      LAYER li1 ;
        RECT 131.650 61.320 134.310 61.490 ;
      LAYER li1 ;
        RECT 134.490 61.420 135.440 61.970 ;
        RECT 135.980 61.550 136.310 62.050 ;
        RECT 137.100 61.420 138.050 62.550 ;
      LAYER li1 ;
        RECT 138.260 61.720 138.600 64.790 ;
      LAYER li1 ;
        RECT 138.970 64.780 140.420 64.810 ;
        RECT 138.970 64.610 139.220 64.780 ;
        RECT 139.390 64.610 139.580 64.780 ;
        RECT 139.750 64.610 140.020 64.780 ;
        RECT 140.190 64.610 140.420 64.780 ;
        RECT 138.970 63.740 140.420 64.610 ;
        RECT 139.200 62.300 139.530 63.080 ;
        RECT 139.740 62.750 140.070 63.740 ;
        RECT 139.200 61.900 140.500 62.300 ;
        RECT 138.890 61.420 140.500 61.900 ;
        RECT 5.760 60.960 5.920 61.140 ;
        RECT 6.090 60.960 6.400 61.140 ;
        RECT 6.570 60.960 6.880 61.140 ;
        RECT 7.050 60.960 7.360 61.140 ;
        RECT 7.530 60.960 7.840 61.140 ;
        RECT 8.010 60.960 8.320 61.140 ;
        RECT 8.490 60.960 8.800 61.140 ;
        RECT 8.970 60.960 9.280 61.140 ;
        RECT 9.450 60.960 9.760 61.140 ;
        RECT 9.930 60.960 10.240 61.140 ;
        RECT 10.410 60.960 10.720 61.140 ;
        RECT 10.890 60.960 11.200 61.140 ;
        RECT 11.370 60.960 11.680 61.140 ;
        RECT 11.850 60.960 12.160 61.140 ;
        RECT 12.330 60.960 12.640 61.140 ;
        RECT 12.810 60.960 13.120 61.140 ;
        RECT 13.290 60.960 13.600 61.140 ;
        RECT 13.770 60.960 14.080 61.140 ;
        RECT 14.250 60.960 14.560 61.140 ;
        RECT 14.730 60.960 15.040 61.140 ;
        RECT 15.210 60.960 15.520 61.140 ;
        RECT 15.690 60.960 16.000 61.140 ;
        RECT 16.170 60.960 16.480 61.140 ;
        RECT 16.650 60.960 16.960 61.140 ;
        RECT 17.130 60.960 17.440 61.140 ;
        RECT 17.610 60.960 17.920 61.140 ;
        RECT 18.090 60.960 18.400 61.140 ;
        RECT 18.570 60.960 18.880 61.140 ;
        RECT 19.050 60.960 19.360 61.140 ;
        RECT 19.530 60.960 19.840 61.140 ;
        RECT 20.010 60.960 20.320 61.140 ;
        RECT 20.490 60.960 20.800 61.140 ;
        RECT 20.970 60.960 21.280 61.140 ;
        RECT 21.450 60.960 21.760 61.140 ;
        RECT 21.930 60.960 22.240 61.140 ;
        RECT 22.410 60.960 22.720 61.140 ;
        RECT 22.890 60.960 23.200 61.140 ;
        RECT 23.370 60.960 23.680 61.140 ;
        RECT 23.850 60.960 24.160 61.140 ;
        RECT 24.330 60.960 24.640 61.140 ;
        RECT 24.810 60.960 25.120 61.140 ;
        RECT 25.290 60.960 25.600 61.140 ;
        RECT 25.770 60.960 26.080 61.140 ;
        RECT 26.250 60.960 26.560 61.140 ;
        RECT 26.730 60.960 27.040 61.140 ;
        RECT 27.210 60.960 27.520 61.140 ;
        RECT 27.690 60.960 28.000 61.140 ;
        RECT 28.170 60.960 28.480 61.140 ;
        RECT 28.650 60.960 28.960 61.140 ;
        RECT 29.130 60.960 29.440 61.140 ;
        RECT 29.610 60.960 29.920 61.140 ;
        RECT 30.090 60.960 30.400 61.140 ;
        RECT 30.570 60.960 30.880 61.140 ;
        RECT 31.050 60.960 31.360 61.140 ;
        RECT 31.530 60.960 31.840 61.140 ;
        RECT 32.010 60.960 32.320 61.140 ;
        RECT 32.490 60.960 32.800 61.140 ;
        RECT 32.970 60.960 33.280 61.140 ;
        RECT 33.450 60.960 33.760 61.140 ;
        RECT 33.930 60.960 34.240 61.140 ;
        RECT 34.410 60.960 34.720 61.140 ;
        RECT 34.890 60.960 35.200 61.140 ;
        RECT 35.370 60.960 35.680 61.140 ;
        RECT 35.850 60.960 36.160 61.140 ;
        RECT 36.330 60.960 36.640 61.140 ;
        RECT 36.810 60.960 37.120 61.140 ;
        RECT 37.290 60.960 37.600 61.140 ;
        RECT 37.770 60.960 38.080 61.140 ;
        RECT 38.250 60.960 38.560 61.140 ;
        RECT 38.730 60.960 39.040 61.140 ;
        RECT 39.210 60.960 39.520 61.140 ;
        RECT 39.690 60.960 40.000 61.140 ;
        RECT 40.170 60.960 40.480 61.140 ;
        RECT 40.650 60.960 40.960 61.140 ;
        RECT 41.130 60.960 41.440 61.140 ;
        RECT 41.610 60.960 41.920 61.140 ;
        RECT 42.090 60.960 42.400 61.140 ;
        RECT 42.570 60.960 42.880 61.140 ;
        RECT 43.050 60.960 43.360 61.140 ;
        RECT 43.530 60.960 43.840 61.140 ;
        RECT 44.010 60.960 44.320 61.140 ;
        RECT 44.490 60.960 44.800 61.140 ;
        RECT 44.970 60.960 45.280 61.140 ;
        RECT 45.450 60.960 45.760 61.140 ;
        RECT 45.930 60.960 46.240 61.140 ;
        RECT 46.410 60.960 46.720 61.140 ;
        RECT 46.890 60.960 47.200 61.140 ;
        RECT 47.370 60.960 47.680 61.140 ;
        RECT 47.850 60.960 48.160 61.140 ;
        RECT 48.330 60.960 48.640 61.140 ;
        RECT 48.810 60.960 49.120 61.140 ;
        RECT 49.290 60.960 49.600 61.140 ;
        RECT 49.770 60.960 50.080 61.140 ;
        RECT 50.250 60.960 50.560 61.140 ;
        RECT 50.730 60.960 51.040 61.140 ;
        RECT 51.210 60.960 51.520 61.140 ;
        RECT 51.690 60.960 52.000 61.140 ;
        RECT 52.170 60.960 52.480 61.140 ;
        RECT 52.650 60.960 52.960 61.140 ;
        RECT 53.130 60.960 53.440 61.140 ;
        RECT 53.610 60.960 53.920 61.140 ;
        RECT 54.090 60.960 54.400 61.140 ;
        RECT 54.570 60.960 54.880 61.140 ;
        RECT 55.050 60.960 55.360 61.140 ;
        RECT 55.530 60.960 55.840 61.140 ;
        RECT 56.010 60.960 56.320 61.140 ;
        RECT 56.490 60.960 56.800 61.140 ;
        RECT 56.970 60.960 57.280 61.140 ;
        RECT 57.450 60.960 57.760 61.140 ;
        RECT 57.930 60.960 58.240 61.140 ;
        RECT 58.410 60.960 58.720 61.140 ;
        RECT 58.890 60.960 59.200 61.140 ;
        RECT 59.370 60.960 59.680 61.140 ;
        RECT 59.850 60.960 60.160 61.140 ;
        RECT 60.330 60.960 60.640 61.140 ;
        RECT 60.810 60.960 61.120 61.140 ;
        RECT 61.290 60.960 61.600 61.140 ;
        RECT 61.770 60.960 62.080 61.140 ;
        RECT 62.250 60.960 62.560 61.140 ;
        RECT 62.730 60.960 63.040 61.140 ;
        RECT 63.210 60.960 63.520 61.140 ;
        RECT 63.690 60.960 64.000 61.140 ;
        RECT 64.170 60.960 64.480 61.140 ;
        RECT 64.650 60.960 64.960 61.140 ;
        RECT 65.130 60.960 65.440 61.140 ;
        RECT 65.610 60.960 65.920 61.140 ;
        RECT 66.090 60.960 66.400 61.140 ;
        RECT 66.570 60.960 66.880 61.140 ;
        RECT 67.050 60.960 67.360 61.140 ;
        RECT 67.530 60.960 67.840 61.140 ;
        RECT 68.010 60.960 68.320 61.140 ;
        RECT 68.490 60.960 68.800 61.140 ;
        RECT 68.970 60.960 69.280 61.140 ;
        RECT 69.450 60.960 69.760 61.140 ;
        RECT 69.930 60.960 70.240 61.140 ;
        RECT 70.410 60.960 70.720 61.140 ;
        RECT 70.890 60.960 71.200 61.140 ;
        RECT 71.370 60.960 71.680 61.140 ;
        RECT 71.850 60.960 72.160 61.140 ;
        RECT 72.330 60.960 72.640 61.140 ;
        RECT 72.810 60.960 73.120 61.140 ;
        RECT 73.290 60.960 73.600 61.140 ;
        RECT 73.770 60.960 74.080 61.140 ;
        RECT 74.250 60.960 74.560 61.140 ;
        RECT 74.730 60.960 75.040 61.140 ;
        RECT 75.210 60.960 75.520 61.140 ;
        RECT 75.690 60.960 76.000 61.140 ;
        RECT 76.170 60.960 76.480 61.140 ;
        RECT 76.650 60.960 76.960 61.140 ;
        RECT 77.130 60.960 77.440 61.140 ;
        RECT 77.610 60.960 77.920 61.140 ;
        RECT 78.090 60.960 78.400 61.140 ;
        RECT 78.570 60.960 78.880 61.140 ;
        RECT 79.050 60.960 79.360 61.140 ;
        RECT 79.530 60.960 79.840 61.140 ;
        RECT 80.010 60.960 80.320 61.140 ;
        RECT 80.490 60.960 80.800 61.140 ;
        RECT 80.970 60.960 81.280 61.140 ;
        RECT 81.450 60.960 81.760 61.140 ;
        RECT 81.930 60.960 82.240 61.140 ;
        RECT 82.410 60.960 82.720 61.140 ;
        RECT 82.890 60.960 83.200 61.140 ;
        RECT 83.370 60.960 83.680 61.140 ;
        RECT 83.850 60.960 84.160 61.140 ;
        RECT 84.330 60.960 84.640 61.140 ;
        RECT 84.810 60.960 85.120 61.140 ;
        RECT 85.290 60.960 85.600 61.140 ;
        RECT 85.770 60.960 86.080 61.140 ;
        RECT 86.250 60.960 86.560 61.140 ;
        RECT 86.730 60.960 87.040 61.140 ;
        RECT 87.210 60.960 87.520 61.140 ;
        RECT 87.690 60.960 88.000 61.140 ;
        RECT 88.170 60.960 88.480 61.140 ;
        RECT 88.650 60.960 88.960 61.140 ;
        RECT 89.130 60.960 89.440 61.140 ;
        RECT 89.610 60.960 89.920 61.140 ;
        RECT 90.090 60.960 90.400 61.140 ;
        RECT 90.570 60.960 90.880 61.140 ;
        RECT 91.050 60.960 91.200 61.140 ;
        RECT 91.680 60.960 91.840 61.140 ;
        RECT 92.010 60.960 92.320 61.140 ;
        RECT 92.490 60.960 92.800 61.140 ;
        RECT 92.970 60.960 93.280 61.140 ;
        RECT 93.450 60.960 93.760 61.140 ;
        RECT 93.930 60.960 94.240 61.140 ;
        RECT 94.410 60.960 94.720 61.140 ;
        RECT 94.890 60.960 95.200 61.140 ;
        RECT 95.370 60.960 95.680 61.140 ;
        RECT 95.850 60.960 96.160 61.140 ;
        RECT 96.330 60.960 96.640 61.140 ;
        RECT 96.810 60.960 97.120 61.140 ;
        RECT 97.290 60.960 97.600 61.140 ;
        RECT 97.770 60.960 98.080 61.140 ;
        RECT 98.250 60.960 98.560 61.140 ;
        RECT 98.730 60.960 99.040 61.140 ;
        RECT 99.210 60.960 99.520 61.140 ;
        RECT 99.690 60.960 100.000 61.140 ;
        RECT 100.170 60.960 100.480 61.140 ;
        RECT 100.650 60.960 100.960 61.140 ;
        RECT 101.130 60.960 101.440 61.140 ;
        RECT 101.610 60.960 101.920 61.140 ;
        RECT 102.090 60.960 102.400 61.140 ;
        RECT 102.570 60.960 102.880 61.140 ;
        RECT 103.050 60.960 103.360 61.140 ;
        RECT 103.530 60.960 103.840 61.140 ;
        RECT 104.010 60.960 104.320 61.140 ;
        RECT 104.490 60.960 104.800 61.140 ;
        RECT 104.970 60.960 105.280 61.140 ;
        RECT 105.450 60.960 105.600 61.140 ;
        RECT 106.080 60.960 106.240 61.140 ;
        RECT 106.410 60.960 106.720 61.140 ;
        RECT 106.890 60.960 107.200 61.140 ;
        RECT 107.370 60.960 107.680 61.140 ;
        RECT 107.850 60.960 108.160 61.140 ;
        RECT 108.330 60.960 108.640 61.140 ;
        RECT 108.810 60.960 109.120 61.140 ;
        RECT 109.290 60.960 109.600 61.140 ;
        RECT 109.770 60.960 110.080 61.140 ;
        RECT 110.250 60.960 110.560 61.140 ;
        RECT 110.730 60.960 111.040 61.140 ;
        RECT 111.210 60.960 111.520 61.140 ;
        RECT 111.690 60.960 112.000 61.140 ;
        RECT 112.170 60.960 112.480 61.140 ;
        RECT 112.650 60.960 112.960 61.140 ;
        RECT 113.130 60.960 113.440 61.140 ;
        RECT 113.610 60.960 113.920 61.140 ;
        RECT 114.090 60.960 114.400 61.140 ;
        RECT 114.570 60.960 114.880 61.140 ;
        RECT 115.050 60.960 115.360 61.140 ;
        RECT 115.530 60.960 115.840 61.140 ;
        RECT 116.010 60.960 116.320 61.140 ;
        RECT 116.490 60.960 116.800 61.140 ;
        RECT 116.970 60.960 117.280 61.140 ;
        RECT 117.450 60.960 117.760 61.140 ;
        RECT 117.930 60.960 118.240 61.140 ;
        RECT 118.410 60.960 118.720 61.140 ;
        RECT 118.890 60.960 119.200 61.140 ;
        RECT 119.370 60.960 119.680 61.140 ;
        RECT 119.850 60.960 120.160 61.140 ;
        RECT 120.330 60.960 120.640 61.140 ;
        RECT 120.810 60.960 121.120 61.140 ;
        RECT 121.290 60.960 121.600 61.140 ;
        RECT 121.770 60.960 122.080 61.140 ;
        RECT 122.250 60.960 122.560 61.140 ;
        RECT 122.730 60.960 123.040 61.140 ;
        RECT 123.210 60.960 123.520 61.140 ;
        RECT 123.690 60.960 124.000 61.140 ;
        RECT 124.170 60.960 124.480 61.140 ;
        RECT 124.650 60.960 124.960 61.140 ;
        RECT 125.130 60.960 125.440 61.140 ;
        RECT 125.610 60.960 125.920 61.140 ;
        RECT 126.090 60.960 126.400 61.140 ;
        RECT 126.570 60.960 126.880 61.140 ;
        RECT 127.050 60.960 127.360 61.140 ;
        RECT 127.530 60.960 127.840 61.140 ;
        RECT 128.010 60.960 128.320 61.140 ;
        RECT 128.490 60.960 128.800 61.140 ;
        RECT 128.970 60.960 129.280 61.140 ;
        RECT 129.450 60.960 129.760 61.140 ;
        RECT 129.930 60.960 130.240 61.140 ;
        RECT 130.410 60.960 130.720 61.140 ;
        RECT 130.890 60.960 131.200 61.140 ;
        RECT 131.370 60.960 131.680 61.140 ;
        RECT 131.850 60.960 132.160 61.140 ;
        RECT 132.330 60.960 132.640 61.140 ;
        RECT 132.810 60.960 133.120 61.140 ;
        RECT 133.290 60.960 133.600 61.140 ;
        RECT 133.770 60.960 134.080 61.140 ;
        RECT 134.250 60.960 134.560 61.140 ;
        RECT 134.730 60.960 135.040 61.140 ;
        RECT 135.210 60.960 135.520 61.140 ;
        RECT 135.690 60.960 136.000 61.140 ;
        RECT 136.170 60.960 136.480 61.140 ;
        RECT 136.650 60.960 136.960 61.140 ;
        RECT 137.130 60.960 137.440 61.140 ;
        RECT 137.610 60.960 137.920 61.140 ;
        RECT 138.090 60.960 138.400 61.140 ;
        RECT 138.570 60.960 138.880 61.140 ;
        RECT 139.050 60.960 139.360 61.140 ;
        RECT 139.530 60.960 139.840 61.140 ;
        RECT 140.010 60.960 140.320 61.140 ;
        RECT 140.490 60.960 140.800 61.140 ;
        RECT 140.970 60.960 141.280 61.140 ;
        RECT 141.450 60.960 141.600 61.140 ;
        RECT 5.930 60.650 7.540 60.680 ;
        RECT 5.930 60.480 5.980 60.650 ;
        RECT 6.150 60.480 6.420 60.650 ;
        RECT 6.590 60.480 6.860 60.650 ;
        RECT 7.030 60.480 7.270 60.650 ;
        RECT 7.440 60.480 7.540 60.650 ;
        RECT 8.240 60.650 9.190 60.680 ;
        RECT 5.930 60.200 7.540 60.480 ;
        RECT 6.240 59.800 7.540 60.200 ;
        RECT 6.240 59.020 6.570 59.800 ;
        RECT 6.780 58.360 7.110 59.350 ;
        RECT 7.790 58.690 8.060 60.550 ;
        RECT 8.240 60.480 8.270 60.650 ;
        RECT 8.440 60.480 8.630 60.650 ;
        RECT 8.800 60.480 8.990 60.650 ;
        RECT 9.160 60.480 9.190 60.650 ;
        RECT 9.880 60.650 10.470 60.680 ;
        RECT 8.240 60.050 9.190 60.480 ;
        RECT 9.370 60.050 9.700 60.550 ;
        RECT 8.920 58.690 9.250 59.190 ;
        RECT 7.790 58.520 9.250 58.690 ;
        RECT 6.010 57.490 7.460 58.360 ;
        RECT 7.790 57.590 8.120 58.520 ;
        RECT 6.010 57.320 6.260 57.490 ;
        RECT 6.430 57.320 6.620 57.490 ;
        RECT 6.790 57.320 7.060 57.490 ;
        RECT 7.230 57.320 7.460 57.490 ;
        RECT 8.310 57.540 8.900 58.320 ;
        RECT 8.310 57.370 8.340 57.540 ;
        RECT 8.510 57.370 8.700 57.540 ;
        RECT 8.870 57.370 8.900 57.540 ;
        RECT 8.310 57.340 8.900 57.370 ;
        RECT 9.080 57.410 9.250 58.520 ;
        RECT 9.430 59.130 9.700 60.050 ;
        RECT 9.880 60.480 9.910 60.650 ;
        RECT 10.080 60.480 10.270 60.650 ;
        RECT 10.440 60.480 10.470 60.650 ;
        RECT 14.840 60.650 15.790 60.680 ;
        RECT 9.880 59.800 10.470 60.480 ;
      LAYER li1 ;
        RECT 10.750 60.420 13.690 60.590 ;
        RECT 10.750 59.430 10.920 60.420 ;
      LAYER li1 ;
        RECT 9.430 58.900 9.960 59.130 ;
        RECT 9.430 57.590 9.680 58.900 ;
      LAYER li1 ;
        RECT 10.380 58.560 10.920 59.430 ;
        RECT 11.100 58.940 11.430 60.240 ;
      LAYER li1 ;
        RECT 11.610 59.720 11.880 60.220 ;
        RECT 12.330 59.970 12.660 60.220 ;
        RECT 12.330 59.800 13.340 59.970 ;
        RECT 11.610 58.730 11.780 59.720 ;
        RECT 12.660 59.130 12.990 59.620 ;
        RECT 11.560 58.560 11.780 58.730 ;
        RECT 11.960 58.900 12.990 59.130 ;
        RECT 13.170 59.570 13.340 59.800 ;
      LAYER li1 ;
        RECT 13.520 59.920 13.690 60.420 ;
      LAYER li1 ;
        RECT 14.840 60.480 14.870 60.650 ;
        RECT 15.040 60.480 15.230 60.650 ;
        RECT 15.400 60.480 15.590 60.650 ;
        RECT 15.760 60.480 15.790 60.650 ;
        RECT 14.840 60.100 15.790 60.480 ;
      LAYER li1 ;
        RECT 15.970 60.610 18.630 60.780 ;
        RECT 15.970 59.920 16.140 60.610 ;
        RECT 13.520 59.750 16.140 59.920 ;
      LAYER li1 ;
        RECT 13.170 59.400 15.790 59.570 ;
        RECT 11.560 58.380 11.730 58.560 ;
        RECT 11.960 58.380 12.130 58.900 ;
        RECT 13.170 58.720 13.340 59.400 ;
      LAYER li1 ;
        RECT 15.970 59.220 16.140 59.750 ;
      LAYER li1 ;
        RECT 9.920 58.210 11.730 58.380 ;
        RECT 9.920 57.590 10.170 58.210 ;
        RECT 10.350 57.860 11.380 58.030 ;
        RECT 10.350 57.410 10.520 57.860 ;
        RECT 6.010 57.290 7.460 57.320 ;
        RECT 9.080 57.240 10.520 57.410 ;
        RECT 10.700 57.540 11.030 57.680 ;
        RECT 10.700 57.370 10.730 57.540 ;
        RECT 10.900 57.370 11.030 57.540 ;
        RECT 10.700 57.340 11.030 57.370 ;
        RECT 11.210 57.410 11.380 57.860 ;
        RECT 11.560 57.590 11.730 58.210 ;
        RECT 11.910 58.050 12.130 58.380 ;
        RECT 12.310 58.550 13.340 58.720 ;
        RECT 13.520 58.870 13.850 59.220 ;
      LAYER li1 ;
        RECT 14.290 59.050 16.140 59.220 ;
      LAYER li1 ;
        RECT 16.320 59.720 16.650 60.430 ;
        RECT 17.110 60.260 18.280 60.430 ;
        RECT 17.110 59.720 17.440 60.260 ;
        RECT 16.320 58.870 16.580 59.720 ;
        RECT 17.650 59.460 17.930 59.960 ;
        RECT 13.520 58.700 16.580 58.870 ;
        RECT 12.310 57.850 12.480 58.550 ;
        RECT 13.170 58.520 13.340 58.550 ;
        RECT 12.660 58.170 12.990 58.370 ;
        RECT 13.170 58.350 14.940 58.520 ;
        RECT 12.660 58.050 14.430 58.170 ;
        RECT 12.780 58.000 14.430 58.050 ;
        RECT 12.260 57.590 12.590 57.850 ;
        RECT 12.780 57.410 12.950 58.000 ;
        RECT 11.210 57.240 12.950 57.410 ;
        RECT 13.130 57.540 14.080 57.820 ;
        RECT 13.130 57.370 13.160 57.540 ;
        RECT 13.330 57.370 13.520 57.540 ;
        RECT 13.690 57.370 13.880 57.540 ;
        RECT 14.050 57.370 14.080 57.540 ;
        RECT 13.130 57.340 14.080 57.370 ;
        RECT 14.260 57.410 14.430 58.000 ;
        RECT 14.610 57.590 14.940 58.350 ;
        RECT 16.250 58.120 16.580 58.700 ;
        RECT 16.760 59.290 17.930 59.460 ;
        RECT 16.760 57.940 16.930 59.290 ;
        RECT 17.310 58.610 17.640 59.110 ;
        RECT 18.110 58.860 18.280 60.260 ;
      LAYER li1 ;
        RECT 18.460 59.950 18.630 60.610 ;
      LAYER li1 ;
        RECT 18.810 60.650 19.760 60.680 ;
        RECT 18.810 60.480 18.840 60.650 ;
        RECT 19.010 60.480 19.200 60.650 ;
        RECT 19.370 60.480 19.560 60.650 ;
        RECT 19.730 60.480 19.760 60.650 ;
        RECT 21.420 60.650 22.370 60.680 ;
        RECT 18.810 60.130 19.760 60.480 ;
        RECT 20.300 60.050 20.630 60.550 ;
        RECT 21.420 60.480 21.450 60.650 ;
        RECT 21.620 60.480 21.810 60.650 ;
        RECT 21.980 60.480 22.170 60.650 ;
        RECT 22.340 60.480 22.370 60.650 ;
      LAYER li1 ;
        RECT 18.460 59.840 19.470 59.950 ;
        RECT 18.460 59.780 19.520 59.840 ;
        RECT 19.140 59.670 19.520 59.780 ;
      LAYER li1 ;
        RECT 18.490 59.210 18.820 59.600 ;
      LAYER li1 ;
        RECT 19.140 59.390 19.470 59.670 ;
      LAYER li1 ;
        RECT 20.300 59.210 20.530 60.050 ;
        RECT 20.910 59.550 21.240 60.050 ;
        RECT 21.420 59.550 22.370 60.480 ;
        RECT 23.210 60.650 24.820 60.680 ;
        RECT 25.510 60.650 26.760 60.680 ;
        RECT 27.530 60.650 29.140 60.680 ;
        RECT 23.210 60.480 23.260 60.650 ;
        RECT 23.430 60.480 23.700 60.650 ;
        RECT 23.870 60.480 24.140 60.650 ;
        RECT 24.310 60.480 24.550 60.650 ;
        RECT 24.720 60.480 24.820 60.650 ;
        RECT 18.490 59.040 20.530 59.210 ;
        RECT 17.820 58.690 20.180 58.860 ;
        RECT 17.820 58.370 17.990 58.690 ;
        RECT 20.360 58.510 20.530 59.040 ;
        RECT 15.120 57.770 16.930 57.940 ;
        RECT 17.110 58.200 17.990 58.370 ;
        RECT 15.120 57.410 15.290 57.770 ;
        RECT 14.260 57.240 15.290 57.410 ;
        RECT 15.470 57.540 16.420 57.590 ;
        RECT 15.470 57.370 15.500 57.540 ;
        RECT 15.670 57.370 15.860 57.540 ;
        RECT 16.030 57.370 16.220 57.540 ;
        RECT 16.390 57.370 16.420 57.540 ;
        RECT 15.470 57.290 16.420 57.370 ;
        RECT 17.110 57.290 17.360 58.200 ;
        RECT 18.170 57.540 19.120 58.370 ;
        RECT 19.520 58.340 20.530 58.510 ;
        RECT 21.030 59.370 21.240 59.550 ;
        RECT 21.030 59.040 22.400 59.370 ;
        RECT 19.520 57.870 19.770 58.340 ;
        RECT 19.950 57.540 20.850 58.160 ;
        RECT 21.030 58.040 21.280 59.040 ;
        RECT 18.170 57.370 18.200 57.540 ;
        RECT 18.370 57.370 18.560 57.540 ;
        RECT 18.730 57.370 18.920 57.540 ;
        RECT 19.090 57.370 19.120 57.540 ;
        RECT 20.120 57.370 20.310 57.540 ;
        RECT 20.480 57.370 20.670 57.540 ;
        RECT 20.840 57.370 20.850 57.540 ;
        RECT 18.170 57.340 19.120 57.370 ;
        RECT 19.950 57.340 20.850 57.370 ;
        RECT 21.460 57.540 22.400 58.850 ;
        RECT 21.460 57.370 21.480 57.540 ;
        RECT 21.650 57.370 21.840 57.540 ;
        RECT 22.010 57.370 22.200 57.540 ;
        RECT 22.370 57.370 22.400 57.540 ;
        RECT 21.460 57.310 22.400 57.370 ;
      LAYER li1 ;
        RECT 22.580 57.310 22.920 60.380 ;
      LAYER li1 ;
        RECT 23.210 60.200 24.820 60.480 ;
        RECT 23.520 59.800 24.820 60.200 ;
        RECT 23.520 59.020 23.850 59.800 ;
        RECT 24.060 58.360 24.390 59.350 ;
      LAYER li1 ;
        RECT 25.080 58.870 25.330 60.550 ;
      LAYER li1 ;
        RECT 25.680 60.480 25.870 60.650 ;
        RECT 26.040 60.480 26.230 60.650 ;
        RECT 26.400 60.480 26.590 60.650 ;
        RECT 25.510 60.110 26.760 60.480 ;
        RECT 26.940 59.930 27.190 60.550 ;
        RECT 27.530 60.480 27.580 60.650 ;
        RECT 27.750 60.480 28.020 60.650 ;
        RECT 28.190 60.480 28.460 60.650 ;
        RECT 28.630 60.480 28.870 60.650 ;
        RECT 29.040 60.480 29.140 60.650 ;
        RECT 27.530 60.200 29.140 60.480 ;
        RECT 25.640 59.760 27.190 59.930 ;
        RECT 25.640 59.300 25.970 59.760 ;
        RECT 23.290 57.490 24.740 58.360 ;
        RECT 23.290 57.320 23.540 57.490 ;
        RECT 23.710 57.320 23.900 57.490 ;
        RECT 24.070 57.320 24.340 57.490 ;
        RECT 24.510 57.320 24.740 57.490 ;
        RECT 23.290 57.290 24.740 57.320 ;
      LAYER li1 ;
        RECT 25.080 57.290 25.510 58.870 ;
      LAYER li1 ;
        RECT 25.690 57.540 26.250 58.870 ;
      LAYER li1 ;
        RECT 26.430 57.790 26.760 59.580 ;
      LAYER li1 ;
        RECT 26.940 58.040 27.190 59.760 ;
        RECT 27.840 59.800 29.140 60.200 ;
        RECT 29.370 60.650 30.320 60.680 ;
        RECT 29.370 60.480 29.400 60.650 ;
        RECT 29.570 60.480 29.760 60.650 ;
        RECT 29.930 60.480 30.120 60.650 ;
        RECT 30.290 60.480 30.320 60.650 ;
        RECT 30.930 60.650 31.880 60.680 ;
        RECT 27.840 59.020 28.170 59.800 ;
        RECT 29.370 59.720 30.320 60.480 ;
      LAYER li1 ;
        RECT 30.500 59.840 30.750 60.550 ;
      LAYER li1 ;
        RECT 30.930 60.480 30.960 60.650 ;
        RECT 31.130 60.480 31.320 60.650 ;
        RECT 31.490 60.480 31.680 60.650 ;
        RECT 31.850 60.480 31.880 60.650 ;
        RECT 32.490 60.650 33.440 60.680 ;
        RECT 30.930 60.020 31.880 60.480 ;
      LAYER li1 ;
        RECT 32.060 59.840 32.310 60.550 ;
        RECT 30.500 59.670 32.310 59.840 ;
      LAYER li1 ;
        RECT 32.490 60.480 32.520 60.650 ;
        RECT 32.690 60.480 32.880 60.650 ;
        RECT 33.050 60.480 33.240 60.650 ;
        RECT 33.410 60.480 33.440 60.650 ;
        RECT 34.250 60.650 35.860 60.680 ;
        RECT 32.490 59.800 33.440 60.480 ;
      LAYER li1 ;
        RECT 30.500 59.500 30.670 59.670 ;
      LAYER li1 ;
        RECT 33.620 59.620 33.950 60.550 ;
        RECT 34.250 60.480 34.300 60.650 ;
        RECT 34.470 60.480 34.740 60.650 ;
        RECT 34.910 60.480 35.180 60.650 ;
        RECT 35.350 60.480 35.590 60.650 ;
        RECT 35.760 60.480 35.860 60.650 ;
        RECT 34.250 60.200 35.860 60.480 ;
        RECT 28.380 58.360 28.710 59.350 ;
      LAYER li1 ;
        RECT 29.410 59.270 30.670 59.500 ;
      LAYER li1 ;
        RECT 32.710 59.490 33.950 59.620 ;
        RECT 30.850 59.450 33.950 59.490 ;
        RECT 30.850 59.320 32.880 59.450 ;
      LAYER li1 ;
        RECT 30.500 59.140 30.670 59.270 ;
        RECT 30.500 58.970 32.390 59.140 ;
      LAYER li1 ;
        RECT 25.690 57.370 25.700 57.540 ;
        RECT 25.870 57.370 26.060 57.540 ;
        RECT 26.230 57.370 26.250 57.540 ;
        RECT 25.690 57.290 26.250 57.370 ;
        RECT 27.610 57.490 29.060 58.360 ;
        RECT 27.610 57.320 27.860 57.490 ;
        RECT 28.030 57.320 28.220 57.490 ;
        RECT 28.390 57.320 28.660 57.490 ;
        RECT 28.830 57.320 29.060 57.490 ;
        RECT 27.610 57.290 29.060 57.320 ;
        RECT 29.370 57.540 30.320 58.870 ;
        RECT 29.370 57.370 29.400 57.540 ;
        RECT 29.570 57.370 29.760 57.540 ;
        RECT 29.930 57.370 30.120 57.540 ;
        RECT 30.290 57.370 30.320 57.540 ;
        RECT 29.370 57.290 30.320 57.370 ;
      LAYER li1 ;
        RECT 30.500 57.290 30.750 58.970 ;
      LAYER li1 ;
        RECT 30.930 57.540 31.880 58.790 ;
        RECT 30.930 57.370 30.960 57.540 ;
        RECT 31.130 57.370 31.320 57.540 ;
        RECT 31.490 57.370 31.680 57.540 ;
        RECT 31.850 57.370 31.880 57.540 ;
        RECT 30.930 57.290 31.880 57.370 ;
      LAYER li1 ;
        RECT 32.060 57.290 32.390 58.970 ;
        RECT 33.170 58.930 33.500 59.270 ;
      LAYER li1 ;
        RECT 32.570 57.540 33.520 58.750 ;
        RECT 32.570 57.370 32.600 57.540 ;
        RECT 32.770 57.370 32.960 57.540 ;
        RECT 33.130 57.370 33.320 57.540 ;
        RECT 33.490 57.370 33.520 57.540 ;
        RECT 32.570 57.290 33.520 57.370 ;
        RECT 33.700 57.290 33.950 59.450 ;
        RECT 34.560 59.800 35.860 60.200 ;
        RECT 36.090 60.650 37.040 60.680 ;
        RECT 36.090 60.480 36.120 60.650 ;
        RECT 36.290 60.480 36.480 60.650 ;
        RECT 36.650 60.480 36.840 60.650 ;
        RECT 37.010 60.480 37.040 60.650 ;
        RECT 37.650 60.650 38.600 60.680 ;
        RECT 34.560 59.020 34.890 59.800 ;
        RECT 36.090 59.720 37.040 60.480 ;
      LAYER li1 ;
        RECT 37.220 59.840 37.470 60.550 ;
      LAYER li1 ;
        RECT 37.650 60.480 37.680 60.650 ;
        RECT 37.850 60.480 38.040 60.650 ;
        RECT 38.210 60.480 38.400 60.650 ;
        RECT 38.570 60.480 38.600 60.650 ;
        RECT 39.210 60.650 40.160 60.680 ;
        RECT 37.650 60.020 38.600 60.480 ;
      LAYER li1 ;
        RECT 38.780 59.840 39.030 60.550 ;
        RECT 37.220 59.670 39.030 59.840 ;
      LAYER li1 ;
        RECT 39.210 60.480 39.240 60.650 ;
        RECT 39.410 60.480 39.600 60.650 ;
        RECT 39.770 60.480 39.960 60.650 ;
        RECT 40.130 60.480 40.160 60.650 ;
        RECT 40.970 60.650 42.580 60.680 ;
        RECT 39.210 59.800 40.160 60.480 ;
      LAYER li1 ;
        RECT 37.220 59.500 37.390 59.670 ;
      LAYER li1 ;
        RECT 40.340 59.620 40.670 60.550 ;
        RECT 40.970 60.480 41.020 60.650 ;
        RECT 41.190 60.480 41.460 60.650 ;
        RECT 41.630 60.480 41.900 60.650 ;
        RECT 42.070 60.480 42.310 60.650 ;
        RECT 42.480 60.480 42.580 60.650 ;
        RECT 40.970 60.200 42.580 60.480 ;
        RECT 35.100 58.360 35.430 59.350 ;
      LAYER li1 ;
        RECT 36.130 59.270 37.390 59.500 ;
      LAYER li1 ;
        RECT 39.430 59.490 40.670 59.620 ;
        RECT 37.570 59.450 40.670 59.490 ;
        RECT 37.570 59.320 39.600 59.450 ;
      LAYER li1 ;
        RECT 37.220 59.140 37.390 59.270 ;
        RECT 37.220 58.970 39.110 59.140 ;
      LAYER li1 ;
        RECT 34.330 57.490 35.780 58.360 ;
        RECT 34.330 57.320 34.580 57.490 ;
        RECT 34.750 57.320 34.940 57.490 ;
        RECT 35.110 57.320 35.380 57.490 ;
        RECT 35.550 57.320 35.780 57.490 ;
        RECT 34.330 57.290 35.780 57.320 ;
        RECT 36.090 57.540 37.040 58.870 ;
        RECT 36.090 57.370 36.120 57.540 ;
        RECT 36.290 57.370 36.480 57.540 ;
        RECT 36.650 57.370 36.840 57.540 ;
        RECT 37.010 57.370 37.040 57.540 ;
        RECT 36.090 57.290 37.040 57.370 ;
      LAYER li1 ;
        RECT 37.220 57.290 37.470 58.970 ;
      LAYER li1 ;
        RECT 37.650 57.540 38.600 58.790 ;
        RECT 37.650 57.370 37.680 57.540 ;
        RECT 37.850 57.370 38.040 57.540 ;
        RECT 38.210 57.370 38.400 57.540 ;
        RECT 38.570 57.370 38.600 57.540 ;
        RECT 37.650 57.290 38.600 57.370 ;
      LAYER li1 ;
        RECT 38.780 57.290 39.110 58.970 ;
        RECT 39.890 58.930 40.220 59.270 ;
      LAYER li1 ;
        RECT 39.290 57.540 40.240 58.750 ;
        RECT 39.290 57.370 39.320 57.540 ;
        RECT 39.490 57.370 39.680 57.540 ;
        RECT 39.850 57.370 40.040 57.540 ;
        RECT 40.210 57.370 40.240 57.540 ;
        RECT 39.290 57.290 40.240 57.370 ;
        RECT 40.420 57.290 40.670 59.450 ;
        RECT 41.280 59.800 42.580 60.200 ;
        RECT 42.810 60.650 43.760 60.680 ;
        RECT 42.810 60.480 42.840 60.650 ;
        RECT 43.010 60.480 43.200 60.650 ;
        RECT 43.370 60.480 43.560 60.650 ;
        RECT 43.730 60.480 43.760 60.650 ;
        RECT 44.370 60.650 45.320 60.680 ;
        RECT 41.280 59.020 41.610 59.800 ;
        RECT 42.810 59.720 43.760 60.480 ;
      LAYER li1 ;
        RECT 43.940 59.840 44.190 60.550 ;
      LAYER li1 ;
        RECT 44.370 60.480 44.400 60.650 ;
        RECT 44.570 60.480 44.760 60.650 ;
        RECT 44.930 60.480 45.120 60.650 ;
        RECT 45.290 60.480 45.320 60.650 ;
        RECT 45.930 60.650 46.880 60.680 ;
        RECT 44.370 60.020 45.320 60.480 ;
      LAYER li1 ;
        RECT 45.500 59.840 45.750 60.550 ;
        RECT 43.940 59.670 45.750 59.840 ;
      LAYER li1 ;
        RECT 45.930 60.480 45.960 60.650 ;
        RECT 46.130 60.480 46.320 60.650 ;
        RECT 46.490 60.480 46.680 60.650 ;
        RECT 46.850 60.480 46.880 60.650 ;
        RECT 47.690 60.650 49.300 60.680 ;
        RECT 45.930 59.800 46.880 60.480 ;
      LAYER li1 ;
        RECT 43.940 59.500 44.110 59.670 ;
      LAYER li1 ;
        RECT 47.060 59.620 47.390 60.550 ;
        RECT 47.690 60.480 47.740 60.650 ;
        RECT 47.910 60.480 48.180 60.650 ;
        RECT 48.350 60.480 48.620 60.650 ;
        RECT 48.790 60.480 49.030 60.650 ;
        RECT 49.200 60.480 49.300 60.650 ;
        RECT 47.690 60.200 49.300 60.480 ;
        RECT 41.820 58.360 42.150 59.350 ;
      LAYER li1 ;
        RECT 42.850 59.270 44.110 59.500 ;
      LAYER li1 ;
        RECT 46.150 59.490 47.390 59.620 ;
        RECT 44.290 59.450 47.390 59.490 ;
        RECT 44.290 59.320 46.320 59.450 ;
      LAYER li1 ;
        RECT 43.940 59.140 44.110 59.270 ;
        RECT 43.940 58.970 45.830 59.140 ;
      LAYER li1 ;
        RECT 41.050 57.490 42.500 58.360 ;
        RECT 41.050 57.320 41.300 57.490 ;
        RECT 41.470 57.320 41.660 57.490 ;
        RECT 41.830 57.320 42.100 57.490 ;
        RECT 42.270 57.320 42.500 57.490 ;
        RECT 41.050 57.290 42.500 57.320 ;
        RECT 42.810 57.540 43.760 58.870 ;
        RECT 42.810 57.370 42.840 57.540 ;
        RECT 43.010 57.370 43.200 57.540 ;
        RECT 43.370 57.370 43.560 57.540 ;
        RECT 43.730 57.370 43.760 57.540 ;
        RECT 42.810 57.290 43.760 57.370 ;
      LAYER li1 ;
        RECT 43.940 57.290 44.190 58.970 ;
      LAYER li1 ;
        RECT 44.370 57.540 45.320 58.790 ;
        RECT 44.370 57.370 44.400 57.540 ;
        RECT 44.570 57.370 44.760 57.540 ;
        RECT 44.930 57.370 45.120 57.540 ;
        RECT 45.290 57.370 45.320 57.540 ;
        RECT 44.370 57.290 45.320 57.370 ;
      LAYER li1 ;
        RECT 45.500 57.290 45.830 58.970 ;
        RECT 46.610 58.930 46.940 59.270 ;
      LAYER li1 ;
        RECT 46.010 57.540 46.960 58.750 ;
        RECT 46.010 57.370 46.040 57.540 ;
        RECT 46.210 57.370 46.400 57.540 ;
        RECT 46.570 57.370 46.760 57.540 ;
        RECT 46.930 57.370 46.960 57.540 ;
        RECT 46.010 57.290 46.960 57.370 ;
        RECT 47.140 57.290 47.390 59.450 ;
        RECT 48.000 59.800 49.300 60.200 ;
        RECT 50.010 60.650 50.960 60.680 ;
        RECT 50.010 60.480 50.040 60.650 ;
        RECT 50.210 60.480 50.400 60.650 ;
        RECT 50.570 60.480 50.760 60.650 ;
        RECT 50.930 60.480 50.960 60.650 ;
        RECT 51.570 60.650 52.520 60.680 ;
        RECT 48.000 59.020 48.330 59.800 ;
        RECT 50.010 59.720 50.960 60.480 ;
      LAYER li1 ;
        RECT 51.140 59.840 51.390 60.550 ;
      LAYER li1 ;
        RECT 51.570 60.480 51.600 60.650 ;
        RECT 51.770 60.480 51.960 60.650 ;
        RECT 52.130 60.480 52.320 60.650 ;
        RECT 52.490 60.480 52.520 60.650 ;
        RECT 53.130 60.650 54.080 60.680 ;
        RECT 51.570 60.020 52.520 60.480 ;
      LAYER li1 ;
        RECT 52.700 59.840 52.950 60.550 ;
        RECT 51.140 59.670 52.950 59.840 ;
      LAYER li1 ;
        RECT 53.130 60.480 53.160 60.650 ;
        RECT 53.330 60.480 53.520 60.650 ;
        RECT 53.690 60.480 53.880 60.650 ;
        RECT 54.050 60.480 54.080 60.650 ;
        RECT 54.890 60.650 56.500 60.680 ;
        RECT 53.130 59.800 54.080 60.480 ;
      LAYER li1 ;
        RECT 51.140 59.500 51.310 59.670 ;
      LAYER li1 ;
        RECT 54.260 59.620 54.590 60.550 ;
        RECT 54.890 60.480 54.940 60.650 ;
        RECT 55.110 60.480 55.380 60.650 ;
        RECT 55.550 60.480 55.820 60.650 ;
        RECT 55.990 60.480 56.230 60.650 ;
        RECT 56.400 60.480 56.500 60.650 ;
        RECT 54.890 60.200 56.500 60.480 ;
        RECT 48.540 58.360 48.870 59.350 ;
      LAYER li1 ;
        RECT 50.050 59.270 51.310 59.500 ;
      LAYER li1 ;
        RECT 53.350 59.490 54.590 59.620 ;
        RECT 51.490 59.450 54.590 59.490 ;
        RECT 51.490 59.320 53.520 59.450 ;
      LAYER li1 ;
        RECT 51.140 59.140 51.310 59.270 ;
        RECT 51.140 58.970 53.030 59.140 ;
      LAYER li1 ;
        RECT 47.770 57.490 49.220 58.360 ;
        RECT 47.770 57.320 48.020 57.490 ;
        RECT 48.190 57.320 48.380 57.490 ;
        RECT 48.550 57.320 48.820 57.490 ;
        RECT 48.990 57.320 49.220 57.490 ;
        RECT 47.770 57.290 49.220 57.320 ;
        RECT 50.010 57.540 50.960 58.870 ;
        RECT 50.010 57.370 50.040 57.540 ;
        RECT 50.210 57.370 50.400 57.540 ;
        RECT 50.570 57.370 50.760 57.540 ;
        RECT 50.930 57.370 50.960 57.540 ;
        RECT 50.010 57.290 50.960 57.370 ;
      LAYER li1 ;
        RECT 51.140 57.290 51.390 58.970 ;
      LAYER li1 ;
        RECT 51.570 57.540 52.520 58.790 ;
        RECT 51.570 57.370 51.600 57.540 ;
        RECT 51.770 57.370 51.960 57.540 ;
        RECT 52.130 57.370 52.320 57.540 ;
        RECT 52.490 57.370 52.520 57.540 ;
        RECT 51.570 57.290 52.520 57.370 ;
      LAYER li1 ;
        RECT 52.700 57.290 53.030 58.970 ;
        RECT 53.810 58.930 54.140 59.270 ;
      LAYER li1 ;
        RECT 53.210 57.540 54.160 58.750 ;
        RECT 53.210 57.370 53.240 57.540 ;
        RECT 53.410 57.370 53.600 57.540 ;
        RECT 53.770 57.370 53.960 57.540 ;
        RECT 54.130 57.370 54.160 57.540 ;
        RECT 53.210 57.290 54.160 57.370 ;
        RECT 54.340 57.290 54.590 59.450 ;
        RECT 55.200 59.800 56.500 60.200 ;
        RECT 56.730 60.650 57.320 60.680 ;
        RECT 56.730 60.480 56.760 60.650 ;
        RECT 56.930 60.480 57.120 60.650 ;
        RECT 57.290 60.480 57.320 60.650 ;
        RECT 58.000 60.650 58.950 60.680 ;
        RECT 55.200 59.020 55.530 59.800 ;
        RECT 56.730 59.720 57.320 60.480 ;
      LAYER li1 ;
        RECT 57.570 59.620 57.820 60.550 ;
      LAYER li1 ;
        RECT 58.000 60.480 58.030 60.650 ;
        RECT 58.200 60.480 58.390 60.650 ;
        RECT 58.560 60.480 58.750 60.650 ;
        RECT 58.920 60.480 58.950 60.650 ;
        RECT 60.170 60.650 61.780 60.680 ;
        RECT 58.000 59.800 58.950 60.480 ;
      LAYER li1 ;
        RECT 59.130 59.620 59.400 60.550 ;
      LAYER li1 ;
        RECT 60.170 60.480 60.220 60.650 ;
        RECT 60.390 60.480 60.660 60.650 ;
        RECT 60.830 60.480 61.100 60.650 ;
        RECT 61.270 60.480 61.510 60.650 ;
        RECT 61.680 60.480 61.780 60.650 ;
        RECT 62.480 60.650 63.430 60.680 ;
        RECT 60.170 60.200 61.780 60.480 ;
        RECT 55.740 58.360 56.070 59.350 ;
      LAYER li1 ;
        RECT 56.770 58.930 57.070 59.520 ;
        RECT 57.570 59.450 59.400 59.620 ;
        RECT 57.250 58.930 58.440 59.270 ;
      LAYER li1 ;
        RECT 54.970 57.490 56.420 58.360 ;
        RECT 54.970 57.320 55.220 57.490 ;
        RECT 55.390 57.320 55.580 57.490 ;
        RECT 55.750 57.320 56.020 57.490 ;
        RECT 56.190 57.320 56.420 57.490 ;
        RECT 54.970 57.290 56.420 57.320 ;
        RECT 56.730 57.540 58.400 58.750 ;
      LAYER li1 ;
        RECT 58.620 57.790 58.950 59.270 ;
      LAYER li1 ;
        RECT 56.730 57.370 56.760 57.540 ;
        RECT 56.930 57.370 57.120 57.540 ;
        RECT 57.290 57.370 57.480 57.540 ;
        RECT 57.650 57.370 57.840 57.540 ;
        RECT 58.010 57.370 58.200 57.540 ;
        RECT 58.370 57.370 58.400 57.540 ;
        RECT 56.730 57.290 58.400 57.370 ;
      LAYER li1 ;
        RECT 59.130 57.290 59.400 59.450 ;
      LAYER li1 ;
        RECT 60.480 59.800 61.780 60.200 ;
        RECT 60.480 59.020 60.810 59.800 ;
        RECT 61.020 58.360 61.350 59.350 ;
        RECT 62.030 58.690 62.300 60.550 ;
        RECT 62.480 60.480 62.510 60.650 ;
        RECT 62.680 60.480 62.870 60.650 ;
        RECT 63.040 60.480 63.230 60.650 ;
        RECT 63.400 60.480 63.430 60.650 ;
        RECT 64.120 60.650 64.710 60.680 ;
        RECT 62.480 60.050 63.430 60.480 ;
        RECT 63.610 60.050 63.940 60.550 ;
        RECT 63.160 58.690 63.490 59.190 ;
        RECT 62.030 58.520 63.490 58.690 ;
        RECT 60.250 57.490 61.700 58.360 ;
        RECT 62.030 57.590 62.360 58.520 ;
        RECT 60.250 57.320 60.500 57.490 ;
        RECT 60.670 57.320 60.860 57.490 ;
        RECT 61.030 57.320 61.300 57.490 ;
        RECT 61.470 57.320 61.700 57.490 ;
        RECT 62.550 57.540 63.140 58.320 ;
        RECT 62.550 57.370 62.580 57.540 ;
        RECT 62.750 57.370 62.940 57.540 ;
        RECT 63.110 57.370 63.140 57.540 ;
        RECT 62.550 57.340 63.140 57.370 ;
        RECT 63.320 57.410 63.490 58.520 ;
        RECT 63.670 59.130 63.940 60.050 ;
        RECT 64.120 60.480 64.150 60.650 ;
        RECT 64.320 60.480 64.510 60.650 ;
        RECT 64.680 60.480 64.710 60.650 ;
        RECT 69.080 60.650 70.030 60.680 ;
        RECT 64.120 59.800 64.710 60.480 ;
      LAYER li1 ;
        RECT 64.990 60.420 67.930 60.590 ;
        RECT 64.990 60.210 65.160 60.420 ;
        RECT 64.950 60.040 65.160 60.210 ;
        RECT 64.990 59.430 65.160 60.040 ;
      LAYER li1 ;
        RECT 63.670 58.900 64.200 59.130 ;
        RECT 63.670 57.590 63.920 58.900 ;
      LAYER li1 ;
        RECT 64.620 58.560 65.160 59.430 ;
        RECT 65.340 58.940 65.670 60.240 ;
      LAYER li1 ;
        RECT 65.850 59.720 66.120 60.220 ;
        RECT 66.570 59.970 66.900 60.220 ;
        RECT 66.570 59.800 67.580 59.970 ;
        RECT 65.850 58.730 66.020 59.720 ;
        RECT 66.900 59.130 67.230 59.620 ;
        RECT 65.800 58.560 66.020 58.730 ;
        RECT 66.200 58.900 67.230 59.130 ;
        RECT 67.410 59.570 67.580 59.800 ;
      LAYER li1 ;
        RECT 67.760 59.920 67.930 60.420 ;
      LAYER li1 ;
        RECT 69.080 60.480 69.110 60.650 ;
        RECT 69.280 60.480 69.470 60.650 ;
        RECT 69.640 60.480 69.830 60.650 ;
        RECT 70.000 60.480 70.030 60.650 ;
        RECT 69.080 60.100 70.030 60.480 ;
      LAYER li1 ;
        RECT 70.210 60.610 72.870 60.780 ;
        RECT 70.210 59.920 70.380 60.610 ;
        RECT 67.760 59.750 70.380 59.920 ;
      LAYER li1 ;
        RECT 67.410 59.400 70.030 59.570 ;
        RECT 65.800 58.380 65.970 58.560 ;
        RECT 66.200 58.380 66.370 58.900 ;
        RECT 67.410 58.720 67.580 59.400 ;
      LAYER li1 ;
        RECT 70.210 59.220 70.380 59.750 ;
      LAYER li1 ;
        RECT 64.160 58.210 65.970 58.380 ;
        RECT 64.160 57.590 64.410 58.210 ;
        RECT 64.590 57.860 65.620 58.030 ;
        RECT 64.590 57.410 64.760 57.860 ;
        RECT 60.250 57.290 61.700 57.320 ;
        RECT 63.320 57.240 64.760 57.410 ;
        RECT 64.940 57.540 65.270 57.680 ;
        RECT 64.940 57.370 64.970 57.540 ;
        RECT 65.140 57.370 65.270 57.540 ;
        RECT 64.940 57.340 65.270 57.370 ;
        RECT 65.450 57.410 65.620 57.860 ;
        RECT 65.800 57.590 65.970 58.210 ;
        RECT 66.150 58.050 66.370 58.380 ;
        RECT 66.550 58.550 67.580 58.720 ;
        RECT 67.760 58.870 68.090 59.220 ;
      LAYER li1 ;
        RECT 68.530 59.050 70.380 59.220 ;
      LAYER li1 ;
        RECT 70.560 59.720 70.890 60.430 ;
        RECT 71.350 60.260 72.520 60.430 ;
        RECT 71.350 59.720 71.680 60.260 ;
        RECT 70.560 58.870 70.820 59.720 ;
        RECT 71.890 59.460 72.170 59.960 ;
        RECT 67.760 58.700 70.820 58.870 ;
        RECT 66.550 57.850 66.720 58.550 ;
        RECT 67.410 58.520 67.580 58.550 ;
        RECT 66.900 58.170 67.230 58.370 ;
        RECT 67.410 58.350 69.180 58.520 ;
        RECT 66.900 58.050 68.670 58.170 ;
        RECT 67.020 58.000 68.670 58.050 ;
        RECT 66.500 57.590 66.830 57.850 ;
        RECT 67.020 57.410 67.190 58.000 ;
        RECT 65.450 57.240 67.190 57.410 ;
        RECT 67.370 57.540 68.320 57.820 ;
        RECT 67.370 57.370 67.400 57.540 ;
        RECT 67.570 57.370 67.760 57.540 ;
        RECT 67.930 57.370 68.120 57.540 ;
        RECT 68.290 57.370 68.320 57.540 ;
        RECT 67.370 57.340 68.320 57.370 ;
        RECT 68.500 57.410 68.670 58.000 ;
        RECT 68.850 57.590 69.180 58.350 ;
        RECT 70.490 58.120 70.820 58.700 ;
        RECT 71.000 59.290 72.170 59.460 ;
        RECT 71.000 57.940 71.170 59.290 ;
        RECT 71.550 58.610 71.880 59.110 ;
        RECT 72.350 58.860 72.520 60.260 ;
      LAYER li1 ;
        RECT 72.700 59.950 72.870 60.610 ;
      LAYER li1 ;
        RECT 73.050 60.650 74.000 60.680 ;
        RECT 73.050 60.480 73.080 60.650 ;
        RECT 73.250 60.480 73.440 60.650 ;
        RECT 73.610 60.480 73.800 60.650 ;
        RECT 73.970 60.480 74.000 60.650 ;
        RECT 75.660 60.650 76.610 60.680 ;
        RECT 73.050 60.130 74.000 60.480 ;
        RECT 74.540 60.050 74.870 60.550 ;
        RECT 75.660 60.480 75.690 60.650 ;
        RECT 75.860 60.480 76.050 60.650 ;
        RECT 76.220 60.480 76.410 60.650 ;
        RECT 76.580 60.480 76.610 60.650 ;
      LAYER li1 ;
        RECT 72.700 59.780 73.710 59.950 ;
      LAYER li1 ;
        RECT 72.730 59.210 73.060 59.600 ;
      LAYER li1 ;
        RECT 73.380 59.390 73.710 59.780 ;
      LAYER li1 ;
        RECT 74.540 59.210 74.770 60.050 ;
        RECT 75.150 59.550 75.480 60.050 ;
        RECT 75.660 59.550 76.610 60.480 ;
        RECT 77.450 60.650 79.060 60.680 ;
        RECT 77.450 60.480 77.500 60.650 ;
        RECT 77.670 60.480 77.940 60.650 ;
        RECT 78.110 60.480 78.380 60.650 ;
        RECT 78.550 60.480 78.790 60.650 ;
        RECT 78.960 60.480 79.060 60.650 ;
        RECT 72.730 59.040 74.770 59.210 ;
        RECT 72.060 58.690 74.420 58.860 ;
        RECT 72.060 58.370 72.230 58.690 ;
        RECT 74.600 58.510 74.770 59.040 ;
        RECT 69.360 57.770 71.170 57.940 ;
        RECT 71.350 58.200 72.230 58.370 ;
        RECT 69.360 57.410 69.530 57.770 ;
        RECT 68.500 57.240 69.530 57.410 ;
        RECT 69.710 57.540 70.660 57.590 ;
        RECT 69.710 57.370 69.740 57.540 ;
        RECT 69.910 57.370 70.100 57.540 ;
        RECT 70.270 57.370 70.460 57.540 ;
        RECT 70.630 57.370 70.660 57.540 ;
        RECT 69.710 57.290 70.660 57.370 ;
        RECT 71.350 57.290 71.600 58.200 ;
        RECT 72.410 57.540 73.360 58.370 ;
        RECT 73.760 58.340 74.770 58.510 ;
        RECT 75.270 59.370 75.480 59.550 ;
        RECT 75.270 59.040 76.640 59.370 ;
        RECT 73.760 57.870 74.010 58.340 ;
        RECT 74.190 57.540 75.090 58.160 ;
        RECT 75.270 58.040 75.520 59.040 ;
        RECT 72.410 57.370 72.440 57.540 ;
        RECT 72.610 57.370 72.800 57.540 ;
        RECT 72.970 57.370 73.160 57.540 ;
        RECT 73.330 57.370 73.360 57.540 ;
        RECT 74.360 57.370 74.550 57.540 ;
        RECT 74.720 57.370 74.910 57.540 ;
        RECT 75.080 57.370 75.090 57.540 ;
        RECT 72.410 57.340 73.360 57.370 ;
        RECT 74.190 57.340 75.090 57.370 ;
        RECT 75.700 57.540 76.640 58.850 ;
        RECT 75.700 57.370 75.720 57.540 ;
        RECT 75.890 57.370 76.080 57.540 ;
        RECT 76.250 57.370 76.440 57.540 ;
        RECT 76.610 57.370 76.640 57.540 ;
        RECT 75.700 57.310 76.640 57.370 ;
      LAYER li1 ;
        RECT 76.820 57.310 77.160 60.380 ;
      LAYER li1 ;
        RECT 77.450 60.200 79.060 60.480 ;
        RECT 77.760 59.800 79.060 60.200 ;
        RECT 79.290 60.650 80.240 60.680 ;
        RECT 79.290 60.480 79.320 60.650 ;
        RECT 79.490 60.480 79.680 60.650 ;
        RECT 79.850 60.480 80.040 60.650 ;
        RECT 80.210 60.480 80.240 60.650 ;
        RECT 80.850 60.650 81.800 60.680 ;
        RECT 77.760 59.020 78.090 59.800 ;
        RECT 79.290 59.720 80.240 60.480 ;
      LAYER li1 ;
        RECT 80.420 59.840 80.670 60.550 ;
      LAYER li1 ;
        RECT 80.850 60.480 80.880 60.650 ;
        RECT 81.050 60.480 81.240 60.650 ;
        RECT 81.410 60.480 81.600 60.650 ;
        RECT 81.770 60.480 81.800 60.650 ;
        RECT 82.410 60.650 83.360 60.680 ;
        RECT 80.850 60.020 81.800 60.480 ;
      LAYER li1 ;
        RECT 81.980 59.840 82.230 60.550 ;
        RECT 80.420 59.670 82.230 59.840 ;
      LAYER li1 ;
        RECT 82.410 60.480 82.440 60.650 ;
        RECT 82.610 60.480 82.800 60.650 ;
        RECT 82.970 60.480 83.160 60.650 ;
        RECT 83.330 60.480 83.360 60.650 ;
        RECT 84.580 60.660 87.310 60.690 ;
        RECT 82.410 59.800 83.360 60.480 ;
      LAYER li1 ;
        RECT 80.420 59.500 80.590 59.670 ;
      LAYER li1 ;
        RECT 83.540 59.620 83.870 60.550 ;
        RECT 84.580 60.490 84.750 60.660 ;
        RECT 84.920 60.490 85.190 60.660 ;
        RECT 85.360 60.490 85.600 60.660 ;
        RECT 85.770 60.490 86.030 60.660 ;
        RECT 86.200 60.490 86.470 60.660 ;
        RECT 86.640 60.490 86.880 60.660 ;
        RECT 87.050 60.490 87.310 60.660 ;
        RECT 84.580 59.690 87.310 60.490 ;
        RECT 87.930 60.650 88.880 60.680 ;
        RECT 87.930 60.480 87.960 60.650 ;
        RECT 88.130 60.480 88.320 60.650 ;
        RECT 88.490 60.480 88.680 60.650 ;
        RECT 88.850 60.480 88.880 60.650 ;
        RECT 89.490 60.650 90.440 60.680 ;
        RECT 87.930 59.720 88.880 60.480 ;
      LAYER li1 ;
        RECT 89.060 59.840 89.310 60.550 ;
      LAYER li1 ;
        RECT 89.490 60.480 89.520 60.650 ;
        RECT 89.690 60.480 89.880 60.650 ;
        RECT 90.050 60.480 90.240 60.650 ;
        RECT 90.410 60.480 90.440 60.650 ;
        RECT 91.050 60.650 92.000 60.680 ;
        RECT 89.490 60.020 90.440 60.480 ;
      LAYER li1 ;
        RECT 90.620 59.840 90.870 60.550 ;
      LAYER li1 ;
        RECT 78.300 58.360 78.630 59.350 ;
      LAYER li1 ;
        RECT 79.330 59.270 80.590 59.500 ;
      LAYER li1 ;
        RECT 82.630 59.490 83.870 59.620 ;
        RECT 80.770 59.450 83.870 59.490 ;
        RECT 80.770 59.320 82.800 59.450 ;
      LAYER li1 ;
        RECT 80.420 59.140 80.590 59.270 ;
        RECT 80.420 58.970 82.310 59.140 ;
      LAYER li1 ;
        RECT 77.530 57.490 78.980 58.360 ;
        RECT 77.530 57.320 77.780 57.490 ;
        RECT 77.950 57.320 78.140 57.490 ;
        RECT 78.310 57.320 78.580 57.490 ;
        RECT 78.750 57.320 78.980 57.490 ;
        RECT 77.530 57.290 78.980 57.320 ;
        RECT 79.290 57.540 80.240 58.870 ;
        RECT 79.290 57.370 79.320 57.540 ;
        RECT 79.490 57.370 79.680 57.540 ;
        RECT 79.850 57.370 80.040 57.540 ;
        RECT 80.210 57.370 80.240 57.540 ;
        RECT 79.290 57.290 80.240 57.370 ;
      LAYER li1 ;
        RECT 80.420 57.290 80.670 58.970 ;
      LAYER li1 ;
        RECT 80.850 57.540 81.800 58.790 ;
        RECT 80.850 57.370 80.880 57.540 ;
        RECT 81.050 57.370 81.240 57.540 ;
        RECT 81.410 57.370 81.600 57.540 ;
        RECT 81.770 57.370 81.800 57.540 ;
        RECT 80.850 57.290 81.800 57.370 ;
      LAYER li1 ;
        RECT 81.980 57.290 82.310 58.970 ;
        RECT 83.090 58.930 83.420 59.270 ;
      LAYER li1 ;
        RECT 82.490 57.540 83.440 58.750 ;
        RECT 82.490 57.370 82.520 57.540 ;
        RECT 82.690 57.370 82.880 57.540 ;
        RECT 83.050 57.370 83.240 57.540 ;
        RECT 83.410 57.370 83.440 57.540 ;
        RECT 82.490 57.290 83.440 57.370 ;
        RECT 83.620 57.290 83.870 59.450 ;
        RECT 84.740 59.020 85.070 59.690 ;
        RECT 85.470 58.370 85.800 59.350 ;
        RECT 86.020 59.020 86.350 59.690 ;
      LAYER li1 ;
        RECT 89.060 59.670 90.870 59.840 ;
      LAYER li1 ;
        RECT 91.050 60.480 91.080 60.650 ;
        RECT 91.250 60.480 91.440 60.650 ;
        RECT 91.610 60.480 91.800 60.650 ;
        RECT 91.970 60.480 92.000 60.650 ;
        RECT 92.810 60.650 94.420 60.680 ;
        RECT 91.050 59.800 92.000 60.480 ;
      LAYER li1 ;
        RECT 89.060 59.500 89.230 59.670 ;
      LAYER li1 ;
        RECT 92.180 59.620 92.510 60.550 ;
        RECT 92.810 60.480 92.860 60.650 ;
        RECT 93.030 60.480 93.300 60.650 ;
        RECT 93.470 60.480 93.740 60.650 ;
        RECT 93.910 60.480 94.150 60.650 ;
        RECT 94.320 60.480 94.420 60.650 ;
        RECT 92.810 60.200 94.420 60.480 ;
        RECT 86.750 58.370 87.080 59.350 ;
      LAYER li1 ;
        RECT 87.970 59.270 89.230 59.500 ;
      LAYER li1 ;
        RECT 91.270 59.490 92.510 59.620 ;
        RECT 89.410 59.450 92.510 59.490 ;
        RECT 89.410 59.320 91.440 59.450 ;
      LAYER li1 ;
        RECT 89.060 59.140 89.230 59.270 ;
        RECT 89.060 58.970 90.950 59.140 ;
      LAYER li1 ;
        RECT 84.500 57.490 87.240 58.370 ;
        RECT 84.500 57.320 84.710 57.490 ;
        RECT 84.880 57.320 85.150 57.490 ;
        RECT 85.320 57.320 85.560 57.490 ;
        RECT 85.730 57.320 85.990 57.490 ;
        RECT 86.160 57.320 86.430 57.490 ;
        RECT 86.600 57.320 86.840 57.490 ;
        RECT 87.010 57.320 87.240 57.490 ;
        RECT 84.500 57.300 87.240 57.320 ;
        RECT 87.930 57.540 88.880 58.870 ;
        RECT 87.930 57.370 87.960 57.540 ;
        RECT 88.130 57.370 88.320 57.540 ;
        RECT 88.490 57.370 88.680 57.540 ;
        RECT 88.850 57.370 88.880 57.540 ;
        RECT 87.930 57.290 88.880 57.370 ;
      LAYER li1 ;
        RECT 89.060 57.290 89.310 58.970 ;
      LAYER li1 ;
        RECT 89.490 57.540 90.440 58.790 ;
        RECT 89.490 57.370 89.520 57.540 ;
        RECT 89.690 57.370 89.880 57.540 ;
        RECT 90.050 57.370 90.240 57.540 ;
        RECT 90.410 57.370 90.440 57.540 ;
        RECT 89.490 57.290 90.440 57.370 ;
      LAYER li1 ;
        RECT 90.620 57.290 90.950 58.970 ;
        RECT 91.730 58.930 92.060 59.270 ;
      LAYER li1 ;
        RECT 91.130 57.540 92.080 58.750 ;
        RECT 91.130 57.370 91.160 57.540 ;
        RECT 91.330 57.370 91.520 57.540 ;
        RECT 91.690 57.370 91.880 57.540 ;
        RECT 92.050 57.370 92.080 57.540 ;
        RECT 91.130 57.290 92.080 57.370 ;
        RECT 92.260 57.290 92.510 59.450 ;
        RECT 93.120 59.800 94.420 60.200 ;
        RECT 94.650 60.650 95.600 60.680 ;
        RECT 94.650 60.480 94.680 60.650 ;
        RECT 94.850 60.480 95.040 60.650 ;
        RECT 95.210 60.480 95.400 60.650 ;
        RECT 95.570 60.480 95.600 60.650 ;
        RECT 96.210 60.650 97.160 60.680 ;
        RECT 93.120 59.020 93.450 59.800 ;
        RECT 94.650 59.720 95.600 60.480 ;
      LAYER li1 ;
        RECT 95.780 59.840 96.030 60.550 ;
      LAYER li1 ;
        RECT 96.210 60.480 96.240 60.650 ;
        RECT 96.410 60.480 96.600 60.650 ;
        RECT 96.770 60.480 96.960 60.650 ;
        RECT 97.130 60.480 97.160 60.650 ;
        RECT 97.770 60.650 98.720 60.680 ;
        RECT 96.210 60.020 97.160 60.480 ;
      LAYER li1 ;
        RECT 97.340 59.840 97.590 60.550 ;
        RECT 95.780 59.670 97.590 59.840 ;
      LAYER li1 ;
        RECT 97.770 60.480 97.800 60.650 ;
        RECT 97.970 60.480 98.160 60.650 ;
        RECT 98.330 60.480 98.520 60.650 ;
        RECT 98.690 60.480 98.720 60.650 ;
        RECT 99.530 60.650 101.140 60.680 ;
        RECT 97.770 59.800 98.720 60.480 ;
      LAYER li1 ;
        RECT 95.780 59.500 95.950 59.670 ;
      LAYER li1 ;
        RECT 98.900 59.620 99.230 60.550 ;
        RECT 99.530 60.480 99.580 60.650 ;
        RECT 99.750 60.480 100.020 60.650 ;
        RECT 100.190 60.480 100.460 60.650 ;
        RECT 100.630 60.480 100.870 60.650 ;
        RECT 101.040 60.480 101.140 60.650 ;
        RECT 102.850 60.650 104.650 60.680 ;
        RECT 105.340 60.650 105.870 60.680 ;
        RECT 107.690 60.650 109.300 60.680 ;
        RECT 99.530 60.200 101.140 60.480 ;
        RECT 93.660 58.360 93.990 59.350 ;
      LAYER li1 ;
        RECT 94.690 59.270 95.950 59.500 ;
      LAYER li1 ;
        RECT 97.990 59.490 99.230 59.620 ;
        RECT 96.130 59.450 99.230 59.490 ;
        RECT 96.130 59.320 98.160 59.450 ;
      LAYER li1 ;
        RECT 95.780 59.140 95.950 59.270 ;
        RECT 95.780 58.970 97.670 59.140 ;
      LAYER li1 ;
        RECT 92.890 57.490 94.340 58.360 ;
        RECT 92.890 57.320 93.140 57.490 ;
        RECT 93.310 57.320 93.500 57.490 ;
        RECT 93.670 57.320 93.940 57.490 ;
        RECT 94.110 57.320 94.340 57.490 ;
        RECT 92.890 57.290 94.340 57.320 ;
        RECT 94.650 57.540 95.600 58.870 ;
        RECT 94.650 57.370 94.680 57.540 ;
        RECT 94.850 57.370 95.040 57.540 ;
        RECT 95.210 57.370 95.400 57.540 ;
        RECT 95.570 57.370 95.600 57.540 ;
        RECT 94.650 57.290 95.600 57.370 ;
      LAYER li1 ;
        RECT 95.780 57.290 96.030 58.970 ;
      LAYER li1 ;
        RECT 96.210 57.540 97.160 58.790 ;
        RECT 96.210 57.370 96.240 57.540 ;
        RECT 96.410 57.370 96.600 57.540 ;
        RECT 96.770 57.370 96.960 57.540 ;
        RECT 97.130 57.370 97.160 57.540 ;
        RECT 96.210 57.290 97.160 57.370 ;
      LAYER li1 ;
        RECT 97.340 57.290 97.670 58.970 ;
        RECT 98.450 58.930 98.780 59.270 ;
      LAYER li1 ;
        RECT 97.850 57.540 98.800 58.750 ;
        RECT 97.850 57.370 97.880 57.540 ;
        RECT 98.050 57.370 98.240 57.540 ;
        RECT 98.410 57.370 98.600 57.540 ;
        RECT 98.770 57.370 98.800 57.540 ;
        RECT 97.850 57.290 98.800 57.370 ;
        RECT 98.980 57.290 99.230 59.450 ;
        RECT 99.840 59.800 101.140 60.200 ;
        RECT 102.350 59.820 102.680 60.550 ;
        RECT 102.850 60.480 103.040 60.650 ;
        RECT 103.210 60.480 103.400 60.650 ;
        RECT 103.570 60.480 103.760 60.650 ;
        RECT 103.930 60.480 104.120 60.650 ;
        RECT 104.290 60.480 104.480 60.650 ;
        RECT 102.850 60.000 104.650 60.480 ;
        RECT 104.830 59.940 105.160 60.550 ;
        RECT 105.510 60.480 105.700 60.650 ;
        RECT 105.340 60.120 105.870 60.480 ;
        RECT 106.210 59.940 106.540 60.510 ;
        RECT 99.840 59.020 100.170 59.800 ;
        RECT 102.350 59.650 104.650 59.820 ;
        RECT 104.830 59.760 106.540 59.940 ;
        RECT 100.380 58.360 100.710 59.350 ;
        RECT 102.350 58.770 102.600 59.650 ;
        RECT 104.480 59.590 104.650 59.650 ;
      LAYER li1 ;
        RECT 102.820 59.120 103.150 59.320 ;
        RECT 103.330 59.300 104.300 59.470 ;
      LAYER li1 ;
        RECT 104.480 59.420 106.220 59.590 ;
      LAYER li1 ;
        RECT 106.990 59.500 107.400 60.510 ;
      LAYER li1 ;
        RECT 107.690 60.480 107.740 60.650 ;
        RECT 107.910 60.480 108.180 60.650 ;
        RECT 108.350 60.480 108.620 60.650 ;
        RECT 108.790 60.480 109.030 60.650 ;
        RECT 109.200 60.480 109.300 60.650 ;
        RECT 107.690 60.200 109.300 60.480 ;
        RECT 105.890 59.320 106.220 59.420 ;
      LAYER li1 ;
        RECT 105.170 59.120 105.500 59.240 ;
        RECT 106.690 59.140 107.400 59.500 ;
        RECT 102.820 58.950 105.500 59.120 ;
        RECT 103.810 58.930 105.500 58.950 ;
        RECT 106.270 58.970 107.400 59.140 ;
      LAYER li1 ;
        RECT 108.000 59.800 109.300 60.200 ;
        RECT 109.530 60.650 110.480 60.680 ;
        RECT 109.530 60.480 109.560 60.650 ;
        RECT 109.730 60.480 109.920 60.650 ;
        RECT 110.090 60.480 110.280 60.650 ;
        RECT 110.450 60.480 110.480 60.650 ;
        RECT 111.090 60.650 112.040 60.680 ;
        RECT 108.000 59.020 108.330 59.800 ;
        RECT 109.530 59.720 110.480 60.480 ;
      LAYER li1 ;
        RECT 110.660 59.840 110.910 60.550 ;
      LAYER li1 ;
        RECT 111.090 60.480 111.120 60.650 ;
        RECT 111.290 60.480 111.480 60.650 ;
        RECT 111.650 60.480 111.840 60.650 ;
        RECT 112.010 60.480 112.040 60.650 ;
        RECT 112.650 60.650 113.600 60.680 ;
        RECT 111.090 60.020 112.040 60.480 ;
      LAYER li1 ;
        RECT 112.220 59.840 112.470 60.550 ;
        RECT 110.660 59.670 112.470 59.840 ;
      LAYER li1 ;
        RECT 112.650 60.480 112.680 60.650 ;
        RECT 112.850 60.480 113.040 60.650 ;
        RECT 113.210 60.480 113.400 60.650 ;
        RECT 113.570 60.480 113.600 60.650 ;
        RECT 114.410 60.650 116.020 60.680 ;
        RECT 112.650 59.800 113.600 60.480 ;
      LAYER li1 ;
        RECT 110.660 59.500 110.830 59.670 ;
      LAYER li1 ;
        RECT 113.780 59.620 114.110 60.550 ;
        RECT 114.410 60.480 114.460 60.650 ;
        RECT 114.630 60.480 114.900 60.650 ;
        RECT 115.070 60.480 115.340 60.650 ;
        RECT 115.510 60.480 115.750 60.650 ;
        RECT 115.920 60.480 116.020 60.650 ;
        RECT 114.410 60.200 116.020 60.480 ;
        RECT 102.350 58.600 103.580 58.770 ;
        RECT 99.610 57.490 101.060 58.360 ;
        RECT 99.610 57.320 99.860 57.490 ;
        RECT 100.030 57.320 100.220 57.490 ;
        RECT 100.390 57.320 100.660 57.490 ;
        RECT 100.830 57.320 101.060 57.490 ;
        RECT 99.610 57.290 101.060 57.320 ;
        RECT 102.330 57.540 103.230 58.420 ;
        RECT 102.330 57.370 102.340 57.540 ;
        RECT 102.510 57.370 102.700 57.540 ;
        RECT 102.870 57.370 103.060 57.540 ;
        RECT 102.330 57.290 103.230 57.370 ;
        RECT 103.410 57.290 103.580 58.600 ;
        RECT 103.760 57.540 106.090 58.750 ;
        RECT 103.930 57.370 104.120 57.540 ;
        RECT 104.290 57.370 104.480 57.540 ;
        RECT 104.650 57.370 104.840 57.540 ;
        RECT 105.010 57.370 105.200 57.540 ;
        RECT 105.370 57.370 105.560 57.540 ;
        RECT 105.730 57.370 105.920 57.540 ;
        RECT 103.760 57.290 106.090 57.370 ;
      LAYER li1 ;
        RECT 106.270 57.290 106.520 58.970 ;
      LAYER li1 ;
        RECT 106.710 57.540 107.300 58.790 ;
        RECT 108.540 58.360 108.870 59.350 ;
      LAYER li1 ;
        RECT 109.570 59.270 110.830 59.500 ;
      LAYER li1 ;
        RECT 112.870 59.490 114.110 59.620 ;
        RECT 111.010 59.450 114.110 59.490 ;
        RECT 111.010 59.320 113.040 59.450 ;
      LAYER li1 ;
        RECT 110.660 59.140 110.830 59.270 ;
        RECT 110.660 58.970 112.550 59.140 ;
      LAYER li1 ;
        RECT 106.710 57.370 106.740 57.540 ;
        RECT 106.910 57.370 107.100 57.540 ;
        RECT 107.270 57.370 107.300 57.540 ;
        RECT 106.710 57.290 107.300 57.370 ;
        RECT 107.770 57.490 109.220 58.360 ;
        RECT 107.770 57.320 108.020 57.490 ;
        RECT 108.190 57.320 108.380 57.490 ;
        RECT 108.550 57.320 108.820 57.490 ;
        RECT 108.990 57.320 109.220 57.490 ;
        RECT 107.770 57.290 109.220 57.320 ;
        RECT 109.530 57.540 110.480 58.870 ;
        RECT 109.530 57.370 109.560 57.540 ;
        RECT 109.730 57.370 109.920 57.540 ;
        RECT 110.090 57.370 110.280 57.540 ;
        RECT 110.450 57.370 110.480 57.540 ;
        RECT 109.530 57.290 110.480 57.370 ;
      LAYER li1 ;
        RECT 110.660 57.290 110.910 58.970 ;
      LAYER li1 ;
        RECT 111.090 57.540 112.040 58.790 ;
        RECT 111.090 57.370 111.120 57.540 ;
        RECT 111.290 57.370 111.480 57.540 ;
        RECT 111.650 57.370 111.840 57.540 ;
        RECT 112.010 57.370 112.040 57.540 ;
        RECT 111.090 57.290 112.040 57.370 ;
      LAYER li1 ;
        RECT 112.220 57.290 112.550 58.970 ;
        RECT 113.330 58.930 113.660 59.270 ;
      LAYER li1 ;
        RECT 112.730 57.540 113.680 58.750 ;
        RECT 112.730 57.370 112.760 57.540 ;
        RECT 112.930 57.370 113.120 57.540 ;
        RECT 113.290 57.370 113.480 57.540 ;
        RECT 113.650 57.370 113.680 57.540 ;
        RECT 112.730 57.290 113.680 57.370 ;
        RECT 113.860 57.290 114.110 59.450 ;
        RECT 114.720 59.800 116.020 60.200 ;
        RECT 116.250 60.650 117.200 60.680 ;
        RECT 116.250 60.480 116.280 60.650 ;
        RECT 116.450 60.480 116.640 60.650 ;
        RECT 116.810 60.480 117.000 60.650 ;
        RECT 117.170 60.480 117.200 60.650 ;
        RECT 117.810 60.650 118.760 60.680 ;
        RECT 114.720 59.020 115.050 59.800 ;
        RECT 116.250 59.720 117.200 60.480 ;
      LAYER li1 ;
        RECT 117.380 59.840 117.630 60.550 ;
      LAYER li1 ;
        RECT 117.810 60.480 117.840 60.650 ;
        RECT 118.010 60.480 118.200 60.650 ;
        RECT 118.370 60.480 118.560 60.650 ;
        RECT 118.730 60.480 118.760 60.650 ;
        RECT 119.370 60.650 120.320 60.680 ;
        RECT 117.810 60.020 118.760 60.480 ;
      LAYER li1 ;
        RECT 118.940 59.840 119.190 60.550 ;
        RECT 117.380 59.670 119.190 59.840 ;
      LAYER li1 ;
        RECT 119.370 60.480 119.400 60.650 ;
        RECT 119.570 60.480 119.760 60.650 ;
        RECT 119.930 60.480 120.120 60.650 ;
        RECT 120.290 60.480 120.320 60.650 ;
        RECT 121.130 60.650 122.740 60.680 ;
        RECT 119.370 59.800 120.320 60.480 ;
      LAYER li1 ;
        RECT 117.380 59.500 117.550 59.670 ;
      LAYER li1 ;
        RECT 120.500 59.620 120.830 60.550 ;
        RECT 121.130 60.480 121.180 60.650 ;
        RECT 121.350 60.480 121.620 60.650 ;
        RECT 121.790 60.480 122.060 60.650 ;
        RECT 122.230 60.480 122.470 60.650 ;
        RECT 122.640 60.480 122.740 60.650 ;
        RECT 121.130 60.200 122.740 60.480 ;
        RECT 115.260 58.360 115.590 59.350 ;
      LAYER li1 ;
        RECT 116.290 59.270 117.550 59.500 ;
      LAYER li1 ;
        RECT 119.590 59.490 120.830 59.620 ;
        RECT 117.730 59.450 120.830 59.490 ;
        RECT 117.730 59.320 119.760 59.450 ;
      LAYER li1 ;
        RECT 117.380 59.140 117.550 59.270 ;
        RECT 117.380 58.970 119.270 59.140 ;
      LAYER li1 ;
        RECT 114.490 57.490 115.940 58.360 ;
        RECT 114.490 57.320 114.740 57.490 ;
        RECT 114.910 57.320 115.100 57.490 ;
        RECT 115.270 57.320 115.540 57.490 ;
        RECT 115.710 57.320 115.940 57.490 ;
        RECT 114.490 57.290 115.940 57.320 ;
        RECT 116.250 57.540 117.200 58.870 ;
        RECT 116.250 57.370 116.280 57.540 ;
        RECT 116.450 57.370 116.640 57.540 ;
        RECT 116.810 57.370 117.000 57.540 ;
        RECT 117.170 57.370 117.200 57.540 ;
        RECT 116.250 57.290 117.200 57.370 ;
      LAYER li1 ;
        RECT 117.380 57.290 117.630 58.970 ;
      LAYER li1 ;
        RECT 117.810 57.540 118.760 58.790 ;
        RECT 117.810 57.370 117.840 57.540 ;
        RECT 118.010 57.370 118.200 57.540 ;
        RECT 118.370 57.370 118.560 57.540 ;
        RECT 118.730 57.370 118.760 57.540 ;
        RECT 117.810 57.290 118.760 57.370 ;
      LAYER li1 ;
        RECT 118.940 57.290 119.270 58.970 ;
        RECT 120.050 58.930 120.380 59.270 ;
      LAYER li1 ;
        RECT 119.450 57.540 120.400 58.750 ;
        RECT 119.450 57.370 119.480 57.540 ;
        RECT 119.650 57.370 119.840 57.540 ;
        RECT 120.010 57.370 120.200 57.540 ;
        RECT 120.370 57.370 120.400 57.540 ;
        RECT 119.450 57.290 120.400 57.370 ;
        RECT 120.580 57.290 120.830 59.450 ;
        RECT 121.440 59.800 122.740 60.200 ;
        RECT 122.970 60.650 123.920 60.680 ;
        RECT 122.970 60.480 123.000 60.650 ;
        RECT 123.170 60.480 123.360 60.650 ;
        RECT 123.530 60.480 123.720 60.650 ;
        RECT 123.890 60.480 123.920 60.650 ;
        RECT 124.530 60.650 125.480 60.680 ;
        RECT 121.440 59.020 121.770 59.800 ;
        RECT 122.970 59.720 123.920 60.480 ;
      LAYER li1 ;
        RECT 124.100 59.840 124.350 60.550 ;
      LAYER li1 ;
        RECT 124.530 60.480 124.560 60.650 ;
        RECT 124.730 60.480 124.920 60.650 ;
        RECT 125.090 60.480 125.280 60.650 ;
        RECT 125.450 60.480 125.480 60.650 ;
        RECT 126.090 60.650 127.040 60.680 ;
        RECT 124.530 60.020 125.480 60.480 ;
      LAYER li1 ;
        RECT 125.660 59.840 125.910 60.550 ;
        RECT 124.100 59.670 125.910 59.840 ;
      LAYER li1 ;
        RECT 126.090 60.480 126.120 60.650 ;
        RECT 126.290 60.480 126.480 60.650 ;
        RECT 126.650 60.480 126.840 60.650 ;
        RECT 127.010 60.480 127.040 60.650 ;
        RECT 127.850 60.650 129.460 60.680 ;
        RECT 126.090 59.800 127.040 60.480 ;
      LAYER li1 ;
        RECT 124.100 59.500 124.270 59.670 ;
      LAYER li1 ;
        RECT 127.220 59.620 127.550 60.550 ;
        RECT 127.850 60.480 127.900 60.650 ;
        RECT 128.070 60.480 128.340 60.650 ;
        RECT 128.510 60.480 128.780 60.650 ;
        RECT 128.950 60.480 129.190 60.650 ;
        RECT 129.360 60.480 129.460 60.650 ;
        RECT 127.850 60.200 129.460 60.480 ;
        RECT 121.980 58.360 122.310 59.350 ;
      LAYER li1 ;
        RECT 123.010 59.270 124.270 59.500 ;
      LAYER li1 ;
        RECT 126.310 59.490 127.550 59.620 ;
        RECT 124.450 59.450 127.550 59.490 ;
        RECT 124.450 59.320 126.480 59.450 ;
      LAYER li1 ;
        RECT 124.100 59.140 124.270 59.270 ;
        RECT 124.100 58.970 125.990 59.140 ;
      LAYER li1 ;
        RECT 121.210 57.490 122.660 58.360 ;
        RECT 121.210 57.320 121.460 57.490 ;
        RECT 121.630 57.320 121.820 57.490 ;
        RECT 121.990 57.320 122.260 57.490 ;
        RECT 122.430 57.320 122.660 57.490 ;
        RECT 121.210 57.290 122.660 57.320 ;
        RECT 122.970 57.540 123.920 58.870 ;
        RECT 122.970 57.370 123.000 57.540 ;
        RECT 123.170 57.370 123.360 57.540 ;
        RECT 123.530 57.370 123.720 57.540 ;
        RECT 123.890 57.370 123.920 57.540 ;
        RECT 122.970 57.290 123.920 57.370 ;
      LAYER li1 ;
        RECT 124.100 57.290 124.350 58.970 ;
      LAYER li1 ;
        RECT 124.530 57.540 125.480 58.790 ;
        RECT 124.530 57.370 124.560 57.540 ;
        RECT 124.730 57.370 124.920 57.540 ;
        RECT 125.090 57.370 125.280 57.540 ;
        RECT 125.450 57.370 125.480 57.540 ;
        RECT 124.530 57.290 125.480 57.370 ;
      LAYER li1 ;
        RECT 125.660 57.290 125.990 58.970 ;
        RECT 126.770 58.930 127.100 59.270 ;
      LAYER li1 ;
        RECT 126.170 57.540 127.120 58.750 ;
        RECT 126.170 57.370 126.200 57.540 ;
        RECT 126.370 57.370 126.560 57.540 ;
        RECT 126.730 57.370 126.920 57.540 ;
        RECT 127.090 57.370 127.120 57.540 ;
        RECT 126.170 57.290 127.120 57.370 ;
        RECT 127.300 57.290 127.550 59.450 ;
        RECT 128.160 59.800 129.460 60.200 ;
        RECT 129.690 60.650 130.640 60.680 ;
        RECT 129.690 60.480 129.720 60.650 ;
        RECT 129.890 60.480 130.080 60.650 ;
        RECT 130.250 60.480 130.440 60.650 ;
        RECT 130.610 60.480 130.640 60.650 ;
        RECT 131.250 60.650 132.200 60.680 ;
        RECT 128.160 59.020 128.490 59.800 ;
        RECT 129.690 59.720 130.640 60.480 ;
      LAYER li1 ;
        RECT 130.820 59.840 131.070 60.550 ;
      LAYER li1 ;
        RECT 131.250 60.480 131.280 60.650 ;
        RECT 131.450 60.480 131.640 60.650 ;
        RECT 131.810 60.480 132.000 60.650 ;
        RECT 132.170 60.480 132.200 60.650 ;
        RECT 132.810 60.650 133.760 60.680 ;
        RECT 131.250 60.020 132.200 60.480 ;
      LAYER li1 ;
        RECT 132.380 59.840 132.630 60.550 ;
        RECT 130.820 59.670 132.630 59.840 ;
      LAYER li1 ;
        RECT 132.810 60.480 132.840 60.650 ;
        RECT 133.010 60.480 133.200 60.650 ;
        RECT 133.370 60.480 133.560 60.650 ;
        RECT 133.730 60.480 133.760 60.650 ;
        RECT 134.570 60.650 136.180 60.680 ;
        RECT 132.810 59.800 133.760 60.480 ;
      LAYER li1 ;
        RECT 130.820 59.500 130.990 59.670 ;
      LAYER li1 ;
        RECT 133.940 59.620 134.270 60.550 ;
        RECT 134.570 60.480 134.620 60.650 ;
        RECT 134.790 60.480 135.060 60.650 ;
        RECT 135.230 60.480 135.500 60.650 ;
        RECT 135.670 60.480 135.910 60.650 ;
        RECT 136.080 60.480 136.180 60.650 ;
        RECT 137.860 60.650 138.510 60.760 ;
        RECT 134.570 60.200 136.180 60.480 ;
        RECT 128.700 58.360 129.030 59.350 ;
      LAYER li1 ;
        RECT 129.730 59.270 130.990 59.500 ;
      LAYER li1 ;
        RECT 133.030 59.490 134.270 59.620 ;
        RECT 131.170 59.450 134.270 59.490 ;
        RECT 131.170 59.320 133.200 59.450 ;
      LAYER li1 ;
        RECT 130.820 59.140 130.990 59.270 ;
        RECT 130.820 58.970 132.710 59.140 ;
      LAYER li1 ;
        RECT 127.930 57.490 129.380 58.360 ;
        RECT 127.930 57.320 128.180 57.490 ;
        RECT 128.350 57.320 128.540 57.490 ;
        RECT 128.710 57.320 128.980 57.490 ;
        RECT 129.150 57.320 129.380 57.490 ;
        RECT 127.930 57.290 129.380 57.320 ;
        RECT 129.690 57.540 130.640 58.870 ;
        RECT 129.690 57.370 129.720 57.540 ;
        RECT 129.890 57.370 130.080 57.540 ;
        RECT 130.250 57.370 130.440 57.540 ;
        RECT 130.610 57.370 130.640 57.540 ;
        RECT 129.690 57.290 130.640 57.370 ;
      LAYER li1 ;
        RECT 130.820 57.290 131.070 58.970 ;
      LAYER li1 ;
        RECT 131.250 57.540 132.200 58.790 ;
        RECT 131.250 57.370 131.280 57.540 ;
        RECT 131.450 57.370 131.640 57.540 ;
        RECT 131.810 57.370 132.000 57.540 ;
        RECT 132.170 57.370 132.200 57.540 ;
        RECT 131.250 57.290 132.200 57.370 ;
      LAYER li1 ;
        RECT 132.380 57.290 132.710 58.970 ;
        RECT 133.490 58.930 133.820 59.270 ;
      LAYER li1 ;
        RECT 132.890 57.540 133.840 58.750 ;
        RECT 132.890 57.370 132.920 57.540 ;
        RECT 133.090 57.370 133.280 57.540 ;
        RECT 133.450 57.370 133.640 57.540 ;
        RECT 133.810 57.370 133.840 57.540 ;
        RECT 132.890 57.290 133.840 57.370 ;
        RECT 134.020 57.290 134.270 59.450 ;
        RECT 134.880 59.800 136.180 60.200 ;
      LAYER li1 ;
        RECT 136.610 59.980 137.190 60.620 ;
      LAYER li1 ;
        RECT 137.860 60.480 137.920 60.650 ;
        RECT 138.090 60.480 138.280 60.650 ;
        RECT 138.450 60.480 138.510 60.650 ;
        RECT 137.860 60.420 138.510 60.480 ;
        RECT 138.100 59.980 138.510 60.420 ;
        RECT 138.890 60.650 140.500 60.680 ;
        RECT 138.890 60.480 138.940 60.650 ;
        RECT 139.110 60.480 139.380 60.650 ;
        RECT 139.550 60.480 139.820 60.650 ;
        RECT 139.990 60.480 140.230 60.650 ;
        RECT 140.400 60.480 140.500 60.650 ;
        RECT 138.890 60.200 140.500 60.480 ;
        RECT 134.880 59.020 135.210 59.800 ;
        RECT 135.420 58.360 135.750 59.350 ;
      LAYER li1 ;
        RECT 136.940 59.110 137.190 59.980 ;
      LAYER li1 ;
        RECT 139.200 59.800 140.500 60.200 ;
      LAYER li1 ;
        RECT 136.940 58.860 137.650 59.110 ;
      LAYER li1 ;
        RECT 139.200 59.020 139.530 59.800 ;
        RECT 134.650 57.490 136.100 58.360 ;
        RECT 134.650 57.320 134.900 57.490 ;
        RECT 135.070 57.320 135.260 57.490 ;
        RECT 135.430 57.320 135.700 57.490 ;
        RECT 135.870 57.320 136.100 57.490 ;
        RECT 134.650 57.290 136.100 57.320 ;
        RECT 136.540 57.600 136.940 57.870 ;
        RECT 136.540 57.540 137.190 57.600 ;
        RECT 136.540 57.370 136.600 57.540 ;
        RECT 136.770 57.370 136.960 57.540 ;
        RECT 137.130 57.370 137.190 57.540 ;
      LAYER li1 ;
        RECT 137.400 57.520 137.650 58.860 ;
      LAYER li1 ;
        RECT 139.740 58.360 140.070 59.350 ;
        RECT 136.540 57.260 137.190 57.370 ;
        RECT 138.970 57.490 140.420 58.360 ;
        RECT 138.970 57.320 139.220 57.490 ;
        RECT 139.390 57.320 139.580 57.490 ;
        RECT 139.750 57.320 140.020 57.490 ;
        RECT 140.190 57.320 140.420 57.490 ;
        RECT 138.970 57.290 140.420 57.320 ;
        RECT 5.760 56.890 5.920 57.070 ;
        RECT 6.090 56.890 6.400 57.070 ;
        RECT 6.570 56.890 6.880 57.070 ;
        RECT 7.050 56.890 7.360 57.070 ;
        RECT 7.530 56.890 7.840 57.070 ;
        RECT 8.010 56.890 8.320 57.070 ;
        RECT 8.490 56.890 8.800 57.070 ;
        RECT 8.970 56.890 9.280 57.070 ;
        RECT 9.450 56.890 9.760 57.070 ;
        RECT 9.930 56.890 10.240 57.070 ;
        RECT 10.410 56.890 10.720 57.070 ;
        RECT 10.890 56.890 11.200 57.070 ;
        RECT 11.370 56.890 11.680 57.070 ;
        RECT 11.850 56.890 12.160 57.070 ;
        RECT 12.330 56.890 12.640 57.070 ;
        RECT 12.810 56.890 13.120 57.070 ;
        RECT 13.290 56.890 13.600 57.070 ;
        RECT 13.770 56.890 14.080 57.070 ;
        RECT 14.250 56.890 14.560 57.070 ;
        RECT 14.730 56.890 15.040 57.070 ;
        RECT 15.210 56.890 15.520 57.070 ;
        RECT 15.690 56.890 16.000 57.070 ;
        RECT 16.170 56.890 16.480 57.070 ;
        RECT 16.650 56.890 16.960 57.070 ;
        RECT 17.130 56.890 17.440 57.070 ;
        RECT 17.610 56.890 17.920 57.070 ;
        RECT 18.090 56.890 18.400 57.070 ;
        RECT 18.570 56.890 18.880 57.070 ;
        RECT 19.050 56.890 19.360 57.070 ;
        RECT 19.530 56.890 19.840 57.070 ;
        RECT 20.010 56.890 20.320 57.070 ;
        RECT 20.490 56.890 20.800 57.070 ;
        RECT 20.970 56.890 21.280 57.070 ;
        RECT 21.450 56.890 21.760 57.070 ;
        RECT 21.930 56.890 22.240 57.070 ;
        RECT 22.410 56.890 22.720 57.070 ;
        RECT 22.890 56.890 23.200 57.070 ;
        RECT 23.370 56.890 23.680 57.070 ;
        RECT 23.850 56.890 24.160 57.070 ;
        RECT 24.330 56.890 24.640 57.070 ;
        RECT 24.810 56.890 25.120 57.070 ;
        RECT 25.290 56.890 25.600 57.070 ;
        RECT 25.770 56.890 26.080 57.070 ;
        RECT 26.250 56.890 26.560 57.070 ;
        RECT 26.730 56.890 27.040 57.070 ;
        RECT 27.210 56.890 27.520 57.070 ;
        RECT 27.690 56.890 28.000 57.070 ;
        RECT 28.170 56.890 28.480 57.070 ;
        RECT 28.650 56.890 28.960 57.070 ;
        RECT 29.130 56.890 29.440 57.070 ;
        RECT 29.610 56.890 29.920 57.070 ;
        RECT 30.090 56.890 30.400 57.070 ;
        RECT 30.570 56.890 30.880 57.070 ;
        RECT 31.050 56.890 31.360 57.070 ;
        RECT 31.530 56.890 31.840 57.070 ;
        RECT 32.010 56.890 32.320 57.070 ;
        RECT 32.490 56.890 32.800 57.070 ;
        RECT 32.970 56.890 33.280 57.070 ;
        RECT 33.450 56.890 33.760 57.070 ;
        RECT 33.930 56.890 34.240 57.070 ;
        RECT 34.410 56.890 34.720 57.070 ;
        RECT 34.890 56.890 35.200 57.070 ;
        RECT 35.370 56.890 35.680 57.070 ;
        RECT 35.850 56.890 36.160 57.070 ;
        RECT 36.330 56.890 36.640 57.070 ;
        RECT 36.810 56.890 37.120 57.070 ;
        RECT 37.290 56.890 37.600 57.070 ;
        RECT 37.770 56.890 38.080 57.070 ;
        RECT 38.250 56.890 38.560 57.070 ;
        RECT 38.730 56.890 39.040 57.070 ;
        RECT 39.210 56.890 39.520 57.070 ;
        RECT 39.690 56.890 40.000 57.070 ;
        RECT 40.170 56.890 40.480 57.070 ;
        RECT 40.650 56.890 40.960 57.070 ;
        RECT 41.130 56.890 41.440 57.070 ;
        RECT 41.610 56.890 41.920 57.070 ;
        RECT 42.090 56.890 42.400 57.070 ;
        RECT 42.570 56.890 42.880 57.070 ;
        RECT 43.050 56.890 43.360 57.070 ;
        RECT 43.530 56.890 43.840 57.070 ;
        RECT 44.010 56.890 44.320 57.070 ;
        RECT 44.490 56.890 44.800 57.070 ;
        RECT 44.970 56.890 45.280 57.070 ;
        RECT 45.450 56.890 45.760 57.070 ;
        RECT 45.930 56.890 46.240 57.070 ;
        RECT 46.410 56.890 46.720 57.070 ;
        RECT 46.890 56.890 47.200 57.070 ;
        RECT 47.370 56.890 47.680 57.070 ;
        RECT 47.850 56.890 48.160 57.070 ;
        RECT 48.330 56.890 48.640 57.070 ;
        RECT 48.810 56.890 49.120 57.070 ;
        RECT 49.290 57.060 49.600 57.070 ;
        RECT 49.770 57.060 50.080 57.070 ;
        RECT 49.290 56.890 49.440 57.060 ;
        RECT 49.920 56.890 50.080 57.060 ;
        RECT 50.250 56.890 50.560 57.070 ;
        RECT 50.730 56.890 51.040 57.070 ;
        RECT 51.210 56.890 51.520 57.070 ;
        RECT 51.690 56.890 52.000 57.070 ;
        RECT 52.170 56.890 52.480 57.070 ;
        RECT 52.650 56.890 52.960 57.070 ;
        RECT 53.130 56.890 53.440 57.070 ;
        RECT 53.610 56.890 53.920 57.070 ;
        RECT 54.090 56.890 54.400 57.070 ;
        RECT 54.570 56.890 54.880 57.070 ;
        RECT 55.050 56.890 55.360 57.070 ;
        RECT 55.530 56.890 55.840 57.070 ;
        RECT 56.010 56.890 56.320 57.070 ;
        RECT 56.490 56.890 56.800 57.070 ;
        RECT 56.970 56.890 57.280 57.070 ;
        RECT 57.450 56.890 57.760 57.070 ;
        RECT 57.930 56.890 58.240 57.070 ;
        RECT 58.410 56.890 58.720 57.070 ;
        RECT 58.890 56.890 59.200 57.070 ;
        RECT 59.370 56.890 59.680 57.070 ;
        RECT 59.850 56.890 60.160 57.070 ;
        RECT 60.330 56.890 60.640 57.070 ;
        RECT 60.810 56.890 61.120 57.070 ;
        RECT 61.290 56.890 61.600 57.070 ;
        RECT 61.770 56.890 62.080 57.070 ;
        RECT 62.250 56.890 62.560 57.070 ;
        RECT 62.730 56.890 63.040 57.070 ;
        RECT 63.210 56.890 63.520 57.070 ;
        RECT 63.690 56.890 64.000 57.070 ;
        RECT 64.170 56.890 64.480 57.070 ;
        RECT 64.650 56.890 64.960 57.070 ;
        RECT 65.130 56.890 65.440 57.070 ;
        RECT 65.610 56.890 65.920 57.070 ;
        RECT 66.090 56.890 66.400 57.070 ;
        RECT 66.570 56.890 66.880 57.070 ;
        RECT 67.050 56.890 67.360 57.070 ;
        RECT 67.530 56.890 67.840 57.070 ;
        RECT 68.010 56.890 68.320 57.070 ;
        RECT 68.490 56.890 68.800 57.070 ;
        RECT 68.970 56.890 69.280 57.070 ;
        RECT 69.450 56.890 69.760 57.070 ;
        RECT 69.930 56.890 70.240 57.070 ;
        RECT 70.410 56.890 70.720 57.070 ;
        RECT 70.890 56.890 71.200 57.070 ;
        RECT 71.370 56.890 71.680 57.070 ;
        RECT 71.850 56.890 72.160 57.070 ;
        RECT 72.330 56.890 72.640 57.070 ;
        RECT 72.810 56.890 73.120 57.070 ;
        RECT 73.290 56.890 73.600 57.070 ;
        RECT 73.770 56.890 74.080 57.070 ;
        RECT 74.250 56.890 74.560 57.070 ;
        RECT 74.730 56.890 75.040 57.070 ;
        RECT 75.210 56.890 75.520 57.070 ;
        RECT 75.690 56.890 76.000 57.070 ;
        RECT 76.170 56.890 76.480 57.070 ;
        RECT 76.650 56.890 76.960 57.070 ;
        RECT 77.130 56.890 77.440 57.070 ;
        RECT 77.610 56.890 77.920 57.070 ;
        RECT 78.090 56.890 78.400 57.070 ;
        RECT 78.570 56.890 78.880 57.070 ;
        RECT 79.050 56.890 79.360 57.070 ;
        RECT 79.530 56.890 79.840 57.070 ;
        RECT 80.010 56.890 80.320 57.070 ;
        RECT 80.490 56.890 80.800 57.070 ;
        RECT 80.970 56.890 81.280 57.070 ;
        RECT 81.450 56.890 81.760 57.070 ;
        RECT 81.930 56.890 82.240 57.070 ;
        RECT 82.410 56.890 82.720 57.070 ;
        RECT 82.890 56.890 83.200 57.070 ;
        RECT 83.370 56.890 83.680 57.070 ;
        RECT 83.850 56.890 84.160 57.070 ;
        RECT 84.330 56.890 84.640 57.070 ;
        RECT 84.810 56.890 85.120 57.070 ;
        RECT 85.290 56.890 85.600 57.070 ;
        RECT 85.770 56.890 86.080 57.070 ;
        RECT 86.250 56.890 86.560 57.070 ;
        RECT 86.730 56.890 87.040 57.070 ;
        RECT 87.210 56.890 87.520 57.070 ;
        RECT 87.690 56.890 88.000 57.070 ;
        RECT 88.170 56.890 88.480 57.070 ;
        RECT 88.650 56.890 88.960 57.070 ;
        RECT 89.130 56.890 89.440 57.070 ;
        RECT 89.610 56.890 89.920 57.070 ;
        RECT 90.090 56.890 90.400 57.070 ;
        RECT 90.570 56.890 90.880 57.070 ;
        RECT 91.050 56.890 91.360 57.070 ;
        RECT 91.530 56.890 91.840 57.070 ;
        RECT 92.010 56.890 92.320 57.070 ;
        RECT 92.490 56.890 92.800 57.070 ;
        RECT 92.970 56.890 93.280 57.070 ;
        RECT 93.450 56.890 93.760 57.070 ;
        RECT 93.930 56.890 94.240 57.070 ;
        RECT 94.410 56.890 94.720 57.070 ;
        RECT 94.890 56.890 95.200 57.070 ;
        RECT 95.370 56.890 95.680 57.070 ;
        RECT 95.850 56.890 96.160 57.070 ;
        RECT 96.330 56.890 96.640 57.070 ;
        RECT 96.810 56.890 97.120 57.070 ;
        RECT 97.290 56.890 97.600 57.070 ;
        RECT 97.770 56.890 98.080 57.070 ;
        RECT 98.250 56.890 98.560 57.070 ;
        RECT 98.730 56.890 99.040 57.070 ;
        RECT 99.210 56.890 99.520 57.070 ;
        RECT 99.690 56.890 100.000 57.070 ;
        RECT 100.170 56.890 100.480 57.070 ;
        RECT 100.650 56.890 100.960 57.070 ;
        RECT 101.130 56.890 101.440 57.070 ;
        RECT 101.610 57.060 101.760 57.070 ;
        RECT 102.240 57.060 102.400 57.070 ;
        RECT 101.610 56.890 101.920 57.060 ;
        RECT 102.090 56.890 102.400 57.060 ;
        RECT 102.570 56.890 102.880 57.070 ;
        RECT 103.050 56.890 103.360 57.070 ;
        RECT 103.530 56.890 103.840 57.070 ;
        RECT 104.010 56.890 104.320 57.070 ;
        RECT 104.490 56.890 104.800 57.070 ;
        RECT 104.970 56.890 105.280 57.070 ;
        RECT 105.450 56.890 105.760 57.070 ;
        RECT 105.930 56.890 106.240 57.070 ;
        RECT 106.410 56.890 106.720 57.070 ;
        RECT 106.890 56.890 107.200 57.070 ;
        RECT 107.370 56.890 107.680 57.070 ;
        RECT 107.850 56.890 108.160 57.070 ;
        RECT 108.330 56.890 108.640 57.070 ;
        RECT 108.810 56.890 109.120 57.070 ;
        RECT 109.290 56.890 109.600 57.070 ;
        RECT 109.770 56.890 110.080 57.070 ;
        RECT 110.250 56.890 110.560 57.070 ;
        RECT 110.730 56.890 111.040 57.070 ;
        RECT 111.210 56.890 111.520 57.070 ;
        RECT 111.690 56.890 112.000 57.070 ;
        RECT 112.170 56.890 112.480 57.070 ;
        RECT 112.650 56.890 112.960 57.070 ;
        RECT 113.130 56.890 113.440 57.070 ;
        RECT 113.610 56.890 113.920 57.070 ;
        RECT 114.090 56.890 114.400 57.070 ;
        RECT 114.570 56.890 114.880 57.070 ;
        RECT 115.050 56.890 115.360 57.070 ;
        RECT 115.530 57.060 115.680 57.070 ;
        RECT 116.160 57.060 116.320 57.070 ;
        RECT 115.530 56.890 115.840 57.060 ;
        RECT 116.010 56.890 116.320 57.060 ;
        RECT 116.490 56.890 116.800 57.070 ;
        RECT 116.970 56.890 117.280 57.070 ;
        RECT 117.450 56.890 117.760 57.070 ;
        RECT 117.930 56.890 118.240 57.070 ;
        RECT 118.410 56.890 118.720 57.070 ;
        RECT 118.890 56.890 119.200 57.070 ;
        RECT 119.370 56.890 119.680 57.070 ;
        RECT 119.850 56.890 120.160 57.070 ;
        RECT 120.330 56.890 120.640 57.070 ;
        RECT 120.810 56.890 121.120 57.070 ;
        RECT 121.290 56.890 121.600 57.070 ;
        RECT 121.770 56.890 122.080 57.070 ;
        RECT 122.250 56.890 122.560 57.070 ;
        RECT 122.730 56.890 123.040 57.070 ;
        RECT 123.210 56.890 123.520 57.070 ;
        RECT 123.690 56.890 124.000 57.070 ;
        RECT 124.170 56.890 124.480 57.070 ;
        RECT 124.650 56.890 124.960 57.070 ;
        RECT 125.130 56.890 125.440 57.070 ;
        RECT 125.610 56.890 125.920 57.070 ;
        RECT 126.090 56.890 126.400 57.070 ;
        RECT 126.570 56.890 126.880 57.070 ;
        RECT 127.050 56.890 127.360 57.070 ;
        RECT 127.530 56.890 127.840 57.070 ;
        RECT 128.010 56.890 128.320 57.070 ;
        RECT 128.490 56.890 128.800 57.070 ;
        RECT 128.970 56.890 129.280 57.070 ;
        RECT 129.450 56.890 129.760 57.070 ;
        RECT 129.930 56.890 130.240 57.070 ;
        RECT 130.410 56.890 130.720 57.070 ;
        RECT 130.890 56.890 131.200 57.070 ;
        RECT 131.370 56.890 131.680 57.070 ;
        RECT 131.850 56.890 132.160 57.070 ;
        RECT 132.330 56.890 132.640 57.070 ;
        RECT 132.810 56.890 133.120 57.070 ;
        RECT 133.290 56.890 133.600 57.070 ;
        RECT 133.770 56.890 134.080 57.070 ;
        RECT 134.250 56.890 134.560 57.070 ;
        RECT 134.730 56.890 135.040 57.070 ;
        RECT 135.210 56.890 135.520 57.070 ;
        RECT 135.690 56.890 136.000 57.070 ;
        RECT 136.170 56.890 136.480 57.070 ;
        RECT 136.650 56.890 136.960 57.070 ;
        RECT 137.130 56.890 137.440 57.070 ;
        RECT 137.610 56.890 137.920 57.070 ;
        RECT 138.090 56.890 138.400 57.070 ;
        RECT 138.570 56.890 138.880 57.070 ;
        RECT 139.050 56.890 139.360 57.070 ;
        RECT 139.530 56.890 139.840 57.070 ;
        RECT 140.010 56.890 140.320 57.070 ;
        RECT 140.490 56.890 140.800 57.070 ;
        RECT 140.970 56.890 141.280 57.070 ;
        RECT 141.450 57.060 141.760 57.070 ;
        RECT 141.930 57.060 142.080 57.070 ;
        RECT 141.450 56.890 141.600 57.060 ;
        RECT 5.850 56.590 6.440 56.670 ;
        RECT 5.850 56.420 5.880 56.590 ;
        RECT 6.050 56.420 6.240 56.590 ;
        RECT 6.410 56.420 6.440 56.590 ;
        RECT 5.850 55.090 6.440 56.420 ;
      LAYER li1 ;
        RECT 6.720 55.090 7.110 56.670 ;
      LAYER li1 ;
        RECT 7.450 56.640 8.900 56.670 ;
        RECT 7.450 56.470 7.700 56.640 ;
        RECT 7.870 56.470 8.060 56.640 ;
        RECT 8.230 56.470 8.500 56.640 ;
        RECT 8.670 56.470 8.900 56.640 ;
        RECT 7.450 55.600 8.900 56.470 ;
        RECT 9.210 56.590 9.800 56.670 ;
        RECT 9.210 56.420 9.240 56.590 ;
        RECT 9.410 56.420 9.600 56.590 ;
        RECT 9.770 56.420 9.800 56.590 ;
      LAYER li1 ;
        RECT 5.890 54.460 6.600 54.850 ;
      LAYER li1 ;
        RECT 5.850 53.280 6.440 54.240 ;
      LAYER li1 ;
        RECT 6.780 53.410 7.110 55.090 ;
      LAYER li1 ;
        RECT 7.680 54.160 8.010 54.940 ;
        RECT 8.220 54.610 8.550 55.600 ;
        RECT 9.210 55.090 9.800 56.420 ;
      LAYER li1 ;
        RECT 10.080 55.090 10.470 56.670 ;
      LAYER li1 ;
        RECT 10.810 56.640 12.260 56.670 ;
        RECT 10.810 56.470 11.060 56.640 ;
        RECT 11.230 56.470 11.420 56.640 ;
        RECT 11.590 56.470 11.860 56.640 ;
        RECT 12.030 56.470 12.260 56.640 ;
        RECT 10.810 55.600 12.260 56.470 ;
      LAYER li1 ;
        RECT 9.250 54.460 9.960 54.850 ;
      LAYER li1 ;
        RECT 7.680 53.760 8.980 54.160 ;
        RECT 7.370 53.280 8.980 53.760 ;
        RECT 9.210 53.280 9.800 54.240 ;
      LAYER li1 ;
        RECT 10.140 53.410 10.470 55.090 ;
      LAYER li1 ;
        RECT 11.040 54.160 11.370 54.940 ;
        RECT 11.580 54.610 11.910 55.600 ;
      LAYER li1 ;
        RECT 12.600 55.090 13.030 56.670 ;
      LAYER li1 ;
        RECT 13.210 56.590 13.770 56.670 ;
        RECT 13.210 56.420 13.220 56.590 ;
        RECT 13.390 56.420 13.580 56.590 ;
        RECT 13.750 56.420 13.770 56.590 ;
        RECT 13.210 55.090 13.770 56.420 ;
        RECT 15.130 56.640 16.580 56.670 ;
        RECT 15.130 56.470 15.380 56.640 ;
        RECT 15.550 56.470 15.740 56.640 ;
        RECT 15.910 56.470 16.180 56.640 ;
        RECT 16.350 56.470 16.580 56.640 ;
        RECT 11.040 53.760 12.340 54.160 ;
        RECT 10.730 53.280 12.340 53.760 ;
      LAYER li1 ;
        RECT 12.600 53.410 12.850 55.090 ;
      LAYER li1 ;
        RECT 13.160 54.200 13.490 54.660 ;
      LAYER li1 ;
        RECT 13.950 54.380 14.280 56.170 ;
      LAYER li1 ;
        RECT 14.460 54.200 14.710 55.920 ;
        RECT 15.130 55.600 16.580 56.470 ;
        RECT 16.890 56.590 18.560 56.670 ;
        RECT 16.890 56.420 16.920 56.590 ;
        RECT 17.090 56.420 17.280 56.590 ;
        RECT 17.450 56.420 17.640 56.590 ;
        RECT 17.810 56.420 18.000 56.590 ;
        RECT 18.170 56.420 18.360 56.590 ;
        RECT 18.530 56.420 18.560 56.590 ;
        RECT 13.160 54.030 14.710 54.200 ;
        RECT 13.030 53.280 14.280 53.850 ;
        RECT 14.460 53.410 14.710 54.030 ;
        RECT 15.360 54.160 15.690 54.940 ;
        RECT 15.900 54.610 16.230 55.600 ;
        RECT 16.890 55.210 18.560 56.420 ;
      LAYER li1 ;
        RECT 16.930 54.440 17.230 55.030 ;
        RECT 17.410 54.690 18.600 55.030 ;
        RECT 18.780 54.690 19.110 56.170 ;
        RECT 19.290 54.510 19.560 56.670 ;
      LAYER li1 ;
        RECT 20.410 56.640 21.860 56.670 ;
        RECT 20.410 56.470 20.660 56.640 ;
        RECT 20.830 56.470 21.020 56.640 ;
        RECT 21.190 56.470 21.460 56.640 ;
        RECT 21.630 56.470 21.860 56.640 ;
        RECT 20.410 55.600 21.860 56.470 ;
        RECT 22.170 56.590 23.430 56.670 ;
        RECT 22.170 56.420 22.180 56.590 ;
        RECT 22.350 56.420 22.540 56.590 ;
        RECT 22.710 56.420 22.900 56.590 ;
        RECT 23.070 56.420 23.260 56.590 ;
      LAYER li1 ;
        RECT 17.730 54.340 19.560 54.510 ;
      LAYER li1 ;
        RECT 15.360 53.760 16.660 54.160 ;
        RECT 15.050 53.280 16.660 53.760 ;
        RECT 16.890 53.280 17.480 54.240 ;
      LAYER li1 ;
        RECT 17.730 53.410 17.980 54.340 ;
      LAYER li1 ;
        RECT 18.160 53.280 19.110 54.160 ;
      LAYER li1 ;
        RECT 19.290 53.410 19.560 54.340 ;
        RECT 19.830 53.750 20.000 55.030 ;
      LAYER li1 ;
        RECT 20.640 54.160 20.970 54.940 ;
        RECT 21.180 54.610 21.510 55.600 ;
        RECT 22.170 55.190 23.430 56.420 ;
      LAYER li1 ;
        RECT 23.960 56.170 24.130 56.670 ;
        RECT 23.610 55.090 24.130 56.170 ;
      LAYER li1 ;
        RECT 24.390 56.590 25.700 56.670 ;
        RECT 24.390 56.420 24.420 56.590 ;
        RECT 24.590 56.420 24.780 56.590 ;
        RECT 24.950 56.420 25.140 56.590 ;
        RECT 25.310 56.420 25.500 56.590 ;
        RECT 25.670 56.420 25.700 56.590 ;
        RECT 24.390 55.210 25.700 56.420 ;
        RECT 26.170 56.640 27.620 56.670 ;
        RECT 26.170 56.470 26.420 56.640 ;
        RECT 26.590 56.470 26.780 56.640 ;
        RECT 26.950 56.470 27.220 56.640 ;
        RECT 27.390 56.470 27.620 56.640 ;
        RECT 26.170 55.600 27.620 56.470 ;
        RECT 27.930 56.590 28.880 56.670 ;
        RECT 27.930 56.420 27.960 56.590 ;
        RECT 28.130 56.420 28.320 56.590 ;
        RECT 28.490 56.420 28.680 56.590 ;
        RECT 28.850 56.420 28.880 56.590 ;
      LAYER li1 ;
        RECT 23.610 55.010 23.880 55.090 ;
        RECT 22.820 54.840 23.880 55.010 ;
        RECT 22.210 54.450 22.630 54.780 ;
        RECT 22.820 54.270 22.990 54.840 ;
        RECT 24.330 54.720 24.840 55.030 ;
        RECT 25.090 54.720 25.800 55.030 ;
        RECT 23.170 54.450 23.680 54.660 ;
      LAYER li1 ;
        RECT 23.880 54.370 25.750 54.540 ;
        RECT 20.640 53.760 21.940 54.160 ;
        RECT 20.330 53.280 21.940 53.760 ;
        RECT 22.240 53.350 22.570 54.270 ;
      LAYER li1 ;
        RECT 22.820 53.530 23.350 54.270 ;
      LAYER li1 ;
        RECT 23.880 53.350 24.050 54.370 ;
        RECT 22.240 53.180 24.050 53.350 ;
        RECT 24.230 53.280 25.330 54.190 ;
        RECT 25.500 53.440 25.750 54.370 ;
        RECT 26.400 54.160 26.730 54.940 ;
        RECT 26.940 54.610 27.270 55.600 ;
        RECT 27.930 55.090 28.880 56.420 ;
      LAYER li1 ;
        RECT 29.060 54.990 29.310 56.670 ;
      LAYER li1 ;
        RECT 29.490 56.590 30.440 56.670 ;
        RECT 29.490 56.420 29.520 56.590 ;
        RECT 29.690 56.420 29.880 56.590 ;
        RECT 30.050 56.420 30.240 56.590 ;
        RECT 30.410 56.420 30.440 56.590 ;
        RECT 29.490 55.170 30.440 56.420 ;
      LAYER li1 ;
        RECT 30.620 54.990 30.950 56.670 ;
      LAYER li1 ;
        RECT 31.130 56.590 32.080 56.670 ;
        RECT 31.130 56.420 31.160 56.590 ;
        RECT 31.330 56.420 31.520 56.590 ;
        RECT 31.690 56.420 31.880 56.590 ;
        RECT 32.050 56.420 32.080 56.590 ;
        RECT 31.130 55.210 32.080 56.420 ;
      LAYER li1 ;
        RECT 29.060 54.820 30.950 54.990 ;
        RECT 29.060 54.690 29.230 54.820 ;
        RECT 31.730 54.690 32.060 55.030 ;
        RECT 27.970 54.460 29.230 54.690 ;
      LAYER li1 ;
        RECT 29.410 54.510 31.440 54.640 ;
        RECT 32.260 54.510 32.510 56.670 ;
        RECT 32.890 56.640 34.340 56.670 ;
        RECT 32.890 56.470 33.140 56.640 ;
        RECT 33.310 56.470 33.500 56.640 ;
        RECT 33.670 56.470 33.940 56.640 ;
        RECT 34.110 56.470 34.340 56.640 ;
        RECT 32.890 55.600 34.340 56.470 ;
        RECT 34.650 56.590 35.600 56.670 ;
        RECT 34.650 56.420 34.680 56.590 ;
        RECT 34.850 56.420 35.040 56.590 ;
        RECT 35.210 56.420 35.400 56.590 ;
        RECT 35.570 56.420 35.600 56.590 ;
        RECT 29.410 54.470 32.510 54.510 ;
      LAYER li1 ;
        RECT 29.060 54.290 29.230 54.460 ;
      LAYER li1 ;
        RECT 31.270 54.340 32.510 54.470 ;
        RECT 26.400 53.760 27.700 54.160 ;
        RECT 26.090 53.280 27.700 53.760 ;
        RECT 27.930 53.280 28.880 54.240 ;
      LAYER li1 ;
        RECT 29.060 54.120 30.870 54.290 ;
        RECT 29.060 53.410 29.310 54.120 ;
      LAYER li1 ;
        RECT 29.490 53.280 30.440 53.940 ;
      LAYER li1 ;
        RECT 30.620 53.410 30.870 54.120 ;
      LAYER li1 ;
        RECT 31.050 53.280 32.000 54.160 ;
        RECT 32.180 53.410 32.510 54.340 ;
        RECT 33.120 54.160 33.450 54.940 ;
        RECT 33.660 54.610 33.990 55.600 ;
        RECT 34.650 55.090 35.600 56.420 ;
      LAYER li1 ;
        RECT 35.780 54.990 36.030 56.670 ;
      LAYER li1 ;
        RECT 36.210 56.590 37.160 56.670 ;
        RECT 36.210 56.420 36.240 56.590 ;
        RECT 36.410 56.420 36.600 56.590 ;
        RECT 36.770 56.420 36.960 56.590 ;
        RECT 37.130 56.420 37.160 56.590 ;
        RECT 36.210 55.170 37.160 56.420 ;
      LAYER li1 ;
        RECT 37.340 54.990 37.670 56.670 ;
      LAYER li1 ;
        RECT 37.850 56.590 38.800 56.670 ;
        RECT 37.850 56.420 37.880 56.590 ;
        RECT 38.050 56.420 38.240 56.590 ;
        RECT 38.410 56.420 38.600 56.590 ;
        RECT 38.770 56.420 38.800 56.590 ;
        RECT 37.850 55.210 38.800 56.420 ;
      LAYER li1 ;
        RECT 35.780 54.820 37.670 54.990 ;
        RECT 35.780 54.690 35.950 54.820 ;
        RECT 38.450 54.690 38.780 55.030 ;
        RECT 34.690 54.460 35.950 54.690 ;
      LAYER li1 ;
        RECT 36.130 54.510 38.160 54.640 ;
        RECT 38.980 54.510 39.230 56.670 ;
        RECT 39.610 56.640 41.060 56.670 ;
        RECT 39.610 56.470 39.860 56.640 ;
        RECT 40.030 56.470 40.220 56.640 ;
        RECT 40.390 56.470 40.660 56.640 ;
        RECT 40.830 56.470 41.060 56.640 ;
        RECT 39.610 55.600 41.060 56.470 ;
        RECT 41.370 56.590 42.320 56.670 ;
        RECT 41.370 56.420 41.400 56.590 ;
        RECT 41.570 56.420 41.760 56.590 ;
        RECT 41.930 56.420 42.120 56.590 ;
        RECT 42.290 56.420 42.320 56.590 ;
        RECT 36.130 54.470 39.230 54.510 ;
      LAYER li1 ;
        RECT 35.780 54.290 35.950 54.460 ;
      LAYER li1 ;
        RECT 37.990 54.340 39.230 54.470 ;
        RECT 33.120 53.760 34.420 54.160 ;
        RECT 32.810 53.280 34.420 53.760 ;
        RECT 34.650 53.280 35.600 54.240 ;
      LAYER li1 ;
        RECT 35.780 54.120 37.590 54.290 ;
        RECT 35.780 53.410 36.030 54.120 ;
      LAYER li1 ;
        RECT 36.210 53.280 37.160 53.940 ;
      LAYER li1 ;
        RECT 37.340 53.410 37.590 54.120 ;
      LAYER li1 ;
        RECT 37.770 53.280 38.720 54.160 ;
        RECT 38.900 53.410 39.230 54.340 ;
        RECT 39.840 54.160 40.170 54.940 ;
        RECT 40.380 54.610 40.710 55.600 ;
        RECT 41.370 55.090 42.320 56.420 ;
      LAYER li1 ;
        RECT 42.500 54.990 42.750 56.670 ;
      LAYER li1 ;
        RECT 42.930 56.590 43.880 56.670 ;
        RECT 42.930 56.420 42.960 56.590 ;
        RECT 43.130 56.420 43.320 56.590 ;
        RECT 43.490 56.420 43.680 56.590 ;
        RECT 43.850 56.420 43.880 56.590 ;
        RECT 42.930 55.170 43.880 56.420 ;
      LAYER li1 ;
        RECT 44.060 54.990 44.390 56.670 ;
      LAYER li1 ;
        RECT 44.570 56.590 45.520 56.670 ;
        RECT 44.570 56.420 44.600 56.590 ;
        RECT 44.770 56.420 44.960 56.590 ;
        RECT 45.130 56.420 45.320 56.590 ;
        RECT 45.490 56.420 45.520 56.590 ;
        RECT 44.570 55.210 45.520 56.420 ;
      LAYER li1 ;
        RECT 42.500 54.820 44.390 54.990 ;
        RECT 42.500 54.690 42.670 54.820 ;
        RECT 45.170 54.690 45.500 55.030 ;
        RECT 41.410 54.460 42.670 54.690 ;
      LAYER li1 ;
        RECT 42.850 54.510 44.880 54.640 ;
        RECT 45.700 54.510 45.950 56.670 ;
        RECT 46.330 56.640 47.780 56.670 ;
        RECT 46.330 56.470 46.580 56.640 ;
        RECT 46.750 56.470 46.940 56.640 ;
        RECT 47.110 56.470 47.380 56.640 ;
        RECT 47.550 56.470 47.780 56.640 ;
        RECT 46.330 55.600 47.780 56.470 ;
        RECT 48.090 56.590 49.040 56.670 ;
        RECT 48.090 56.420 48.120 56.590 ;
        RECT 48.290 56.420 48.480 56.590 ;
        RECT 48.650 56.420 48.840 56.590 ;
        RECT 49.010 56.420 49.040 56.590 ;
        RECT 42.850 54.470 45.950 54.510 ;
      LAYER li1 ;
        RECT 42.500 54.290 42.670 54.460 ;
      LAYER li1 ;
        RECT 44.710 54.340 45.950 54.470 ;
        RECT 39.840 53.760 41.140 54.160 ;
        RECT 39.530 53.280 41.140 53.760 ;
        RECT 41.370 53.280 42.320 54.240 ;
      LAYER li1 ;
        RECT 42.500 54.120 44.310 54.290 ;
        RECT 42.500 53.410 42.750 54.120 ;
      LAYER li1 ;
        RECT 42.930 53.280 43.880 53.940 ;
      LAYER li1 ;
        RECT 44.060 53.410 44.310 54.120 ;
      LAYER li1 ;
        RECT 44.490 53.280 45.440 54.160 ;
        RECT 45.620 53.410 45.950 54.340 ;
        RECT 46.560 54.160 46.890 54.940 ;
        RECT 47.100 54.610 47.430 55.600 ;
        RECT 48.090 55.090 49.040 56.420 ;
      LAYER li1 ;
        RECT 49.220 54.990 49.470 56.670 ;
      LAYER li1 ;
        RECT 49.650 56.590 50.600 56.670 ;
        RECT 49.650 56.420 49.680 56.590 ;
        RECT 49.850 56.420 50.040 56.590 ;
        RECT 50.210 56.420 50.400 56.590 ;
        RECT 50.570 56.420 50.600 56.590 ;
        RECT 49.650 55.170 50.600 56.420 ;
      LAYER li1 ;
        RECT 50.780 54.990 51.110 56.670 ;
      LAYER li1 ;
        RECT 51.290 56.590 52.240 56.670 ;
        RECT 51.290 56.420 51.320 56.590 ;
        RECT 51.490 56.420 51.680 56.590 ;
        RECT 51.850 56.420 52.040 56.590 ;
        RECT 52.210 56.420 52.240 56.590 ;
        RECT 51.290 55.210 52.240 56.420 ;
      LAYER li1 ;
        RECT 49.220 54.820 51.110 54.990 ;
        RECT 49.220 54.690 49.390 54.820 ;
        RECT 51.890 54.690 52.220 55.030 ;
        RECT 48.130 54.460 49.390 54.690 ;
      LAYER li1 ;
        RECT 49.570 54.510 51.600 54.640 ;
        RECT 52.420 54.510 52.670 56.670 ;
        RECT 53.050 56.640 54.500 56.670 ;
        RECT 53.050 56.470 53.300 56.640 ;
        RECT 53.470 56.470 53.660 56.640 ;
        RECT 53.830 56.470 54.100 56.640 ;
        RECT 54.270 56.470 54.500 56.640 ;
        RECT 53.050 55.600 54.500 56.470 ;
        RECT 54.810 56.590 55.760 56.670 ;
        RECT 54.810 56.420 54.840 56.590 ;
        RECT 55.010 56.420 55.200 56.590 ;
        RECT 55.370 56.420 55.560 56.590 ;
        RECT 55.730 56.420 55.760 56.590 ;
        RECT 49.570 54.470 52.670 54.510 ;
      LAYER li1 ;
        RECT 49.220 54.290 49.390 54.460 ;
      LAYER li1 ;
        RECT 51.430 54.340 52.670 54.470 ;
        RECT 46.560 53.760 47.860 54.160 ;
        RECT 46.250 53.280 47.860 53.760 ;
        RECT 48.090 53.280 49.040 54.240 ;
      LAYER li1 ;
        RECT 49.220 54.120 51.030 54.290 ;
        RECT 49.220 53.410 49.470 54.120 ;
      LAYER li1 ;
        RECT 49.650 53.280 50.600 53.940 ;
      LAYER li1 ;
        RECT 50.780 53.410 51.030 54.120 ;
      LAYER li1 ;
        RECT 51.210 53.280 52.160 54.160 ;
        RECT 52.340 53.410 52.670 54.340 ;
        RECT 53.280 54.160 53.610 54.940 ;
        RECT 53.820 54.610 54.150 55.600 ;
        RECT 54.810 55.090 55.760 56.420 ;
      LAYER li1 ;
        RECT 55.940 54.990 56.190 56.670 ;
      LAYER li1 ;
        RECT 56.370 56.590 57.320 56.670 ;
        RECT 56.370 56.420 56.400 56.590 ;
        RECT 56.570 56.420 56.760 56.590 ;
        RECT 56.930 56.420 57.120 56.590 ;
        RECT 57.290 56.420 57.320 56.590 ;
        RECT 56.370 55.170 57.320 56.420 ;
      LAYER li1 ;
        RECT 57.500 54.990 57.830 56.670 ;
      LAYER li1 ;
        RECT 58.010 56.590 58.960 56.670 ;
        RECT 58.010 56.420 58.040 56.590 ;
        RECT 58.210 56.420 58.400 56.590 ;
        RECT 58.570 56.420 58.760 56.590 ;
        RECT 58.930 56.420 58.960 56.590 ;
        RECT 58.010 55.210 58.960 56.420 ;
      LAYER li1 ;
        RECT 55.940 54.820 57.830 54.990 ;
        RECT 55.940 54.690 56.110 54.820 ;
        RECT 58.610 54.690 58.940 55.030 ;
        RECT 54.850 54.460 56.110 54.690 ;
      LAYER li1 ;
        RECT 56.290 54.510 58.320 54.640 ;
        RECT 59.140 54.510 59.390 56.670 ;
        RECT 59.770 56.640 61.220 56.670 ;
        RECT 59.770 56.470 60.020 56.640 ;
        RECT 60.190 56.470 60.380 56.640 ;
        RECT 60.550 56.470 60.820 56.640 ;
        RECT 60.990 56.470 61.220 56.640 ;
        RECT 59.770 55.600 61.220 56.470 ;
        RECT 61.530 56.590 62.480 56.670 ;
        RECT 61.530 56.420 61.560 56.590 ;
        RECT 61.730 56.420 61.920 56.590 ;
        RECT 62.090 56.420 62.280 56.590 ;
        RECT 62.450 56.420 62.480 56.590 ;
        RECT 56.290 54.470 59.390 54.510 ;
      LAYER li1 ;
        RECT 55.940 54.290 56.110 54.460 ;
      LAYER li1 ;
        RECT 58.150 54.340 59.390 54.470 ;
        RECT 53.280 53.760 54.580 54.160 ;
        RECT 52.970 53.280 54.580 53.760 ;
        RECT 54.810 53.280 55.760 54.240 ;
      LAYER li1 ;
        RECT 55.940 54.120 57.750 54.290 ;
        RECT 55.940 53.410 56.190 54.120 ;
      LAYER li1 ;
        RECT 56.370 53.280 57.320 53.940 ;
      LAYER li1 ;
        RECT 57.500 53.410 57.750 54.120 ;
      LAYER li1 ;
        RECT 57.930 53.280 58.880 54.160 ;
        RECT 59.060 53.410 59.390 54.340 ;
        RECT 60.000 54.160 60.330 54.940 ;
        RECT 60.540 54.610 60.870 55.600 ;
        RECT 61.530 55.090 62.480 56.420 ;
      LAYER li1 ;
        RECT 62.660 54.990 62.910 56.670 ;
      LAYER li1 ;
        RECT 63.090 56.590 64.040 56.670 ;
        RECT 63.090 56.420 63.120 56.590 ;
        RECT 63.290 56.420 63.480 56.590 ;
        RECT 63.650 56.420 63.840 56.590 ;
        RECT 64.010 56.420 64.040 56.590 ;
        RECT 63.090 55.170 64.040 56.420 ;
      LAYER li1 ;
        RECT 64.220 54.990 64.550 56.670 ;
      LAYER li1 ;
        RECT 64.730 56.590 65.680 56.670 ;
        RECT 64.730 56.420 64.760 56.590 ;
        RECT 64.930 56.420 65.120 56.590 ;
        RECT 65.290 56.420 65.480 56.590 ;
        RECT 65.650 56.420 65.680 56.590 ;
        RECT 64.730 55.210 65.680 56.420 ;
      LAYER li1 ;
        RECT 62.660 54.820 64.550 54.990 ;
        RECT 62.660 54.690 62.830 54.820 ;
        RECT 65.330 54.690 65.660 55.030 ;
        RECT 61.570 54.460 62.830 54.690 ;
      LAYER li1 ;
        RECT 63.010 54.510 65.040 54.640 ;
        RECT 65.860 54.510 66.110 56.670 ;
        RECT 66.490 56.640 67.940 56.670 ;
        RECT 66.490 56.470 66.740 56.640 ;
        RECT 66.910 56.470 67.100 56.640 ;
        RECT 67.270 56.470 67.540 56.640 ;
        RECT 67.710 56.470 67.940 56.640 ;
        RECT 66.490 55.600 67.940 56.470 ;
        RECT 68.250 56.590 69.200 56.670 ;
        RECT 68.250 56.420 68.280 56.590 ;
        RECT 68.450 56.420 68.640 56.590 ;
        RECT 68.810 56.420 69.000 56.590 ;
        RECT 69.170 56.420 69.200 56.590 ;
        RECT 63.010 54.470 66.110 54.510 ;
      LAYER li1 ;
        RECT 62.660 54.290 62.830 54.460 ;
      LAYER li1 ;
        RECT 64.870 54.340 66.110 54.470 ;
        RECT 60.000 53.760 61.300 54.160 ;
        RECT 59.690 53.280 61.300 53.760 ;
        RECT 61.530 53.280 62.480 54.240 ;
      LAYER li1 ;
        RECT 62.660 54.120 64.470 54.290 ;
        RECT 62.660 53.410 62.910 54.120 ;
      LAYER li1 ;
        RECT 63.090 53.280 64.040 53.940 ;
      LAYER li1 ;
        RECT 64.220 53.410 64.470 54.120 ;
      LAYER li1 ;
        RECT 64.650 53.280 65.600 54.160 ;
        RECT 65.780 53.410 66.110 54.340 ;
        RECT 66.720 54.160 67.050 54.940 ;
        RECT 67.260 54.610 67.590 55.600 ;
        RECT 68.250 55.090 69.200 56.420 ;
      LAYER li1 ;
        RECT 69.380 54.990 69.630 56.670 ;
      LAYER li1 ;
        RECT 69.810 56.590 70.760 56.670 ;
        RECT 69.810 56.420 69.840 56.590 ;
        RECT 70.010 56.420 70.200 56.590 ;
        RECT 70.370 56.420 70.560 56.590 ;
        RECT 70.730 56.420 70.760 56.590 ;
        RECT 69.810 55.170 70.760 56.420 ;
      LAYER li1 ;
        RECT 70.940 54.990 71.270 56.670 ;
      LAYER li1 ;
        RECT 71.450 56.590 72.400 56.670 ;
        RECT 71.450 56.420 71.480 56.590 ;
        RECT 71.650 56.420 71.840 56.590 ;
        RECT 72.010 56.420 72.200 56.590 ;
        RECT 72.370 56.420 72.400 56.590 ;
        RECT 71.450 55.210 72.400 56.420 ;
      LAYER li1 ;
        RECT 69.380 54.820 71.270 54.990 ;
        RECT 69.380 54.690 69.550 54.820 ;
        RECT 72.050 54.690 72.380 55.030 ;
        RECT 68.290 54.460 69.550 54.690 ;
      LAYER li1 ;
        RECT 69.730 54.510 71.760 54.640 ;
        RECT 72.580 54.510 72.830 56.670 ;
        RECT 73.210 56.640 74.660 56.670 ;
        RECT 73.210 56.470 73.460 56.640 ;
        RECT 73.630 56.470 73.820 56.640 ;
        RECT 73.990 56.470 74.260 56.640 ;
        RECT 74.430 56.470 74.660 56.640 ;
        RECT 73.210 55.600 74.660 56.470 ;
        RECT 74.970 56.590 75.920 56.670 ;
        RECT 74.970 56.420 75.000 56.590 ;
        RECT 75.170 56.420 75.360 56.590 ;
        RECT 75.530 56.420 75.720 56.590 ;
        RECT 75.890 56.420 75.920 56.590 ;
        RECT 69.730 54.470 72.830 54.510 ;
      LAYER li1 ;
        RECT 69.380 54.290 69.550 54.460 ;
      LAYER li1 ;
        RECT 71.590 54.340 72.830 54.470 ;
        RECT 66.720 53.760 68.020 54.160 ;
        RECT 66.410 53.280 68.020 53.760 ;
        RECT 68.250 53.280 69.200 54.240 ;
      LAYER li1 ;
        RECT 69.380 54.120 71.190 54.290 ;
        RECT 69.380 53.410 69.630 54.120 ;
      LAYER li1 ;
        RECT 69.810 53.280 70.760 53.940 ;
      LAYER li1 ;
        RECT 70.940 53.410 71.190 54.120 ;
      LAYER li1 ;
        RECT 71.370 53.280 72.320 54.160 ;
        RECT 72.500 53.410 72.830 54.340 ;
        RECT 73.440 54.160 73.770 54.940 ;
        RECT 73.980 54.610 74.310 55.600 ;
        RECT 74.970 55.090 75.920 56.420 ;
      LAYER li1 ;
        RECT 76.100 54.990 76.350 56.670 ;
      LAYER li1 ;
        RECT 76.530 56.590 77.480 56.670 ;
        RECT 76.530 56.420 76.560 56.590 ;
        RECT 76.730 56.420 76.920 56.590 ;
        RECT 77.090 56.420 77.280 56.590 ;
        RECT 77.450 56.420 77.480 56.590 ;
        RECT 76.530 55.170 77.480 56.420 ;
      LAYER li1 ;
        RECT 77.660 54.990 77.990 56.670 ;
      LAYER li1 ;
        RECT 78.170 56.590 79.120 56.670 ;
        RECT 78.170 56.420 78.200 56.590 ;
        RECT 78.370 56.420 78.560 56.590 ;
        RECT 78.730 56.420 78.920 56.590 ;
        RECT 79.090 56.420 79.120 56.590 ;
        RECT 78.170 55.210 79.120 56.420 ;
      LAYER li1 ;
        RECT 76.100 54.820 77.990 54.990 ;
        RECT 76.100 54.690 76.270 54.820 ;
        RECT 78.770 54.690 79.100 55.030 ;
        RECT 75.010 54.460 76.270 54.690 ;
      LAYER li1 ;
        RECT 76.450 54.510 78.480 54.640 ;
        RECT 79.300 54.510 79.550 56.670 ;
        RECT 79.930 56.640 81.380 56.670 ;
        RECT 79.930 56.470 80.180 56.640 ;
        RECT 80.350 56.470 80.540 56.640 ;
        RECT 80.710 56.470 80.980 56.640 ;
        RECT 81.150 56.470 81.380 56.640 ;
        RECT 79.930 55.600 81.380 56.470 ;
        RECT 82.650 56.590 83.600 56.670 ;
        RECT 82.650 56.420 82.680 56.590 ;
        RECT 82.850 56.420 83.040 56.590 ;
        RECT 83.210 56.420 83.400 56.590 ;
        RECT 83.570 56.420 83.600 56.590 ;
        RECT 76.450 54.470 79.550 54.510 ;
      LAYER li1 ;
        RECT 76.100 54.290 76.270 54.460 ;
      LAYER li1 ;
        RECT 78.310 54.340 79.550 54.470 ;
        RECT 73.440 53.760 74.740 54.160 ;
        RECT 73.130 53.280 74.740 53.760 ;
        RECT 74.970 53.280 75.920 54.240 ;
      LAYER li1 ;
        RECT 76.100 54.120 77.910 54.290 ;
        RECT 76.100 53.410 76.350 54.120 ;
      LAYER li1 ;
        RECT 76.530 53.280 77.480 53.940 ;
      LAYER li1 ;
        RECT 77.660 53.410 77.910 54.120 ;
      LAYER li1 ;
        RECT 78.090 53.280 79.040 54.160 ;
        RECT 79.220 53.410 79.550 54.340 ;
        RECT 80.160 54.160 80.490 54.940 ;
        RECT 80.700 54.610 81.030 55.600 ;
        RECT 82.650 55.090 83.600 56.420 ;
      LAYER li1 ;
        RECT 83.780 54.990 84.030 56.670 ;
      LAYER li1 ;
        RECT 84.210 56.590 85.160 56.670 ;
        RECT 84.210 56.420 84.240 56.590 ;
        RECT 84.410 56.420 84.600 56.590 ;
        RECT 84.770 56.420 84.960 56.590 ;
        RECT 85.130 56.420 85.160 56.590 ;
        RECT 84.210 55.170 85.160 56.420 ;
      LAYER li1 ;
        RECT 85.340 54.990 85.670 56.670 ;
      LAYER li1 ;
        RECT 85.850 56.590 86.800 56.670 ;
        RECT 85.850 56.420 85.880 56.590 ;
        RECT 86.050 56.420 86.240 56.590 ;
        RECT 86.410 56.420 86.600 56.590 ;
        RECT 86.770 56.420 86.800 56.590 ;
        RECT 85.850 55.210 86.800 56.420 ;
      LAYER li1 ;
        RECT 83.780 54.820 85.670 54.990 ;
        RECT 83.780 54.690 83.950 54.820 ;
        RECT 86.450 54.690 86.780 55.030 ;
        RECT 82.690 54.460 83.950 54.690 ;
      LAYER li1 ;
        RECT 84.130 54.510 86.160 54.640 ;
        RECT 86.980 54.510 87.230 56.670 ;
        RECT 87.610 56.640 89.060 56.670 ;
        RECT 87.610 56.470 87.860 56.640 ;
        RECT 88.030 56.470 88.220 56.640 ;
        RECT 88.390 56.470 88.660 56.640 ;
        RECT 88.830 56.470 89.060 56.640 ;
        RECT 87.610 55.600 89.060 56.470 ;
        RECT 89.370 56.590 90.630 56.670 ;
        RECT 89.370 56.420 89.380 56.590 ;
        RECT 89.550 56.420 89.740 56.590 ;
        RECT 89.910 56.420 90.100 56.590 ;
        RECT 90.270 56.420 90.460 56.590 ;
        RECT 84.130 54.470 87.230 54.510 ;
      LAYER li1 ;
        RECT 83.780 54.290 83.950 54.460 ;
      LAYER li1 ;
        RECT 85.990 54.340 87.230 54.470 ;
        RECT 80.160 53.760 81.460 54.160 ;
        RECT 79.850 53.280 81.460 53.760 ;
        RECT 82.650 53.280 83.600 54.240 ;
      LAYER li1 ;
        RECT 83.780 54.120 85.590 54.290 ;
        RECT 83.780 53.410 84.030 54.120 ;
      LAYER li1 ;
        RECT 84.210 53.280 85.160 53.940 ;
      LAYER li1 ;
        RECT 85.340 53.410 85.590 54.120 ;
      LAYER li1 ;
        RECT 85.770 53.280 86.720 54.160 ;
        RECT 86.900 53.410 87.230 54.340 ;
        RECT 87.840 54.160 88.170 54.940 ;
        RECT 88.380 54.610 88.710 55.600 ;
        RECT 89.370 55.190 90.630 56.420 ;
      LAYER li1 ;
        RECT 91.160 56.170 91.330 56.670 ;
        RECT 90.810 55.090 91.330 56.170 ;
      LAYER li1 ;
        RECT 91.590 56.590 92.900 56.670 ;
        RECT 91.590 56.420 91.620 56.590 ;
        RECT 91.790 56.420 91.980 56.590 ;
        RECT 92.150 56.420 92.340 56.590 ;
        RECT 92.510 56.420 92.700 56.590 ;
        RECT 92.870 56.420 92.900 56.590 ;
        RECT 91.590 55.210 92.900 56.420 ;
        RECT 93.370 56.640 94.820 56.670 ;
        RECT 93.370 56.470 93.620 56.640 ;
        RECT 93.790 56.470 93.980 56.640 ;
        RECT 94.150 56.470 94.420 56.640 ;
        RECT 94.590 56.470 94.820 56.640 ;
        RECT 93.370 55.600 94.820 56.470 ;
        RECT 95.190 56.550 97.000 56.720 ;
      LAYER li1 ;
        RECT 90.810 55.010 91.080 55.090 ;
        RECT 90.020 54.840 91.080 55.010 ;
        RECT 89.410 54.450 89.830 54.780 ;
        RECT 90.020 54.270 90.190 54.840 ;
        RECT 91.530 54.720 92.040 55.030 ;
        RECT 90.370 54.450 90.880 54.660 ;
      LAYER li1 ;
        RECT 91.080 54.370 92.950 54.540 ;
        RECT 87.840 53.760 89.140 54.160 ;
        RECT 87.530 53.280 89.140 53.760 ;
        RECT 89.440 53.350 89.770 54.270 ;
      LAYER li1 ;
        RECT 90.020 53.530 90.550 54.270 ;
      LAYER li1 ;
        RECT 91.080 53.350 91.250 54.370 ;
        RECT 89.440 53.180 91.250 53.350 ;
        RECT 91.430 53.280 92.530 54.190 ;
        RECT 92.700 53.440 92.950 54.370 ;
        RECT 93.600 54.160 93.930 54.940 ;
        RECT 94.140 54.610 94.470 55.600 ;
        RECT 95.190 55.090 95.520 56.550 ;
      LAYER li1 ;
        RECT 95.970 55.090 96.330 56.370 ;
        RECT 95.170 54.420 95.880 54.750 ;
      LAYER li1 ;
        RECT 93.600 53.760 94.900 54.160 ;
        RECT 93.290 53.280 94.900 53.760 ;
        RECT 95.130 53.280 95.720 54.240 ;
      LAYER li1 ;
        RECT 96.130 53.890 96.330 55.090 ;
      LAYER li1 ;
        RECT 96.750 55.010 97.000 56.550 ;
        RECT 97.180 56.590 98.130 56.670 ;
        RECT 97.180 56.420 97.210 56.590 ;
        RECT 97.380 56.420 97.570 56.590 ;
        RECT 97.740 56.420 97.930 56.590 ;
        RECT 98.100 56.420 98.130 56.590 ;
        RECT 97.180 55.190 98.130 56.420 ;
        RECT 98.310 55.010 98.640 56.670 ;
        RECT 99.130 56.640 100.580 56.670 ;
        RECT 99.130 56.470 99.380 56.640 ;
        RECT 99.550 56.470 99.740 56.640 ;
        RECT 99.910 56.470 100.180 56.640 ;
        RECT 100.350 56.470 100.580 56.640 ;
        RECT 99.130 55.600 100.580 56.470 ;
        RECT 102.330 56.590 103.280 56.670 ;
        RECT 102.330 56.420 102.360 56.590 ;
        RECT 102.530 56.420 102.720 56.590 ;
        RECT 102.890 56.420 103.080 56.590 ;
        RECT 103.250 56.420 103.280 56.590 ;
        RECT 96.750 54.840 98.640 55.010 ;
      LAYER li1 ;
        RECT 96.510 54.420 96.840 54.660 ;
        RECT 97.090 54.420 97.800 54.660 ;
        RECT 97.980 54.420 98.760 54.660 ;
        RECT 96.750 53.890 97.000 54.240 ;
        RECT 96.130 53.720 97.000 53.890 ;
        RECT 96.750 53.410 97.000 53.720 ;
      LAYER li1 ;
        RECT 97.180 53.280 98.790 54.240 ;
        RECT 99.360 54.160 99.690 54.940 ;
        RECT 99.900 54.610 100.230 55.600 ;
        RECT 102.330 55.090 103.280 56.420 ;
      LAYER li1 ;
        RECT 103.460 54.990 103.710 56.670 ;
      LAYER li1 ;
        RECT 103.890 56.590 104.840 56.670 ;
        RECT 103.890 56.420 103.920 56.590 ;
        RECT 104.090 56.420 104.280 56.590 ;
        RECT 104.450 56.420 104.640 56.590 ;
        RECT 104.810 56.420 104.840 56.590 ;
        RECT 103.890 55.170 104.840 56.420 ;
      LAYER li1 ;
        RECT 105.020 54.990 105.350 56.670 ;
      LAYER li1 ;
        RECT 105.530 56.590 106.480 56.670 ;
        RECT 105.530 56.420 105.560 56.590 ;
        RECT 105.730 56.420 105.920 56.590 ;
        RECT 106.090 56.420 106.280 56.590 ;
        RECT 106.450 56.420 106.480 56.590 ;
        RECT 105.530 55.210 106.480 56.420 ;
      LAYER li1 ;
        RECT 103.460 54.820 105.350 54.990 ;
        RECT 103.460 54.690 103.630 54.820 ;
        RECT 106.130 54.690 106.460 55.030 ;
        RECT 102.370 54.460 103.630 54.690 ;
      LAYER li1 ;
        RECT 103.810 54.510 105.840 54.640 ;
        RECT 106.660 54.510 106.910 56.670 ;
        RECT 107.290 56.640 108.740 56.670 ;
        RECT 107.290 56.470 107.540 56.640 ;
        RECT 107.710 56.470 107.900 56.640 ;
        RECT 108.070 56.470 108.340 56.640 ;
        RECT 108.510 56.470 108.740 56.640 ;
        RECT 107.290 55.600 108.740 56.470 ;
        RECT 109.050 56.590 110.000 56.670 ;
        RECT 109.050 56.420 109.080 56.590 ;
        RECT 109.250 56.420 109.440 56.590 ;
        RECT 109.610 56.420 109.800 56.590 ;
        RECT 109.970 56.420 110.000 56.590 ;
        RECT 103.810 54.470 106.910 54.510 ;
      LAYER li1 ;
        RECT 103.460 54.290 103.630 54.460 ;
      LAYER li1 ;
        RECT 105.670 54.340 106.910 54.470 ;
        RECT 99.360 53.760 100.660 54.160 ;
        RECT 99.050 53.280 100.660 53.760 ;
        RECT 102.330 53.280 103.280 54.240 ;
      LAYER li1 ;
        RECT 103.460 54.120 105.270 54.290 ;
        RECT 103.460 53.410 103.710 54.120 ;
      LAYER li1 ;
        RECT 103.890 53.280 104.840 53.940 ;
      LAYER li1 ;
        RECT 105.020 53.410 105.270 54.120 ;
      LAYER li1 ;
        RECT 105.450 53.280 106.400 54.160 ;
        RECT 106.580 53.410 106.910 54.340 ;
        RECT 107.520 54.160 107.850 54.940 ;
        RECT 108.060 54.610 108.390 55.600 ;
        RECT 109.050 55.090 110.000 56.420 ;
      LAYER li1 ;
        RECT 110.180 54.990 110.430 56.670 ;
      LAYER li1 ;
        RECT 110.610 56.590 111.560 56.670 ;
        RECT 110.610 56.420 110.640 56.590 ;
        RECT 110.810 56.420 111.000 56.590 ;
        RECT 111.170 56.420 111.360 56.590 ;
        RECT 111.530 56.420 111.560 56.590 ;
        RECT 110.610 55.170 111.560 56.420 ;
      LAYER li1 ;
        RECT 111.740 54.990 112.070 56.670 ;
      LAYER li1 ;
        RECT 112.250 56.590 113.200 56.670 ;
        RECT 112.250 56.420 112.280 56.590 ;
        RECT 112.450 56.420 112.640 56.590 ;
        RECT 112.810 56.420 113.000 56.590 ;
        RECT 113.170 56.420 113.200 56.590 ;
        RECT 112.250 55.210 113.200 56.420 ;
      LAYER li1 ;
        RECT 110.180 54.820 112.070 54.990 ;
        RECT 110.180 54.690 110.350 54.820 ;
        RECT 112.850 54.690 113.180 55.030 ;
        RECT 109.090 54.460 110.350 54.690 ;
      LAYER li1 ;
        RECT 110.530 54.510 112.560 54.640 ;
        RECT 113.380 54.510 113.630 56.670 ;
        RECT 114.010 56.640 115.460 56.670 ;
        RECT 114.010 56.470 114.260 56.640 ;
        RECT 114.430 56.470 114.620 56.640 ;
        RECT 114.790 56.470 115.060 56.640 ;
        RECT 115.230 56.470 115.460 56.640 ;
        RECT 114.010 55.600 115.460 56.470 ;
        RECT 116.250 56.590 117.200 56.670 ;
        RECT 116.250 56.420 116.280 56.590 ;
        RECT 116.450 56.420 116.640 56.590 ;
        RECT 116.810 56.420 117.000 56.590 ;
        RECT 117.170 56.420 117.200 56.590 ;
        RECT 110.530 54.470 113.630 54.510 ;
      LAYER li1 ;
        RECT 110.180 54.290 110.350 54.460 ;
      LAYER li1 ;
        RECT 112.390 54.340 113.630 54.470 ;
        RECT 107.520 53.760 108.820 54.160 ;
        RECT 107.210 53.280 108.820 53.760 ;
        RECT 109.050 53.280 110.000 54.240 ;
      LAYER li1 ;
        RECT 110.180 54.120 111.990 54.290 ;
        RECT 110.180 53.410 110.430 54.120 ;
      LAYER li1 ;
        RECT 110.610 53.280 111.560 53.940 ;
      LAYER li1 ;
        RECT 111.740 53.410 111.990 54.120 ;
      LAYER li1 ;
        RECT 112.170 53.280 113.120 54.160 ;
        RECT 113.300 53.410 113.630 54.340 ;
        RECT 114.240 54.160 114.570 54.940 ;
        RECT 114.780 54.610 115.110 55.600 ;
        RECT 116.250 55.090 117.200 56.420 ;
      LAYER li1 ;
        RECT 117.380 54.990 117.630 56.670 ;
      LAYER li1 ;
        RECT 117.810 56.590 118.760 56.670 ;
        RECT 117.810 56.420 117.840 56.590 ;
        RECT 118.010 56.420 118.200 56.590 ;
        RECT 118.370 56.420 118.560 56.590 ;
        RECT 118.730 56.420 118.760 56.590 ;
        RECT 117.810 55.170 118.760 56.420 ;
      LAYER li1 ;
        RECT 118.940 54.990 119.270 56.670 ;
      LAYER li1 ;
        RECT 119.450 56.590 120.400 56.670 ;
        RECT 119.450 56.420 119.480 56.590 ;
        RECT 119.650 56.420 119.840 56.590 ;
        RECT 120.010 56.420 120.200 56.590 ;
        RECT 120.370 56.420 120.400 56.590 ;
        RECT 119.450 55.210 120.400 56.420 ;
      LAYER li1 ;
        RECT 117.380 54.820 119.270 54.990 ;
        RECT 117.380 54.690 117.550 54.820 ;
        RECT 120.050 54.690 120.380 55.030 ;
        RECT 116.290 54.460 117.550 54.690 ;
      LAYER li1 ;
        RECT 117.730 54.510 119.760 54.640 ;
        RECT 120.580 54.510 120.830 56.670 ;
        RECT 121.210 56.640 122.660 56.670 ;
        RECT 121.210 56.470 121.460 56.640 ;
        RECT 121.630 56.470 121.820 56.640 ;
        RECT 121.990 56.470 122.260 56.640 ;
        RECT 122.430 56.470 122.660 56.640 ;
        RECT 121.210 55.600 122.660 56.470 ;
        RECT 122.970 56.590 123.920 56.670 ;
        RECT 122.970 56.420 123.000 56.590 ;
        RECT 123.170 56.420 123.360 56.590 ;
        RECT 123.530 56.420 123.720 56.590 ;
        RECT 123.890 56.420 123.920 56.590 ;
        RECT 117.730 54.470 120.830 54.510 ;
      LAYER li1 ;
        RECT 117.380 54.290 117.550 54.460 ;
      LAYER li1 ;
        RECT 119.590 54.340 120.830 54.470 ;
        RECT 114.240 53.760 115.540 54.160 ;
        RECT 113.930 53.280 115.540 53.760 ;
        RECT 116.250 53.280 117.200 54.240 ;
      LAYER li1 ;
        RECT 117.380 54.120 119.190 54.290 ;
        RECT 117.380 53.410 117.630 54.120 ;
      LAYER li1 ;
        RECT 117.810 53.280 118.760 53.940 ;
      LAYER li1 ;
        RECT 118.940 53.410 119.190 54.120 ;
      LAYER li1 ;
        RECT 119.370 53.280 120.320 54.160 ;
        RECT 120.500 53.410 120.830 54.340 ;
        RECT 121.440 54.160 121.770 54.940 ;
        RECT 121.980 54.610 122.310 55.600 ;
        RECT 122.970 55.090 123.920 56.420 ;
      LAYER li1 ;
        RECT 124.100 54.990 124.350 56.670 ;
      LAYER li1 ;
        RECT 124.530 56.590 125.480 56.670 ;
        RECT 124.530 56.420 124.560 56.590 ;
        RECT 124.730 56.420 124.920 56.590 ;
        RECT 125.090 56.420 125.280 56.590 ;
        RECT 125.450 56.420 125.480 56.590 ;
        RECT 124.530 55.170 125.480 56.420 ;
      LAYER li1 ;
        RECT 125.660 54.990 125.990 56.670 ;
      LAYER li1 ;
        RECT 126.170 56.590 127.120 56.670 ;
        RECT 126.170 56.420 126.200 56.590 ;
        RECT 126.370 56.420 126.560 56.590 ;
        RECT 126.730 56.420 126.920 56.590 ;
        RECT 127.090 56.420 127.120 56.590 ;
        RECT 126.170 55.210 127.120 56.420 ;
      LAYER li1 ;
        RECT 124.100 54.820 125.990 54.990 ;
        RECT 124.100 54.690 124.270 54.820 ;
        RECT 126.770 54.690 127.100 55.030 ;
        RECT 123.010 54.460 124.270 54.690 ;
      LAYER li1 ;
        RECT 124.450 54.510 126.480 54.640 ;
        RECT 127.300 54.510 127.550 56.670 ;
        RECT 127.930 56.640 129.380 56.670 ;
        RECT 127.930 56.470 128.180 56.640 ;
        RECT 128.350 56.470 128.540 56.640 ;
        RECT 128.710 56.470 128.980 56.640 ;
        RECT 129.150 56.470 129.380 56.640 ;
        RECT 127.930 55.600 129.380 56.470 ;
        RECT 129.690 56.590 130.640 56.670 ;
        RECT 129.690 56.420 129.720 56.590 ;
        RECT 129.890 56.420 130.080 56.590 ;
        RECT 130.250 56.420 130.440 56.590 ;
        RECT 130.610 56.420 130.640 56.590 ;
        RECT 124.450 54.470 127.550 54.510 ;
      LAYER li1 ;
        RECT 124.100 54.290 124.270 54.460 ;
      LAYER li1 ;
        RECT 126.310 54.340 127.550 54.470 ;
        RECT 121.440 53.760 122.740 54.160 ;
        RECT 121.130 53.280 122.740 53.760 ;
        RECT 122.970 53.280 123.920 54.240 ;
      LAYER li1 ;
        RECT 124.100 54.120 125.910 54.290 ;
        RECT 124.100 53.410 124.350 54.120 ;
      LAYER li1 ;
        RECT 124.530 53.280 125.480 53.940 ;
      LAYER li1 ;
        RECT 125.660 53.410 125.910 54.120 ;
      LAYER li1 ;
        RECT 126.090 53.280 127.040 54.160 ;
        RECT 127.220 53.410 127.550 54.340 ;
        RECT 128.160 54.160 128.490 54.940 ;
        RECT 128.700 54.610 129.030 55.600 ;
        RECT 129.690 55.090 130.640 56.420 ;
      LAYER li1 ;
        RECT 130.820 54.990 131.070 56.670 ;
      LAYER li1 ;
        RECT 131.250 56.590 132.200 56.670 ;
        RECT 131.250 56.420 131.280 56.590 ;
        RECT 131.450 56.420 131.640 56.590 ;
        RECT 131.810 56.420 132.000 56.590 ;
        RECT 132.170 56.420 132.200 56.590 ;
        RECT 131.250 55.170 132.200 56.420 ;
      LAYER li1 ;
        RECT 132.380 54.990 132.710 56.670 ;
      LAYER li1 ;
        RECT 132.890 56.590 133.840 56.670 ;
        RECT 132.890 56.420 132.920 56.590 ;
        RECT 133.090 56.420 133.280 56.590 ;
        RECT 133.450 56.420 133.640 56.590 ;
        RECT 133.810 56.420 133.840 56.590 ;
        RECT 132.890 55.210 133.840 56.420 ;
      LAYER li1 ;
        RECT 130.820 54.820 132.710 54.990 ;
        RECT 130.820 54.690 130.990 54.820 ;
        RECT 133.490 54.690 133.820 55.030 ;
        RECT 129.730 54.460 130.990 54.690 ;
      LAYER li1 ;
        RECT 131.170 54.510 133.200 54.640 ;
        RECT 134.020 54.510 134.270 56.670 ;
        RECT 134.650 56.640 136.100 56.670 ;
        RECT 134.650 56.470 134.900 56.640 ;
        RECT 135.070 56.470 135.260 56.640 ;
        RECT 135.430 56.470 135.700 56.640 ;
        RECT 135.870 56.470 136.100 56.640 ;
        RECT 134.650 55.600 136.100 56.470 ;
        RECT 136.410 56.590 137.670 56.670 ;
        RECT 136.410 56.420 136.420 56.590 ;
        RECT 136.590 56.420 136.780 56.590 ;
        RECT 136.950 56.420 137.140 56.590 ;
        RECT 137.310 56.420 137.500 56.590 ;
        RECT 131.170 54.470 134.270 54.510 ;
      LAYER li1 ;
        RECT 130.820 54.290 130.990 54.460 ;
      LAYER li1 ;
        RECT 133.030 54.340 134.270 54.470 ;
        RECT 128.160 53.760 129.460 54.160 ;
        RECT 127.850 53.280 129.460 53.760 ;
        RECT 129.690 53.280 130.640 54.240 ;
      LAYER li1 ;
        RECT 130.820 54.120 132.630 54.290 ;
        RECT 130.820 53.410 131.070 54.120 ;
      LAYER li1 ;
        RECT 131.250 53.280 132.200 53.940 ;
      LAYER li1 ;
        RECT 132.380 53.410 132.630 54.120 ;
      LAYER li1 ;
        RECT 132.810 53.280 133.760 54.160 ;
        RECT 133.940 53.410 134.270 54.340 ;
        RECT 134.880 54.160 135.210 54.940 ;
        RECT 135.420 54.610 135.750 55.600 ;
        RECT 136.410 55.190 137.670 56.420 ;
      LAYER li1 ;
        RECT 138.200 56.170 138.370 56.670 ;
        RECT 137.850 55.090 138.370 56.170 ;
      LAYER li1 ;
        RECT 138.630 56.590 139.940 56.670 ;
        RECT 138.630 56.420 138.660 56.590 ;
        RECT 138.830 56.420 139.020 56.590 ;
        RECT 139.190 56.420 139.380 56.590 ;
        RECT 139.550 56.420 139.740 56.590 ;
        RECT 139.910 56.420 139.940 56.590 ;
        RECT 138.630 55.210 139.940 56.420 ;
        RECT 140.410 56.640 141.860 56.670 ;
        RECT 140.410 56.470 140.660 56.640 ;
        RECT 140.830 56.470 141.020 56.640 ;
        RECT 141.190 56.470 141.460 56.640 ;
        RECT 141.630 56.470 141.860 56.640 ;
        RECT 140.410 55.600 141.860 56.470 ;
      LAYER li1 ;
        RECT 137.850 55.010 138.120 55.090 ;
        RECT 137.060 54.840 138.120 55.010 ;
        RECT 136.450 54.450 136.870 54.780 ;
        RECT 137.060 54.270 137.230 54.840 ;
        RECT 138.570 54.720 139.080 55.030 ;
        RECT 139.330 54.720 140.040 55.030 ;
        RECT 137.410 54.450 137.920 54.660 ;
      LAYER li1 ;
        RECT 138.120 54.370 139.990 54.540 ;
        RECT 134.880 53.760 136.180 54.160 ;
        RECT 134.570 53.280 136.180 53.760 ;
        RECT 136.480 53.350 136.810 54.270 ;
      LAYER li1 ;
        RECT 137.060 53.530 137.590 54.270 ;
      LAYER li1 ;
        RECT 138.120 53.350 138.290 54.370 ;
        RECT 136.480 53.180 138.290 53.350 ;
        RECT 138.470 53.280 139.570 54.190 ;
        RECT 139.740 53.440 139.990 54.370 ;
        RECT 140.640 54.160 140.970 54.940 ;
        RECT 141.180 54.610 141.510 55.600 ;
        RECT 140.640 53.760 141.940 54.160 ;
        RECT 140.330 53.280 141.940 53.760 ;
        RECT 5.760 52.820 5.920 53.000 ;
        RECT 6.090 52.820 6.400 53.000 ;
        RECT 6.570 52.820 6.880 53.000 ;
        RECT 7.050 52.820 7.360 53.000 ;
        RECT 7.530 52.820 7.680 53.000 ;
        RECT 8.160 52.820 8.320 53.000 ;
        RECT 8.490 52.820 8.800 53.000 ;
        RECT 8.970 52.820 9.280 53.000 ;
        RECT 9.450 52.820 9.760 53.000 ;
        RECT 9.930 52.820 10.240 53.000 ;
        RECT 10.410 52.820 10.720 53.000 ;
        RECT 10.890 52.820 11.200 53.000 ;
        RECT 11.370 52.820 11.680 53.000 ;
        RECT 11.850 52.820 12.160 53.000 ;
        RECT 12.330 52.820 12.640 53.000 ;
        RECT 12.810 52.820 13.120 53.000 ;
        RECT 13.290 52.820 13.600 53.000 ;
        RECT 13.770 52.820 14.080 53.000 ;
        RECT 14.250 52.820 14.560 53.000 ;
        RECT 14.730 52.820 15.040 53.000 ;
        RECT 15.210 52.820 15.520 53.000 ;
        RECT 15.690 52.820 16.000 53.000 ;
        RECT 16.170 52.820 16.480 53.000 ;
        RECT 16.650 52.820 16.960 53.000 ;
        RECT 17.130 52.820 17.440 53.000 ;
        RECT 17.610 52.820 17.920 53.000 ;
        RECT 18.090 52.820 18.400 53.000 ;
        RECT 18.570 52.820 18.880 53.000 ;
        RECT 19.050 52.820 19.360 53.000 ;
        RECT 19.530 52.820 19.840 53.000 ;
        RECT 20.010 52.820 20.320 53.000 ;
        RECT 20.490 52.820 20.800 53.000 ;
        RECT 20.970 52.820 21.280 53.000 ;
        RECT 21.450 52.820 21.760 53.000 ;
        RECT 21.930 52.820 22.240 53.000 ;
        RECT 22.410 52.820 22.720 53.000 ;
        RECT 22.890 52.820 23.200 53.000 ;
        RECT 23.370 52.820 23.680 53.000 ;
        RECT 23.850 52.820 24.160 53.000 ;
        RECT 24.330 52.820 24.640 53.000 ;
        RECT 24.810 52.820 25.120 53.000 ;
        RECT 25.290 52.820 25.600 53.000 ;
        RECT 25.770 52.820 26.080 53.000 ;
        RECT 26.250 52.820 26.560 53.000 ;
        RECT 26.730 52.820 27.040 53.000 ;
        RECT 27.210 52.820 27.520 53.000 ;
        RECT 27.690 52.820 28.000 53.000 ;
        RECT 28.170 52.820 28.480 53.000 ;
        RECT 28.650 52.820 28.960 53.000 ;
        RECT 29.130 52.820 29.440 53.000 ;
        RECT 29.610 52.820 29.920 53.000 ;
        RECT 30.090 52.820 30.400 53.000 ;
        RECT 30.570 52.820 30.880 53.000 ;
        RECT 31.050 52.820 31.360 53.000 ;
        RECT 31.530 52.820 31.840 53.000 ;
        RECT 32.010 52.820 32.320 53.000 ;
        RECT 32.490 52.820 32.800 53.000 ;
        RECT 32.970 52.820 33.280 53.000 ;
        RECT 33.450 52.820 33.760 53.000 ;
        RECT 33.930 52.820 34.240 53.000 ;
        RECT 34.410 52.820 34.720 53.000 ;
        RECT 34.890 52.820 35.200 53.000 ;
        RECT 35.370 52.820 35.680 53.000 ;
        RECT 35.850 52.820 36.160 53.000 ;
        RECT 36.330 52.820 36.640 53.000 ;
        RECT 36.810 52.820 37.120 53.000 ;
        RECT 37.290 52.820 37.600 53.000 ;
        RECT 37.770 52.820 38.080 53.000 ;
        RECT 38.250 52.820 38.560 53.000 ;
        RECT 38.730 52.820 39.040 53.000 ;
        RECT 39.210 52.820 39.520 53.000 ;
        RECT 39.690 52.820 40.000 53.000 ;
        RECT 40.170 52.820 40.480 53.000 ;
        RECT 40.650 52.820 40.960 53.000 ;
        RECT 41.130 52.820 41.440 53.000 ;
        RECT 41.610 52.820 41.920 53.000 ;
        RECT 42.090 52.820 42.400 53.000 ;
        RECT 42.570 52.820 42.880 53.000 ;
        RECT 43.050 52.820 43.360 53.000 ;
        RECT 43.530 52.820 43.840 53.000 ;
        RECT 44.010 52.820 44.320 53.000 ;
        RECT 44.490 52.820 44.800 53.000 ;
        RECT 44.970 52.820 45.280 53.000 ;
        RECT 45.450 52.820 45.760 53.000 ;
        RECT 45.930 52.820 46.240 53.000 ;
        RECT 46.410 52.820 46.720 53.000 ;
        RECT 46.890 52.820 47.200 53.000 ;
        RECT 47.370 52.820 47.520 53.000 ;
        RECT 48.000 52.820 48.160 53.000 ;
        RECT 48.330 52.820 48.640 53.000 ;
        RECT 48.810 52.820 49.120 53.000 ;
        RECT 49.290 52.820 49.600 53.000 ;
        RECT 49.770 52.820 50.080 53.000 ;
        RECT 50.250 52.820 50.560 53.000 ;
        RECT 50.730 52.820 51.040 53.000 ;
        RECT 51.210 52.820 51.520 53.000 ;
        RECT 51.690 52.820 52.000 53.000 ;
        RECT 52.170 52.820 52.480 53.000 ;
        RECT 52.650 52.820 52.960 53.000 ;
        RECT 53.130 52.820 53.440 53.000 ;
        RECT 53.610 52.820 53.920 53.000 ;
        RECT 54.090 52.820 54.400 53.000 ;
        RECT 54.570 52.820 54.880 53.000 ;
        RECT 55.050 52.820 55.360 53.000 ;
        RECT 55.530 52.820 55.840 53.000 ;
        RECT 56.010 52.820 56.320 53.000 ;
        RECT 56.490 52.820 56.800 53.000 ;
        RECT 56.970 52.820 57.280 53.000 ;
        RECT 57.450 52.820 57.760 53.000 ;
        RECT 57.930 52.820 58.240 53.000 ;
        RECT 58.410 52.820 58.720 53.000 ;
        RECT 58.890 52.820 59.200 53.000 ;
        RECT 59.370 52.820 59.680 53.000 ;
        RECT 59.850 52.820 60.160 53.000 ;
        RECT 60.330 52.820 60.640 53.000 ;
        RECT 60.810 52.820 61.120 53.000 ;
        RECT 61.290 52.820 61.600 53.000 ;
        RECT 61.770 52.820 62.080 53.000 ;
        RECT 62.250 52.820 62.560 53.000 ;
        RECT 62.730 52.820 63.040 53.000 ;
        RECT 63.210 52.820 63.520 53.000 ;
        RECT 63.690 52.820 64.000 53.000 ;
        RECT 64.170 52.820 64.480 53.000 ;
        RECT 64.650 52.820 64.960 53.000 ;
        RECT 65.130 52.820 65.440 53.000 ;
        RECT 65.610 52.820 65.920 53.000 ;
        RECT 66.090 52.820 66.400 53.000 ;
        RECT 66.570 52.820 66.880 53.000 ;
        RECT 67.050 52.820 67.360 53.000 ;
        RECT 67.530 52.820 67.840 53.000 ;
        RECT 68.010 52.820 68.320 53.000 ;
        RECT 68.490 52.820 68.800 53.000 ;
        RECT 68.970 52.820 69.280 53.000 ;
        RECT 69.450 52.820 69.760 53.000 ;
        RECT 69.930 52.820 70.240 53.000 ;
        RECT 70.410 52.820 70.720 53.000 ;
        RECT 70.890 52.820 71.200 53.000 ;
        RECT 71.370 52.820 71.680 53.000 ;
        RECT 71.850 52.820 72.160 53.000 ;
        RECT 72.330 52.820 72.640 53.000 ;
        RECT 72.810 52.820 73.120 53.000 ;
        RECT 73.290 52.820 73.600 53.000 ;
        RECT 73.770 52.820 74.080 53.000 ;
        RECT 74.250 52.820 74.560 53.000 ;
        RECT 74.730 52.820 75.040 53.000 ;
        RECT 75.210 52.820 75.520 53.000 ;
        RECT 75.690 52.820 76.000 53.000 ;
        RECT 76.170 52.820 76.480 53.000 ;
        RECT 76.650 52.820 76.960 53.000 ;
        RECT 77.130 52.820 77.440 53.000 ;
        RECT 77.610 52.820 77.920 53.000 ;
        RECT 78.090 52.820 78.400 53.000 ;
        RECT 78.570 52.820 78.880 53.000 ;
        RECT 79.050 52.820 79.360 53.000 ;
        RECT 79.530 52.820 79.840 53.000 ;
        RECT 80.010 52.820 80.320 53.000 ;
        RECT 80.490 52.820 80.800 53.000 ;
        RECT 80.970 52.820 81.120 53.000 ;
        RECT 81.600 52.820 81.760 53.000 ;
        RECT 81.930 52.820 82.240 53.000 ;
        RECT 82.410 52.820 82.720 53.000 ;
        RECT 82.890 52.820 83.200 53.000 ;
        RECT 83.370 52.820 83.680 53.000 ;
        RECT 83.850 52.820 84.160 53.000 ;
        RECT 84.330 52.820 84.640 53.000 ;
        RECT 84.810 52.820 85.120 53.000 ;
        RECT 85.290 52.820 85.600 53.000 ;
        RECT 85.770 52.820 86.080 53.000 ;
        RECT 86.250 52.820 86.560 53.000 ;
        RECT 86.730 52.820 87.040 53.000 ;
        RECT 87.210 52.820 87.520 53.000 ;
        RECT 87.690 52.820 88.000 53.000 ;
        RECT 88.170 52.820 88.480 53.000 ;
        RECT 88.650 52.820 88.960 53.000 ;
        RECT 89.130 52.820 89.440 53.000 ;
        RECT 89.610 52.820 89.920 53.000 ;
        RECT 90.090 52.820 90.400 53.000 ;
        RECT 90.570 52.820 90.880 53.000 ;
        RECT 91.050 52.820 91.360 53.000 ;
        RECT 91.530 52.820 91.840 53.000 ;
        RECT 92.010 52.820 92.320 53.000 ;
        RECT 92.490 52.820 92.800 53.000 ;
        RECT 92.970 52.820 93.280 53.000 ;
        RECT 93.450 52.820 93.760 53.000 ;
        RECT 93.930 52.820 94.240 53.000 ;
        RECT 94.410 52.820 94.720 53.000 ;
        RECT 94.890 52.820 95.200 53.000 ;
        RECT 95.370 52.820 95.680 53.000 ;
        RECT 95.850 52.820 96.160 53.000 ;
        RECT 96.330 52.820 96.640 53.000 ;
        RECT 96.810 52.820 97.120 53.000 ;
        RECT 97.290 52.820 97.600 53.000 ;
        RECT 97.770 52.820 98.080 53.000 ;
        RECT 98.250 52.820 98.560 53.000 ;
        RECT 98.730 52.820 99.040 53.000 ;
        RECT 99.210 52.820 99.520 53.000 ;
        RECT 99.690 52.820 100.000 53.000 ;
        RECT 100.170 52.820 100.480 53.000 ;
        RECT 100.650 52.820 100.960 53.000 ;
        RECT 101.130 52.820 101.440 53.000 ;
        RECT 101.610 52.820 101.920 53.000 ;
        RECT 102.090 52.820 102.400 53.000 ;
        RECT 102.570 52.820 102.880 53.000 ;
        RECT 103.050 52.820 103.360 53.000 ;
        RECT 103.530 52.820 103.840 53.000 ;
        RECT 104.010 52.820 104.320 53.000 ;
        RECT 104.490 52.820 104.800 53.000 ;
        RECT 104.970 52.820 105.280 53.000 ;
        RECT 105.450 52.820 105.760 53.000 ;
        RECT 105.930 52.820 106.240 53.000 ;
        RECT 106.410 52.820 106.720 53.000 ;
        RECT 106.890 52.820 107.040 53.000 ;
        RECT 107.520 52.820 107.680 53.000 ;
        RECT 107.850 52.820 108.160 53.000 ;
        RECT 108.330 52.820 108.640 53.000 ;
        RECT 108.810 52.820 109.120 53.000 ;
        RECT 109.290 52.820 109.600 53.000 ;
        RECT 109.770 52.820 110.080 53.000 ;
        RECT 110.250 52.820 110.560 53.000 ;
        RECT 110.730 52.820 111.040 53.000 ;
        RECT 111.210 52.820 111.520 53.000 ;
        RECT 111.690 52.820 112.000 53.000 ;
        RECT 112.170 52.820 112.480 53.000 ;
        RECT 112.650 52.820 112.960 53.000 ;
        RECT 113.130 52.820 113.440 53.000 ;
        RECT 113.610 52.820 113.920 53.000 ;
        RECT 114.090 52.820 114.400 53.000 ;
        RECT 114.570 52.820 114.880 53.000 ;
        RECT 115.050 52.820 115.360 53.000 ;
        RECT 115.530 52.820 115.840 53.000 ;
        RECT 116.010 52.820 116.320 53.000 ;
        RECT 116.490 52.820 116.800 53.000 ;
        RECT 116.970 52.820 117.280 53.000 ;
        RECT 117.450 52.820 117.760 53.000 ;
        RECT 117.930 52.820 118.240 53.000 ;
        RECT 118.410 52.820 118.720 53.000 ;
        RECT 118.890 52.820 119.200 53.000 ;
        RECT 119.370 52.820 119.680 53.000 ;
        RECT 119.850 52.820 120.160 53.000 ;
        RECT 120.330 52.820 120.640 53.000 ;
        RECT 120.810 52.820 121.120 53.000 ;
        RECT 121.290 52.820 121.600 53.000 ;
        RECT 121.770 52.820 122.080 53.000 ;
        RECT 122.250 52.820 122.560 53.000 ;
        RECT 122.730 52.820 122.880 53.000 ;
        RECT 123.360 52.820 123.520 53.000 ;
        RECT 123.690 52.820 124.000 53.000 ;
        RECT 124.170 52.820 124.480 53.000 ;
        RECT 124.650 52.820 124.960 53.000 ;
        RECT 125.130 52.820 125.440 53.000 ;
        RECT 125.610 52.820 125.920 53.000 ;
        RECT 126.090 52.820 126.400 53.000 ;
        RECT 126.570 52.820 126.880 53.000 ;
        RECT 127.050 52.820 127.360 53.000 ;
        RECT 127.530 52.820 127.840 53.000 ;
        RECT 128.010 52.820 128.320 53.000 ;
        RECT 128.490 52.820 128.800 53.000 ;
        RECT 128.970 52.820 129.280 53.000 ;
        RECT 129.450 52.820 129.760 53.000 ;
        RECT 129.930 52.820 130.240 53.000 ;
        RECT 130.410 52.820 130.720 53.000 ;
        RECT 130.890 52.820 131.200 53.000 ;
        RECT 131.370 52.820 131.680 53.000 ;
        RECT 131.850 52.820 132.160 53.000 ;
        RECT 132.330 52.820 132.640 53.000 ;
        RECT 132.810 52.820 133.120 53.000 ;
        RECT 133.290 52.820 133.600 53.000 ;
        RECT 133.770 52.820 134.080 53.000 ;
        RECT 134.250 52.820 134.560 53.000 ;
        RECT 134.730 52.820 135.040 53.000 ;
        RECT 135.210 52.820 135.520 53.000 ;
        RECT 135.690 52.820 136.000 53.000 ;
        RECT 136.170 52.820 136.480 53.000 ;
        RECT 136.650 52.820 136.960 53.000 ;
        RECT 137.130 52.820 137.440 53.000 ;
        RECT 137.610 52.820 137.920 53.000 ;
        RECT 138.090 52.820 138.400 53.000 ;
        RECT 138.570 52.820 138.880 53.000 ;
        RECT 139.050 52.820 139.360 53.000 ;
        RECT 139.530 52.820 139.840 53.000 ;
        RECT 140.010 52.820 140.320 53.000 ;
        RECT 140.490 52.820 140.800 53.000 ;
        RECT 140.970 52.820 141.280 53.000 ;
        RECT 141.450 52.820 141.760 53.000 ;
        RECT 141.930 52.820 142.080 53.000 ;
        RECT 5.930 52.510 7.540 52.540 ;
        RECT 5.930 52.340 5.980 52.510 ;
        RECT 6.150 52.340 6.420 52.510 ;
        RECT 6.590 52.340 6.860 52.510 ;
        RECT 7.030 52.340 7.270 52.510 ;
        RECT 7.440 52.340 7.540 52.510 ;
        RECT 5.930 52.060 7.540 52.340 ;
        RECT 6.240 51.660 7.540 52.060 ;
        RECT 8.250 52.510 8.840 52.540 ;
        RECT 8.250 52.340 8.280 52.510 ;
        RECT 8.450 52.340 8.640 52.510 ;
        RECT 8.810 52.340 8.840 52.510 ;
        RECT 9.770 52.510 11.380 52.540 ;
        RECT 12.070 52.510 13.320 52.540 ;
        RECT 14.090 52.510 15.700 52.540 ;
        RECT 6.240 50.880 6.570 51.660 ;
        RECT 8.250 51.580 8.840 52.340 ;
        RECT 6.780 50.220 7.110 51.210 ;
      LAYER li1 ;
        RECT 9.180 50.730 9.510 52.410 ;
      LAYER li1 ;
        RECT 9.770 52.340 9.820 52.510 ;
        RECT 9.990 52.340 10.260 52.510 ;
        RECT 10.430 52.340 10.700 52.510 ;
        RECT 10.870 52.340 11.110 52.510 ;
        RECT 11.280 52.340 11.380 52.510 ;
        RECT 9.770 52.060 11.380 52.340 ;
        RECT 10.080 51.660 11.380 52.060 ;
        RECT 10.080 50.880 10.410 51.660 ;
        RECT 6.010 49.350 7.460 50.220 ;
        RECT 6.010 49.180 6.260 49.350 ;
        RECT 6.430 49.180 6.620 49.350 ;
        RECT 6.790 49.180 7.060 49.350 ;
        RECT 7.230 49.180 7.460 49.350 ;
        RECT 6.010 49.150 7.460 49.180 ;
        RECT 8.250 49.400 8.840 50.730 ;
        RECT 8.250 49.230 8.280 49.400 ;
        RECT 8.450 49.230 8.640 49.400 ;
        RECT 8.810 49.230 8.840 49.400 ;
        RECT 8.250 49.150 8.840 49.230 ;
      LAYER li1 ;
        RECT 9.120 49.150 9.510 50.730 ;
      LAYER li1 ;
        RECT 10.620 50.220 10.950 51.210 ;
      LAYER li1 ;
        RECT 11.640 50.730 11.890 52.410 ;
      LAYER li1 ;
        RECT 12.240 52.340 12.430 52.510 ;
        RECT 12.600 52.340 12.790 52.510 ;
        RECT 12.960 52.340 13.150 52.510 ;
        RECT 12.070 51.970 13.320 52.340 ;
        RECT 13.500 51.790 13.750 52.410 ;
        RECT 14.090 52.340 14.140 52.510 ;
        RECT 14.310 52.340 14.580 52.510 ;
        RECT 14.750 52.340 15.020 52.510 ;
        RECT 15.190 52.340 15.430 52.510 ;
        RECT 15.600 52.340 15.700 52.510 ;
        RECT 14.090 52.060 15.700 52.340 ;
        RECT 12.200 51.620 13.750 51.790 ;
        RECT 12.200 51.160 12.530 51.620 ;
        RECT 9.850 49.350 11.300 50.220 ;
        RECT 9.850 49.180 10.100 49.350 ;
        RECT 10.270 49.180 10.460 49.350 ;
        RECT 10.630 49.180 10.900 49.350 ;
        RECT 11.070 49.180 11.300 49.350 ;
        RECT 9.850 49.150 11.300 49.180 ;
      LAYER li1 ;
        RECT 11.640 49.150 12.070 50.730 ;
      LAYER li1 ;
        RECT 12.250 49.400 12.810 50.730 ;
      LAYER li1 ;
        RECT 12.990 49.650 13.320 51.440 ;
      LAYER li1 ;
        RECT 13.500 49.900 13.750 51.620 ;
        RECT 14.400 51.660 15.700 52.060 ;
        RECT 15.930 52.510 17.240 52.540 ;
        RECT 15.930 52.340 15.960 52.510 ;
        RECT 16.130 52.340 16.320 52.510 ;
        RECT 16.490 52.340 16.680 52.510 ;
        RECT 16.850 52.340 17.040 52.510 ;
        RECT 17.210 52.340 17.240 52.510 ;
        RECT 18.410 52.510 20.020 52.540 ;
        RECT 14.400 50.880 14.730 51.660 ;
        RECT 15.930 51.560 17.240 52.340 ;
      LAYER li1 ;
        RECT 17.690 51.730 18.020 52.390 ;
      LAYER li1 ;
        RECT 18.410 52.340 18.460 52.510 ;
        RECT 18.630 52.340 18.900 52.510 ;
        RECT 19.070 52.340 19.340 52.510 ;
        RECT 19.510 52.340 19.750 52.510 ;
        RECT 19.920 52.340 20.020 52.510 ;
        RECT 18.410 52.060 20.020 52.340 ;
      LAYER li1 ;
        RECT 17.420 51.560 18.020 51.730 ;
      LAYER li1 ;
        RECT 18.720 51.660 20.020 52.060 ;
        RECT 20.250 52.510 20.840 52.540 ;
        RECT 22.300 52.510 23.910 52.540 ;
        RECT 24.170 52.510 25.780 52.540 ;
        RECT 20.250 52.340 20.280 52.510 ;
        RECT 20.450 52.340 20.640 52.510 ;
        RECT 20.810 52.340 20.840 52.510 ;
      LAYER li1 ;
        RECT 17.420 51.380 17.640 51.560 ;
      LAYER li1 ;
        RECT 14.940 50.220 15.270 51.210 ;
      LAYER li1 ;
        RECT 15.970 50.970 16.860 51.360 ;
        RECT 17.060 51.210 17.640 51.380 ;
      LAYER li1 ;
        RECT 12.250 49.230 12.260 49.400 ;
        RECT 12.430 49.230 12.620 49.400 ;
        RECT 12.790 49.230 12.810 49.400 ;
        RECT 12.250 49.150 12.810 49.230 ;
        RECT 14.170 49.350 15.620 50.220 ;
        RECT 14.170 49.180 14.420 49.350 ;
        RECT 14.590 49.180 14.780 49.350 ;
        RECT 14.950 49.180 15.220 49.350 ;
        RECT 15.390 49.180 15.620 49.350 ;
        RECT 14.170 49.150 15.620 49.180 ;
        RECT 15.930 49.400 16.880 50.730 ;
        RECT 15.930 49.230 15.960 49.400 ;
        RECT 16.130 49.230 16.320 49.400 ;
        RECT 16.490 49.230 16.680 49.400 ;
        RECT 16.850 49.230 16.880 49.400 ;
        RECT 15.930 49.150 16.880 49.230 ;
      LAYER li1 ;
        RECT 17.060 49.150 17.310 51.210 ;
        RECT 17.820 51.050 18.120 51.380 ;
      LAYER li1 ;
        RECT 18.720 50.880 19.050 51.660 ;
        RECT 20.250 51.580 20.840 52.340 ;
      LAYER li1 ;
        RECT 21.870 52.100 22.120 52.410 ;
      LAYER li1 ;
        RECT 22.470 52.340 22.660 52.510 ;
        RECT 22.830 52.340 23.020 52.510 ;
        RECT 23.190 52.340 23.380 52.510 ;
        RECT 23.550 52.340 23.740 52.510 ;
        RECT 24.170 52.340 24.220 52.510 ;
        RECT 24.390 52.340 24.660 52.510 ;
        RECT 24.830 52.340 25.100 52.510 ;
        RECT 25.270 52.340 25.510 52.510 ;
        RECT 25.680 52.340 25.780 52.510 ;
        RECT 26.470 52.510 27.240 52.540 ;
        RECT 28.710 52.510 29.600 52.540 ;
        RECT 30.410 52.510 32.020 52.540 ;
      LAYER li1 ;
        RECT 21.250 51.930 22.120 52.100 ;
      LAYER li1 ;
        RECT 17.500 49.400 18.090 50.730 ;
        RECT 19.260 50.220 19.590 51.210 ;
      LAYER li1 ;
        RECT 20.290 51.070 21.000 51.400 ;
        RECT 21.250 50.730 21.450 51.930 ;
        RECT 21.870 51.580 22.120 51.930 ;
      LAYER li1 ;
        RECT 22.300 51.580 23.910 52.340 ;
        RECT 24.170 52.060 25.780 52.340 ;
        RECT 24.480 51.660 25.780 52.060 ;
      LAYER li1 ;
        RECT 21.630 51.160 21.960 51.400 ;
        RECT 22.210 51.160 22.920 51.400 ;
        RECT 23.100 51.160 23.880 51.400 ;
      LAYER li1 ;
        RECT 17.500 49.230 17.530 49.400 ;
        RECT 17.700 49.230 17.890 49.400 ;
        RECT 18.060 49.230 18.090 49.400 ;
        RECT 17.500 49.150 18.090 49.230 ;
        RECT 18.490 49.350 19.940 50.220 ;
        RECT 18.490 49.180 18.740 49.350 ;
        RECT 18.910 49.180 19.100 49.350 ;
        RECT 19.270 49.180 19.540 49.350 ;
        RECT 19.710 49.180 19.940 49.350 ;
        RECT 18.490 49.150 19.940 49.180 ;
        RECT 20.310 49.270 20.640 50.730 ;
      LAYER li1 ;
        RECT 21.090 49.450 21.450 50.730 ;
      LAYER li1 ;
        RECT 21.870 50.810 23.760 50.980 ;
        RECT 24.480 50.880 24.810 51.660 ;
        RECT 21.870 49.270 22.120 50.810 ;
        RECT 20.310 49.100 22.120 49.270 ;
        RECT 22.300 49.400 23.250 50.630 ;
        RECT 22.300 49.230 22.330 49.400 ;
        RECT 22.500 49.230 22.690 49.400 ;
        RECT 22.860 49.230 23.050 49.400 ;
        RECT 23.220 49.230 23.250 49.400 ;
        RECT 22.300 49.150 23.250 49.230 ;
        RECT 23.430 49.150 23.760 50.810 ;
        RECT 25.020 50.220 25.350 51.210 ;
      LAYER li1 ;
        RECT 26.050 50.930 26.300 52.380 ;
      LAYER li1 ;
        RECT 26.470 52.340 26.520 52.510 ;
        RECT 26.690 52.340 27.030 52.510 ;
        RECT 27.200 52.340 27.240 52.510 ;
        RECT 26.470 51.630 27.240 52.340 ;
        RECT 27.420 51.450 27.750 52.410 ;
        RECT 28.200 51.800 28.530 52.410 ;
        RECT 28.880 52.340 29.070 52.510 ;
        RECT 29.240 52.340 29.430 52.510 ;
        RECT 28.710 51.980 29.600 52.340 ;
        RECT 29.780 51.800 30.110 52.410 ;
        RECT 30.410 52.340 30.460 52.510 ;
        RECT 30.630 52.340 30.900 52.510 ;
        RECT 31.070 52.340 31.340 52.510 ;
        RECT 31.510 52.340 31.750 52.510 ;
        RECT 31.920 52.340 32.020 52.510 ;
        RECT 30.410 52.060 32.020 52.340 ;
        RECT 28.200 51.630 30.110 51.800 ;
        RECT 29.780 51.580 30.110 51.630 ;
        RECT 30.720 51.660 32.020 52.060 ;
        RECT 32.250 52.510 33.200 52.540 ;
        RECT 32.250 52.340 32.280 52.510 ;
        RECT 32.450 52.340 32.640 52.510 ;
        RECT 32.810 52.340 33.000 52.510 ;
        RECT 33.170 52.340 33.200 52.510 ;
        RECT 33.810 52.510 34.760 52.540 ;
        RECT 26.470 51.280 28.300 51.450 ;
        RECT 26.470 51.110 26.760 51.280 ;
        RECT 24.250 49.350 25.700 50.220 ;
        RECT 24.250 49.180 24.500 49.350 ;
        RECT 24.670 49.180 24.860 49.350 ;
        RECT 25.030 49.180 25.300 49.350 ;
        RECT 25.470 49.180 25.700 49.350 ;
        RECT 24.250 49.150 25.700 49.180 ;
      LAYER li1 ;
        RECT 26.050 49.150 26.520 50.930 ;
        RECT 27.010 50.790 27.920 51.100 ;
      LAYER li1 ;
        RECT 26.700 49.400 27.950 50.610 ;
        RECT 26.870 49.230 27.060 49.400 ;
        RECT 27.230 49.230 27.420 49.400 ;
        RECT 27.590 49.230 27.780 49.400 ;
        RECT 26.700 49.150 27.950 49.230 ;
        RECT 28.130 49.150 28.300 51.280 ;
      LAYER li1 ;
        RECT 28.480 50.960 28.710 51.360 ;
        RECT 28.930 51.070 30.120 51.400 ;
        RECT 28.470 50.790 28.710 50.960 ;
      LAYER li1 ;
        RECT 30.720 50.880 31.050 51.660 ;
        RECT 32.250 51.580 33.200 52.340 ;
      LAYER li1 ;
        RECT 33.380 51.700 33.630 52.410 ;
      LAYER li1 ;
        RECT 33.810 52.340 33.840 52.510 ;
        RECT 34.010 52.340 34.200 52.510 ;
        RECT 34.370 52.340 34.560 52.510 ;
        RECT 34.730 52.340 34.760 52.510 ;
        RECT 35.370 52.510 36.320 52.540 ;
        RECT 33.810 51.880 34.760 52.340 ;
      LAYER li1 ;
        RECT 34.940 51.700 35.190 52.410 ;
        RECT 33.380 51.530 35.190 51.700 ;
      LAYER li1 ;
        RECT 35.370 52.340 35.400 52.510 ;
        RECT 35.570 52.340 35.760 52.510 ;
        RECT 35.930 52.340 36.120 52.510 ;
        RECT 36.290 52.340 36.320 52.510 ;
        RECT 37.130 52.510 38.740 52.540 ;
        RECT 35.370 51.660 36.320 52.340 ;
      LAYER li1 ;
        RECT 33.380 51.360 33.550 51.530 ;
      LAYER li1 ;
        RECT 36.500 51.480 36.830 52.410 ;
        RECT 37.130 52.340 37.180 52.510 ;
        RECT 37.350 52.340 37.620 52.510 ;
        RECT 37.790 52.340 38.060 52.510 ;
        RECT 38.230 52.340 38.470 52.510 ;
        RECT 38.640 52.340 38.740 52.510 ;
        RECT 37.130 52.060 38.740 52.340 ;
      LAYER li1 ;
        RECT 28.480 49.650 28.710 50.790 ;
      LAYER li1 ;
        RECT 28.890 49.400 30.150 50.730 ;
        RECT 31.260 50.220 31.590 51.210 ;
      LAYER li1 ;
        RECT 32.290 51.130 33.550 51.360 ;
      LAYER li1 ;
        RECT 35.590 51.350 36.830 51.480 ;
        RECT 33.730 51.310 36.830 51.350 ;
        RECT 33.730 51.180 35.760 51.310 ;
      LAYER li1 ;
        RECT 33.380 51.000 33.550 51.130 ;
        RECT 33.380 50.830 35.270 51.000 ;
      LAYER li1 ;
        RECT 29.060 49.230 29.250 49.400 ;
        RECT 29.420 49.230 29.610 49.400 ;
        RECT 29.780 49.230 29.970 49.400 ;
        RECT 30.140 49.230 30.150 49.400 ;
        RECT 28.890 49.150 30.150 49.230 ;
        RECT 30.490 49.350 31.940 50.220 ;
        RECT 30.490 49.180 30.740 49.350 ;
        RECT 30.910 49.180 31.100 49.350 ;
        RECT 31.270 49.180 31.540 49.350 ;
        RECT 31.710 49.180 31.940 49.350 ;
        RECT 30.490 49.150 31.940 49.180 ;
        RECT 32.250 49.400 33.200 50.730 ;
        RECT 32.250 49.230 32.280 49.400 ;
        RECT 32.450 49.230 32.640 49.400 ;
        RECT 32.810 49.230 33.000 49.400 ;
        RECT 33.170 49.230 33.200 49.400 ;
        RECT 32.250 49.150 33.200 49.230 ;
      LAYER li1 ;
        RECT 33.380 49.150 33.630 50.830 ;
      LAYER li1 ;
        RECT 33.810 49.400 34.760 50.650 ;
        RECT 33.810 49.230 33.840 49.400 ;
        RECT 34.010 49.230 34.200 49.400 ;
        RECT 34.370 49.230 34.560 49.400 ;
        RECT 34.730 49.230 34.760 49.400 ;
        RECT 33.810 49.150 34.760 49.230 ;
      LAYER li1 ;
        RECT 34.940 49.150 35.270 50.830 ;
        RECT 36.050 50.790 36.380 51.130 ;
      LAYER li1 ;
        RECT 35.450 49.400 36.400 50.610 ;
        RECT 35.450 49.230 35.480 49.400 ;
        RECT 35.650 49.230 35.840 49.400 ;
        RECT 36.010 49.230 36.200 49.400 ;
        RECT 36.370 49.230 36.400 49.400 ;
        RECT 35.450 49.150 36.400 49.230 ;
        RECT 36.580 49.150 36.830 51.310 ;
        RECT 37.440 51.660 38.740 52.060 ;
        RECT 38.970 52.510 39.920 52.540 ;
        RECT 38.970 52.340 39.000 52.510 ;
        RECT 39.170 52.340 39.360 52.510 ;
        RECT 39.530 52.340 39.720 52.510 ;
        RECT 39.890 52.340 39.920 52.510 ;
        RECT 40.530 52.510 41.480 52.540 ;
        RECT 37.440 50.880 37.770 51.660 ;
        RECT 38.970 51.580 39.920 52.340 ;
      LAYER li1 ;
        RECT 40.100 51.700 40.350 52.410 ;
      LAYER li1 ;
        RECT 40.530 52.340 40.560 52.510 ;
        RECT 40.730 52.340 40.920 52.510 ;
        RECT 41.090 52.340 41.280 52.510 ;
        RECT 41.450 52.340 41.480 52.510 ;
        RECT 42.090 52.510 43.040 52.540 ;
        RECT 40.530 51.880 41.480 52.340 ;
      LAYER li1 ;
        RECT 41.660 51.700 41.910 52.410 ;
        RECT 40.100 51.530 41.910 51.700 ;
      LAYER li1 ;
        RECT 42.090 52.340 42.120 52.510 ;
        RECT 42.290 52.340 42.480 52.510 ;
        RECT 42.650 52.340 42.840 52.510 ;
        RECT 43.010 52.340 43.040 52.510 ;
        RECT 44.260 52.520 46.990 52.550 ;
        RECT 42.090 51.660 43.040 52.340 ;
      LAYER li1 ;
        RECT 40.100 51.360 40.270 51.530 ;
      LAYER li1 ;
        RECT 43.220 51.480 43.550 52.410 ;
        RECT 44.260 52.350 44.430 52.520 ;
        RECT 44.600 52.350 44.870 52.520 ;
        RECT 45.040 52.350 45.280 52.520 ;
        RECT 45.450 52.350 45.710 52.520 ;
        RECT 45.880 52.350 46.150 52.520 ;
        RECT 46.320 52.350 46.560 52.520 ;
        RECT 46.730 52.350 46.990 52.520 ;
        RECT 44.260 51.550 46.990 52.350 ;
        RECT 48.090 52.510 49.040 52.540 ;
        RECT 48.090 52.340 48.120 52.510 ;
        RECT 48.290 52.340 48.480 52.510 ;
        RECT 48.650 52.340 48.840 52.510 ;
        RECT 49.010 52.340 49.040 52.510 ;
        RECT 49.650 52.510 50.600 52.540 ;
        RECT 48.090 51.580 49.040 52.340 ;
      LAYER li1 ;
        RECT 49.220 51.700 49.470 52.410 ;
      LAYER li1 ;
        RECT 49.650 52.340 49.680 52.510 ;
        RECT 49.850 52.340 50.040 52.510 ;
        RECT 50.210 52.340 50.400 52.510 ;
        RECT 50.570 52.340 50.600 52.510 ;
        RECT 51.210 52.510 52.160 52.540 ;
        RECT 49.650 51.880 50.600 52.340 ;
      LAYER li1 ;
        RECT 50.780 51.700 51.030 52.410 ;
      LAYER li1 ;
        RECT 37.980 50.220 38.310 51.210 ;
      LAYER li1 ;
        RECT 39.010 51.130 40.270 51.360 ;
      LAYER li1 ;
        RECT 42.310 51.350 43.550 51.480 ;
        RECT 40.450 51.310 43.550 51.350 ;
        RECT 40.450 51.180 42.480 51.310 ;
      LAYER li1 ;
        RECT 40.100 51.000 40.270 51.130 ;
        RECT 40.100 50.830 41.990 51.000 ;
      LAYER li1 ;
        RECT 37.210 49.350 38.660 50.220 ;
        RECT 37.210 49.180 37.460 49.350 ;
        RECT 37.630 49.180 37.820 49.350 ;
        RECT 37.990 49.180 38.260 49.350 ;
        RECT 38.430 49.180 38.660 49.350 ;
        RECT 37.210 49.150 38.660 49.180 ;
        RECT 38.970 49.400 39.920 50.730 ;
        RECT 38.970 49.230 39.000 49.400 ;
        RECT 39.170 49.230 39.360 49.400 ;
        RECT 39.530 49.230 39.720 49.400 ;
        RECT 39.890 49.230 39.920 49.400 ;
        RECT 38.970 49.150 39.920 49.230 ;
      LAYER li1 ;
        RECT 40.100 49.150 40.350 50.830 ;
      LAYER li1 ;
        RECT 40.530 49.400 41.480 50.650 ;
        RECT 40.530 49.230 40.560 49.400 ;
        RECT 40.730 49.230 40.920 49.400 ;
        RECT 41.090 49.230 41.280 49.400 ;
        RECT 41.450 49.230 41.480 49.400 ;
        RECT 40.530 49.150 41.480 49.230 ;
      LAYER li1 ;
        RECT 41.660 49.150 41.990 50.830 ;
        RECT 42.770 50.790 43.100 51.130 ;
      LAYER li1 ;
        RECT 42.170 49.400 43.120 50.610 ;
        RECT 42.170 49.230 42.200 49.400 ;
        RECT 42.370 49.230 42.560 49.400 ;
        RECT 42.730 49.230 42.920 49.400 ;
        RECT 43.090 49.230 43.120 49.400 ;
        RECT 42.170 49.150 43.120 49.230 ;
        RECT 43.300 49.150 43.550 51.310 ;
        RECT 44.420 50.880 44.750 51.550 ;
        RECT 45.150 50.230 45.480 51.210 ;
        RECT 45.700 50.880 46.030 51.550 ;
      LAYER li1 ;
        RECT 49.220 51.530 51.030 51.700 ;
      LAYER li1 ;
        RECT 51.210 52.340 51.240 52.510 ;
        RECT 51.410 52.340 51.600 52.510 ;
        RECT 51.770 52.340 51.960 52.510 ;
        RECT 52.130 52.340 52.160 52.510 ;
        RECT 53.380 52.520 56.110 52.550 ;
        RECT 51.210 51.660 52.160 52.340 ;
      LAYER li1 ;
        RECT 49.220 51.360 49.390 51.530 ;
      LAYER li1 ;
        RECT 52.340 51.480 52.670 52.410 ;
        RECT 53.380 52.350 53.550 52.520 ;
        RECT 53.720 52.350 53.990 52.520 ;
        RECT 54.160 52.350 54.400 52.520 ;
        RECT 54.570 52.350 54.830 52.520 ;
        RECT 55.000 52.350 55.270 52.520 ;
        RECT 55.440 52.350 55.680 52.520 ;
        RECT 55.850 52.350 56.110 52.520 ;
        RECT 53.380 51.550 56.110 52.350 ;
        RECT 57.690 52.510 58.640 52.540 ;
        RECT 57.690 52.340 57.720 52.510 ;
        RECT 57.890 52.340 58.080 52.510 ;
        RECT 58.250 52.340 58.440 52.510 ;
        RECT 58.610 52.340 58.640 52.510 ;
        RECT 59.250 52.510 60.200 52.540 ;
        RECT 57.690 51.580 58.640 52.340 ;
      LAYER li1 ;
        RECT 58.820 51.700 59.070 52.410 ;
      LAYER li1 ;
        RECT 59.250 52.340 59.280 52.510 ;
        RECT 59.450 52.340 59.640 52.510 ;
        RECT 59.810 52.340 60.000 52.510 ;
        RECT 60.170 52.340 60.200 52.510 ;
        RECT 60.810 52.510 61.760 52.540 ;
        RECT 59.250 51.880 60.200 52.340 ;
      LAYER li1 ;
        RECT 60.380 51.700 60.630 52.410 ;
      LAYER li1 ;
        RECT 46.430 50.230 46.760 51.210 ;
      LAYER li1 ;
        RECT 48.130 51.130 49.390 51.360 ;
      LAYER li1 ;
        RECT 51.430 51.350 52.670 51.480 ;
        RECT 49.570 51.310 52.670 51.350 ;
        RECT 49.570 51.180 51.600 51.310 ;
      LAYER li1 ;
        RECT 49.220 51.000 49.390 51.130 ;
        RECT 49.220 50.830 51.110 51.000 ;
      LAYER li1 ;
        RECT 44.180 49.350 46.920 50.230 ;
        RECT 44.180 49.180 44.390 49.350 ;
        RECT 44.560 49.180 44.830 49.350 ;
        RECT 45.000 49.180 45.240 49.350 ;
        RECT 45.410 49.180 45.670 49.350 ;
        RECT 45.840 49.180 46.110 49.350 ;
        RECT 46.280 49.180 46.520 49.350 ;
        RECT 46.690 49.180 46.920 49.350 ;
        RECT 44.180 49.160 46.920 49.180 ;
        RECT 48.090 49.400 49.040 50.730 ;
        RECT 48.090 49.230 48.120 49.400 ;
        RECT 48.290 49.230 48.480 49.400 ;
        RECT 48.650 49.230 48.840 49.400 ;
        RECT 49.010 49.230 49.040 49.400 ;
        RECT 48.090 49.150 49.040 49.230 ;
      LAYER li1 ;
        RECT 49.220 49.150 49.470 50.830 ;
      LAYER li1 ;
        RECT 49.650 49.400 50.600 50.650 ;
        RECT 49.650 49.230 49.680 49.400 ;
        RECT 49.850 49.230 50.040 49.400 ;
        RECT 50.210 49.230 50.400 49.400 ;
        RECT 50.570 49.230 50.600 49.400 ;
        RECT 49.650 49.150 50.600 49.230 ;
      LAYER li1 ;
        RECT 50.780 49.150 51.110 50.830 ;
        RECT 51.890 50.790 52.220 51.130 ;
      LAYER li1 ;
        RECT 51.290 49.400 52.240 50.610 ;
        RECT 51.290 49.230 51.320 49.400 ;
        RECT 51.490 49.230 51.680 49.400 ;
        RECT 51.850 49.230 52.040 49.400 ;
        RECT 52.210 49.230 52.240 49.400 ;
        RECT 51.290 49.150 52.240 49.230 ;
        RECT 52.420 49.150 52.670 51.310 ;
        RECT 53.540 50.880 53.870 51.550 ;
        RECT 54.270 50.230 54.600 51.210 ;
        RECT 54.820 50.880 55.150 51.550 ;
      LAYER li1 ;
        RECT 58.820 51.530 60.630 51.700 ;
      LAYER li1 ;
        RECT 60.810 52.340 60.840 52.510 ;
        RECT 61.010 52.340 61.200 52.510 ;
        RECT 61.370 52.340 61.560 52.510 ;
        RECT 61.730 52.340 61.760 52.510 ;
        RECT 62.570 52.510 64.180 52.540 ;
        RECT 60.810 51.660 61.760 52.340 ;
      LAYER li1 ;
        RECT 58.820 51.360 58.990 51.530 ;
      LAYER li1 ;
        RECT 61.940 51.480 62.270 52.410 ;
        RECT 62.570 52.340 62.620 52.510 ;
        RECT 62.790 52.340 63.060 52.510 ;
        RECT 63.230 52.340 63.500 52.510 ;
        RECT 63.670 52.340 63.910 52.510 ;
        RECT 64.080 52.340 64.180 52.510 ;
        RECT 62.570 52.060 64.180 52.340 ;
        RECT 55.550 50.230 55.880 51.210 ;
      LAYER li1 ;
        RECT 57.730 51.130 58.990 51.360 ;
      LAYER li1 ;
        RECT 61.030 51.350 62.270 51.480 ;
        RECT 59.170 51.310 62.270 51.350 ;
        RECT 59.170 51.180 61.200 51.310 ;
      LAYER li1 ;
        RECT 58.820 51.000 58.990 51.130 ;
        RECT 58.820 50.830 60.710 51.000 ;
      LAYER li1 ;
        RECT 53.300 49.350 56.040 50.230 ;
        RECT 53.300 49.180 53.510 49.350 ;
        RECT 53.680 49.180 53.950 49.350 ;
        RECT 54.120 49.180 54.360 49.350 ;
        RECT 54.530 49.180 54.790 49.350 ;
        RECT 54.960 49.180 55.230 49.350 ;
        RECT 55.400 49.180 55.640 49.350 ;
        RECT 55.810 49.180 56.040 49.350 ;
        RECT 53.300 49.160 56.040 49.180 ;
        RECT 57.690 49.400 58.640 50.730 ;
        RECT 57.690 49.230 57.720 49.400 ;
        RECT 57.890 49.230 58.080 49.400 ;
        RECT 58.250 49.230 58.440 49.400 ;
        RECT 58.610 49.230 58.640 49.400 ;
        RECT 57.690 49.150 58.640 49.230 ;
      LAYER li1 ;
        RECT 58.820 49.150 59.070 50.830 ;
      LAYER li1 ;
        RECT 59.250 49.400 60.200 50.650 ;
        RECT 59.250 49.230 59.280 49.400 ;
        RECT 59.450 49.230 59.640 49.400 ;
        RECT 59.810 49.230 60.000 49.400 ;
        RECT 60.170 49.230 60.200 49.400 ;
        RECT 59.250 49.150 60.200 49.230 ;
      LAYER li1 ;
        RECT 60.380 49.150 60.710 50.830 ;
        RECT 61.490 50.790 61.820 51.130 ;
      LAYER li1 ;
        RECT 60.890 49.400 61.840 50.610 ;
        RECT 60.890 49.230 60.920 49.400 ;
        RECT 61.090 49.230 61.280 49.400 ;
        RECT 61.450 49.230 61.640 49.400 ;
        RECT 61.810 49.230 61.840 49.400 ;
        RECT 60.890 49.150 61.840 49.230 ;
        RECT 62.020 49.150 62.270 51.310 ;
        RECT 62.880 51.660 64.180 52.060 ;
        RECT 64.410 52.510 65.360 52.540 ;
        RECT 64.410 52.340 64.440 52.510 ;
        RECT 64.610 52.340 64.800 52.510 ;
        RECT 64.970 52.340 65.160 52.510 ;
        RECT 65.330 52.340 65.360 52.510 ;
        RECT 65.970 52.510 66.920 52.540 ;
        RECT 62.880 50.880 63.210 51.660 ;
        RECT 64.410 51.580 65.360 52.340 ;
      LAYER li1 ;
        RECT 65.540 51.700 65.790 52.410 ;
      LAYER li1 ;
        RECT 65.970 52.340 66.000 52.510 ;
        RECT 66.170 52.340 66.360 52.510 ;
        RECT 66.530 52.340 66.720 52.510 ;
        RECT 66.890 52.340 66.920 52.510 ;
        RECT 67.530 52.510 68.480 52.540 ;
        RECT 65.970 51.880 66.920 52.340 ;
      LAYER li1 ;
        RECT 67.100 51.700 67.350 52.410 ;
        RECT 65.540 51.530 67.350 51.700 ;
      LAYER li1 ;
        RECT 67.530 52.340 67.560 52.510 ;
        RECT 67.730 52.340 67.920 52.510 ;
        RECT 68.090 52.340 68.280 52.510 ;
        RECT 68.450 52.340 68.480 52.510 ;
        RECT 69.290 52.510 70.900 52.540 ;
        RECT 67.530 51.660 68.480 52.340 ;
      LAYER li1 ;
        RECT 65.540 51.360 65.710 51.530 ;
      LAYER li1 ;
        RECT 68.660 51.480 68.990 52.410 ;
        RECT 69.290 52.340 69.340 52.510 ;
        RECT 69.510 52.340 69.780 52.510 ;
        RECT 69.950 52.340 70.220 52.510 ;
        RECT 70.390 52.340 70.630 52.510 ;
        RECT 70.800 52.340 70.900 52.510 ;
        RECT 69.290 52.060 70.900 52.340 ;
        RECT 63.420 50.220 63.750 51.210 ;
      LAYER li1 ;
        RECT 64.450 51.130 65.710 51.360 ;
      LAYER li1 ;
        RECT 67.750 51.350 68.990 51.480 ;
        RECT 65.890 51.310 68.990 51.350 ;
        RECT 65.890 51.180 67.920 51.310 ;
      LAYER li1 ;
        RECT 65.540 51.000 65.710 51.130 ;
        RECT 65.540 50.830 67.430 51.000 ;
      LAYER li1 ;
        RECT 62.650 49.350 64.100 50.220 ;
        RECT 62.650 49.180 62.900 49.350 ;
        RECT 63.070 49.180 63.260 49.350 ;
        RECT 63.430 49.180 63.700 49.350 ;
        RECT 63.870 49.180 64.100 49.350 ;
        RECT 62.650 49.150 64.100 49.180 ;
        RECT 64.410 49.400 65.360 50.730 ;
        RECT 64.410 49.230 64.440 49.400 ;
        RECT 64.610 49.230 64.800 49.400 ;
        RECT 64.970 49.230 65.160 49.400 ;
        RECT 65.330 49.230 65.360 49.400 ;
        RECT 64.410 49.150 65.360 49.230 ;
      LAYER li1 ;
        RECT 65.540 49.150 65.790 50.830 ;
      LAYER li1 ;
        RECT 65.970 49.400 66.920 50.650 ;
        RECT 65.970 49.230 66.000 49.400 ;
        RECT 66.170 49.230 66.360 49.400 ;
        RECT 66.530 49.230 66.720 49.400 ;
        RECT 66.890 49.230 66.920 49.400 ;
        RECT 65.970 49.150 66.920 49.230 ;
      LAYER li1 ;
        RECT 67.100 49.150 67.430 50.830 ;
        RECT 68.210 50.790 68.540 51.130 ;
      LAYER li1 ;
        RECT 67.610 49.400 68.560 50.610 ;
        RECT 67.610 49.230 67.640 49.400 ;
        RECT 67.810 49.230 68.000 49.400 ;
        RECT 68.170 49.230 68.360 49.400 ;
        RECT 68.530 49.230 68.560 49.400 ;
        RECT 67.610 49.150 68.560 49.230 ;
        RECT 68.740 49.150 68.990 51.310 ;
        RECT 69.600 51.660 70.900 52.060 ;
        RECT 71.130 52.510 72.080 52.540 ;
        RECT 71.130 52.340 71.160 52.510 ;
        RECT 71.330 52.340 71.520 52.510 ;
        RECT 71.690 52.340 71.880 52.510 ;
        RECT 72.050 52.340 72.080 52.510 ;
        RECT 72.690 52.510 73.640 52.540 ;
        RECT 69.600 50.880 69.930 51.660 ;
        RECT 71.130 51.580 72.080 52.340 ;
      LAYER li1 ;
        RECT 72.260 51.700 72.510 52.410 ;
      LAYER li1 ;
        RECT 72.690 52.340 72.720 52.510 ;
        RECT 72.890 52.340 73.080 52.510 ;
        RECT 73.250 52.340 73.440 52.510 ;
        RECT 73.610 52.340 73.640 52.510 ;
        RECT 74.250 52.510 75.200 52.540 ;
        RECT 72.690 51.880 73.640 52.340 ;
      LAYER li1 ;
        RECT 73.820 51.700 74.070 52.410 ;
        RECT 72.260 51.530 74.070 51.700 ;
      LAYER li1 ;
        RECT 74.250 52.340 74.280 52.510 ;
        RECT 74.450 52.340 74.640 52.510 ;
        RECT 74.810 52.340 75.000 52.510 ;
        RECT 75.170 52.340 75.200 52.510 ;
        RECT 76.010 52.510 77.620 52.540 ;
        RECT 74.250 51.660 75.200 52.340 ;
      LAYER li1 ;
        RECT 72.260 51.360 72.430 51.530 ;
      LAYER li1 ;
        RECT 75.380 51.480 75.710 52.410 ;
        RECT 76.010 52.340 76.060 52.510 ;
        RECT 76.230 52.340 76.500 52.510 ;
        RECT 76.670 52.340 76.940 52.510 ;
        RECT 77.110 52.340 77.350 52.510 ;
        RECT 77.520 52.340 77.620 52.510 ;
        RECT 76.010 52.060 77.620 52.340 ;
        RECT 70.140 50.220 70.470 51.210 ;
      LAYER li1 ;
        RECT 71.170 51.130 72.430 51.360 ;
      LAYER li1 ;
        RECT 74.470 51.350 75.710 51.480 ;
        RECT 72.610 51.310 75.710 51.350 ;
        RECT 72.610 51.180 74.640 51.310 ;
      LAYER li1 ;
        RECT 72.260 51.000 72.430 51.130 ;
        RECT 72.260 50.830 74.150 51.000 ;
      LAYER li1 ;
        RECT 69.370 49.350 70.820 50.220 ;
        RECT 69.370 49.180 69.620 49.350 ;
        RECT 69.790 49.180 69.980 49.350 ;
        RECT 70.150 49.180 70.420 49.350 ;
        RECT 70.590 49.180 70.820 49.350 ;
        RECT 69.370 49.150 70.820 49.180 ;
        RECT 71.130 49.400 72.080 50.730 ;
        RECT 71.130 49.230 71.160 49.400 ;
        RECT 71.330 49.230 71.520 49.400 ;
        RECT 71.690 49.230 71.880 49.400 ;
        RECT 72.050 49.230 72.080 49.400 ;
        RECT 71.130 49.150 72.080 49.230 ;
      LAYER li1 ;
        RECT 72.260 49.150 72.510 50.830 ;
      LAYER li1 ;
        RECT 72.690 49.400 73.640 50.650 ;
        RECT 72.690 49.230 72.720 49.400 ;
        RECT 72.890 49.230 73.080 49.400 ;
        RECT 73.250 49.230 73.440 49.400 ;
        RECT 73.610 49.230 73.640 49.400 ;
        RECT 72.690 49.150 73.640 49.230 ;
      LAYER li1 ;
        RECT 73.820 49.150 74.150 50.830 ;
        RECT 74.930 50.790 75.260 51.130 ;
      LAYER li1 ;
        RECT 74.330 49.400 75.280 50.610 ;
        RECT 74.330 49.230 74.360 49.400 ;
        RECT 74.530 49.230 74.720 49.400 ;
        RECT 74.890 49.230 75.080 49.400 ;
        RECT 75.250 49.230 75.280 49.400 ;
        RECT 74.330 49.150 75.280 49.230 ;
        RECT 75.460 49.150 75.710 51.310 ;
        RECT 76.320 51.660 77.620 52.060 ;
        RECT 77.850 52.510 78.440 52.540 ;
        RECT 77.850 52.340 77.880 52.510 ;
        RECT 78.050 52.340 78.240 52.510 ;
        RECT 78.410 52.340 78.440 52.510 ;
        RECT 79.370 52.510 80.980 52.540 ;
        RECT 76.320 50.880 76.650 51.660 ;
        RECT 77.850 51.580 78.440 52.340 ;
        RECT 76.860 50.220 77.190 51.210 ;
      LAYER li1 ;
        RECT 77.890 50.970 78.600 51.360 ;
        RECT 78.780 50.730 79.110 52.410 ;
      LAYER li1 ;
        RECT 79.370 52.340 79.420 52.510 ;
        RECT 79.590 52.340 79.860 52.510 ;
        RECT 80.030 52.340 80.300 52.510 ;
        RECT 80.470 52.340 80.710 52.510 ;
        RECT 80.880 52.340 80.980 52.510 ;
        RECT 79.370 52.060 80.980 52.340 ;
        RECT 79.680 51.660 80.980 52.060 ;
        RECT 81.690 52.510 82.640 52.540 ;
        RECT 81.690 52.340 81.720 52.510 ;
        RECT 81.890 52.340 82.080 52.510 ;
        RECT 82.250 52.340 82.440 52.510 ;
        RECT 82.610 52.340 82.640 52.510 ;
        RECT 83.250 52.510 84.200 52.540 ;
        RECT 79.680 50.880 80.010 51.660 ;
        RECT 81.690 51.580 82.640 52.340 ;
      LAYER li1 ;
        RECT 82.820 51.700 83.070 52.410 ;
      LAYER li1 ;
        RECT 83.250 52.340 83.280 52.510 ;
        RECT 83.450 52.340 83.640 52.510 ;
        RECT 83.810 52.340 84.000 52.510 ;
        RECT 84.170 52.340 84.200 52.510 ;
        RECT 84.810 52.510 85.760 52.540 ;
        RECT 83.250 51.880 84.200 52.340 ;
      LAYER li1 ;
        RECT 84.380 51.700 84.630 52.410 ;
        RECT 82.820 51.530 84.630 51.700 ;
      LAYER li1 ;
        RECT 84.810 52.340 84.840 52.510 ;
        RECT 85.010 52.340 85.200 52.510 ;
        RECT 85.370 52.340 85.560 52.510 ;
        RECT 85.730 52.340 85.760 52.510 ;
        RECT 86.570 52.510 88.180 52.540 ;
        RECT 84.810 51.660 85.760 52.340 ;
      LAYER li1 ;
        RECT 82.820 51.360 82.990 51.530 ;
      LAYER li1 ;
        RECT 85.940 51.480 86.270 52.410 ;
        RECT 86.570 52.340 86.620 52.510 ;
        RECT 86.790 52.340 87.060 52.510 ;
        RECT 87.230 52.340 87.500 52.510 ;
        RECT 87.670 52.340 87.910 52.510 ;
        RECT 88.080 52.340 88.180 52.510 ;
        RECT 86.570 52.060 88.180 52.340 ;
        RECT 76.090 49.350 77.540 50.220 ;
        RECT 76.090 49.180 76.340 49.350 ;
        RECT 76.510 49.180 76.700 49.350 ;
        RECT 76.870 49.180 77.140 49.350 ;
        RECT 77.310 49.180 77.540 49.350 ;
        RECT 76.090 49.150 77.540 49.180 ;
        RECT 77.850 49.400 78.440 50.730 ;
        RECT 77.850 49.230 77.880 49.400 ;
        RECT 78.050 49.230 78.240 49.400 ;
        RECT 78.410 49.230 78.440 49.400 ;
        RECT 77.850 49.150 78.440 49.230 ;
      LAYER li1 ;
        RECT 78.720 49.150 79.110 50.730 ;
      LAYER li1 ;
        RECT 80.220 50.220 80.550 51.210 ;
      LAYER li1 ;
        RECT 81.730 51.130 82.990 51.360 ;
      LAYER li1 ;
        RECT 85.030 51.350 86.270 51.480 ;
        RECT 83.170 51.310 86.270 51.350 ;
        RECT 83.170 51.180 85.200 51.310 ;
      LAYER li1 ;
        RECT 82.820 51.000 82.990 51.130 ;
        RECT 82.820 50.830 84.710 51.000 ;
      LAYER li1 ;
        RECT 79.450 49.350 80.900 50.220 ;
        RECT 79.450 49.180 79.700 49.350 ;
        RECT 79.870 49.180 80.060 49.350 ;
        RECT 80.230 49.180 80.500 49.350 ;
        RECT 80.670 49.180 80.900 49.350 ;
        RECT 79.450 49.150 80.900 49.180 ;
        RECT 81.690 49.400 82.640 50.730 ;
        RECT 81.690 49.230 81.720 49.400 ;
        RECT 81.890 49.230 82.080 49.400 ;
        RECT 82.250 49.230 82.440 49.400 ;
        RECT 82.610 49.230 82.640 49.400 ;
        RECT 81.690 49.150 82.640 49.230 ;
      LAYER li1 ;
        RECT 82.820 49.150 83.070 50.830 ;
      LAYER li1 ;
        RECT 83.250 49.400 84.200 50.650 ;
        RECT 83.250 49.230 83.280 49.400 ;
        RECT 83.450 49.230 83.640 49.400 ;
        RECT 83.810 49.230 84.000 49.400 ;
        RECT 84.170 49.230 84.200 49.400 ;
        RECT 83.250 49.150 84.200 49.230 ;
      LAYER li1 ;
        RECT 84.380 49.150 84.710 50.830 ;
        RECT 85.490 50.790 85.820 51.130 ;
      LAYER li1 ;
        RECT 84.890 49.400 85.840 50.610 ;
        RECT 84.890 49.230 84.920 49.400 ;
        RECT 85.090 49.230 85.280 49.400 ;
        RECT 85.450 49.230 85.640 49.400 ;
        RECT 85.810 49.230 85.840 49.400 ;
        RECT 84.890 49.150 85.840 49.230 ;
        RECT 86.020 49.150 86.270 51.310 ;
        RECT 86.880 51.660 88.180 52.060 ;
        RECT 88.410 52.510 89.360 52.540 ;
        RECT 88.410 52.340 88.440 52.510 ;
        RECT 88.610 52.340 88.800 52.510 ;
        RECT 88.970 52.340 89.160 52.510 ;
        RECT 89.330 52.340 89.360 52.510 ;
        RECT 89.970 52.510 90.920 52.540 ;
        RECT 86.880 50.880 87.210 51.660 ;
        RECT 88.410 51.580 89.360 52.340 ;
      LAYER li1 ;
        RECT 89.540 51.700 89.790 52.410 ;
      LAYER li1 ;
        RECT 89.970 52.340 90.000 52.510 ;
        RECT 90.170 52.340 90.360 52.510 ;
        RECT 90.530 52.340 90.720 52.510 ;
        RECT 90.890 52.340 90.920 52.510 ;
        RECT 91.530 52.510 92.480 52.540 ;
        RECT 89.970 51.880 90.920 52.340 ;
      LAYER li1 ;
        RECT 91.100 51.700 91.350 52.410 ;
        RECT 89.540 51.530 91.350 51.700 ;
      LAYER li1 ;
        RECT 91.530 52.340 91.560 52.510 ;
        RECT 91.730 52.340 91.920 52.510 ;
        RECT 92.090 52.340 92.280 52.510 ;
        RECT 92.450 52.340 92.480 52.510 ;
        RECT 93.290 52.510 94.900 52.540 ;
        RECT 91.530 51.660 92.480 52.340 ;
      LAYER li1 ;
        RECT 89.540 51.360 89.710 51.530 ;
      LAYER li1 ;
        RECT 92.660 51.480 92.990 52.410 ;
        RECT 93.290 52.340 93.340 52.510 ;
        RECT 93.510 52.340 93.780 52.510 ;
        RECT 93.950 52.340 94.220 52.510 ;
        RECT 94.390 52.340 94.630 52.510 ;
        RECT 94.800 52.340 94.900 52.510 ;
        RECT 93.290 52.060 94.900 52.340 ;
        RECT 87.420 50.220 87.750 51.210 ;
      LAYER li1 ;
        RECT 88.450 51.130 89.710 51.360 ;
      LAYER li1 ;
        RECT 91.750 51.350 92.990 51.480 ;
        RECT 89.890 51.310 92.990 51.350 ;
        RECT 89.890 51.180 91.920 51.310 ;
      LAYER li1 ;
        RECT 89.540 51.000 89.710 51.130 ;
        RECT 89.540 50.830 91.430 51.000 ;
      LAYER li1 ;
        RECT 86.650 49.350 88.100 50.220 ;
        RECT 86.650 49.180 86.900 49.350 ;
        RECT 87.070 49.180 87.260 49.350 ;
        RECT 87.430 49.180 87.700 49.350 ;
        RECT 87.870 49.180 88.100 49.350 ;
        RECT 86.650 49.150 88.100 49.180 ;
        RECT 88.410 49.400 89.360 50.730 ;
        RECT 88.410 49.230 88.440 49.400 ;
        RECT 88.610 49.230 88.800 49.400 ;
        RECT 88.970 49.230 89.160 49.400 ;
        RECT 89.330 49.230 89.360 49.400 ;
        RECT 88.410 49.150 89.360 49.230 ;
      LAYER li1 ;
        RECT 89.540 49.150 89.790 50.830 ;
      LAYER li1 ;
        RECT 89.970 49.400 90.920 50.650 ;
        RECT 89.970 49.230 90.000 49.400 ;
        RECT 90.170 49.230 90.360 49.400 ;
        RECT 90.530 49.230 90.720 49.400 ;
        RECT 90.890 49.230 90.920 49.400 ;
        RECT 89.970 49.150 90.920 49.230 ;
      LAYER li1 ;
        RECT 91.100 49.150 91.430 50.830 ;
        RECT 92.210 50.790 92.540 51.130 ;
      LAYER li1 ;
        RECT 91.610 49.400 92.560 50.610 ;
        RECT 91.610 49.230 91.640 49.400 ;
        RECT 91.810 49.230 92.000 49.400 ;
        RECT 92.170 49.230 92.360 49.400 ;
        RECT 92.530 49.230 92.560 49.400 ;
        RECT 91.610 49.150 92.560 49.230 ;
        RECT 92.740 49.150 92.990 51.310 ;
        RECT 93.600 51.660 94.900 52.060 ;
        RECT 95.130 52.510 95.720 52.540 ;
        RECT 95.130 52.340 95.160 52.510 ;
        RECT 95.330 52.340 95.520 52.510 ;
        RECT 95.690 52.340 95.720 52.510 ;
        RECT 96.650 52.510 98.260 52.540 ;
        RECT 93.600 50.880 93.930 51.660 ;
        RECT 95.130 51.580 95.720 52.340 ;
        RECT 94.140 50.220 94.470 51.210 ;
      LAYER li1 ;
        RECT 95.170 50.970 95.880 51.360 ;
        RECT 96.060 50.730 96.390 52.410 ;
      LAYER li1 ;
        RECT 96.650 52.340 96.700 52.510 ;
        RECT 96.870 52.340 97.140 52.510 ;
        RECT 97.310 52.340 97.580 52.510 ;
        RECT 97.750 52.340 97.990 52.510 ;
        RECT 98.160 52.340 98.260 52.510 ;
        RECT 96.650 52.060 98.260 52.340 ;
        RECT 96.960 51.660 98.260 52.060 ;
        RECT 98.490 52.510 99.440 52.540 ;
        RECT 98.490 52.340 98.520 52.510 ;
        RECT 98.690 52.340 98.880 52.510 ;
        RECT 99.050 52.340 99.240 52.510 ;
        RECT 99.410 52.340 99.440 52.510 ;
        RECT 100.050 52.510 101.000 52.540 ;
        RECT 96.960 50.880 97.290 51.660 ;
        RECT 98.490 51.580 99.440 52.340 ;
      LAYER li1 ;
        RECT 99.620 51.700 99.870 52.410 ;
      LAYER li1 ;
        RECT 100.050 52.340 100.080 52.510 ;
        RECT 100.250 52.340 100.440 52.510 ;
        RECT 100.610 52.340 100.800 52.510 ;
        RECT 100.970 52.340 101.000 52.510 ;
        RECT 101.610 52.510 102.560 52.540 ;
        RECT 100.050 51.880 101.000 52.340 ;
      LAYER li1 ;
        RECT 101.180 51.700 101.430 52.410 ;
        RECT 99.620 51.530 101.430 51.700 ;
      LAYER li1 ;
        RECT 101.610 52.340 101.640 52.510 ;
        RECT 101.810 52.340 102.000 52.510 ;
        RECT 102.170 52.340 102.360 52.510 ;
        RECT 102.530 52.340 102.560 52.510 ;
        RECT 103.780 52.520 106.510 52.550 ;
        RECT 101.610 51.660 102.560 52.340 ;
      LAYER li1 ;
        RECT 99.620 51.360 99.790 51.530 ;
      LAYER li1 ;
        RECT 102.740 51.480 103.070 52.410 ;
        RECT 103.780 52.350 103.950 52.520 ;
        RECT 104.120 52.350 104.390 52.520 ;
        RECT 104.560 52.350 104.800 52.520 ;
        RECT 104.970 52.350 105.230 52.520 ;
        RECT 105.400 52.350 105.670 52.520 ;
        RECT 105.840 52.350 106.080 52.520 ;
        RECT 106.250 52.350 106.510 52.520 ;
        RECT 103.780 51.550 106.510 52.350 ;
        RECT 107.610 52.510 108.560 52.540 ;
        RECT 107.610 52.340 107.640 52.510 ;
        RECT 107.810 52.340 108.000 52.510 ;
        RECT 108.170 52.340 108.360 52.510 ;
        RECT 108.530 52.340 108.560 52.510 ;
        RECT 109.170 52.510 110.120 52.540 ;
        RECT 107.610 51.580 108.560 52.340 ;
      LAYER li1 ;
        RECT 108.740 51.700 108.990 52.410 ;
      LAYER li1 ;
        RECT 109.170 52.340 109.200 52.510 ;
        RECT 109.370 52.340 109.560 52.510 ;
        RECT 109.730 52.340 109.920 52.510 ;
        RECT 110.090 52.340 110.120 52.510 ;
        RECT 110.730 52.510 111.680 52.540 ;
        RECT 109.170 51.880 110.120 52.340 ;
      LAYER li1 ;
        RECT 110.300 51.700 110.550 52.410 ;
      LAYER li1 ;
        RECT 93.370 49.350 94.820 50.220 ;
        RECT 93.370 49.180 93.620 49.350 ;
        RECT 93.790 49.180 93.980 49.350 ;
        RECT 94.150 49.180 94.420 49.350 ;
        RECT 94.590 49.180 94.820 49.350 ;
        RECT 93.370 49.150 94.820 49.180 ;
        RECT 95.130 49.400 95.720 50.730 ;
        RECT 95.130 49.230 95.160 49.400 ;
        RECT 95.330 49.230 95.520 49.400 ;
        RECT 95.690 49.230 95.720 49.400 ;
        RECT 95.130 49.150 95.720 49.230 ;
      LAYER li1 ;
        RECT 96.000 49.150 96.390 50.730 ;
      LAYER li1 ;
        RECT 97.500 50.220 97.830 51.210 ;
      LAYER li1 ;
        RECT 98.530 51.130 99.790 51.360 ;
      LAYER li1 ;
        RECT 101.830 51.350 103.070 51.480 ;
        RECT 99.970 51.310 103.070 51.350 ;
        RECT 99.970 51.180 102.000 51.310 ;
      LAYER li1 ;
        RECT 99.620 51.000 99.790 51.130 ;
        RECT 99.620 50.830 101.510 51.000 ;
      LAYER li1 ;
        RECT 96.730 49.350 98.180 50.220 ;
        RECT 96.730 49.180 96.980 49.350 ;
        RECT 97.150 49.180 97.340 49.350 ;
        RECT 97.510 49.180 97.780 49.350 ;
        RECT 97.950 49.180 98.180 49.350 ;
        RECT 96.730 49.150 98.180 49.180 ;
        RECT 98.490 49.400 99.440 50.730 ;
        RECT 98.490 49.230 98.520 49.400 ;
        RECT 98.690 49.230 98.880 49.400 ;
        RECT 99.050 49.230 99.240 49.400 ;
        RECT 99.410 49.230 99.440 49.400 ;
        RECT 98.490 49.150 99.440 49.230 ;
      LAYER li1 ;
        RECT 99.620 49.150 99.870 50.830 ;
      LAYER li1 ;
        RECT 100.050 49.400 101.000 50.650 ;
        RECT 100.050 49.230 100.080 49.400 ;
        RECT 100.250 49.230 100.440 49.400 ;
        RECT 100.610 49.230 100.800 49.400 ;
        RECT 100.970 49.230 101.000 49.400 ;
        RECT 100.050 49.150 101.000 49.230 ;
      LAYER li1 ;
        RECT 101.180 49.150 101.510 50.830 ;
        RECT 102.290 50.790 102.620 51.130 ;
      LAYER li1 ;
        RECT 101.690 49.400 102.640 50.610 ;
        RECT 101.690 49.230 101.720 49.400 ;
        RECT 101.890 49.230 102.080 49.400 ;
        RECT 102.250 49.230 102.440 49.400 ;
        RECT 102.610 49.230 102.640 49.400 ;
        RECT 101.690 49.150 102.640 49.230 ;
        RECT 102.820 49.150 103.070 51.310 ;
        RECT 103.940 50.880 104.270 51.550 ;
        RECT 104.670 50.230 105.000 51.210 ;
        RECT 105.220 50.880 105.550 51.550 ;
      LAYER li1 ;
        RECT 108.740 51.530 110.550 51.700 ;
      LAYER li1 ;
        RECT 110.730 52.340 110.760 52.510 ;
        RECT 110.930 52.340 111.120 52.510 ;
        RECT 111.290 52.340 111.480 52.510 ;
        RECT 111.650 52.340 111.680 52.510 ;
        RECT 112.490 52.510 114.100 52.540 ;
        RECT 110.730 51.660 111.680 52.340 ;
      LAYER li1 ;
        RECT 108.740 51.360 108.910 51.530 ;
      LAYER li1 ;
        RECT 111.860 51.480 112.190 52.410 ;
        RECT 112.490 52.340 112.540 52.510 ;
        RECT 112.710 52.340 112.980 52.510 ;
        RECT 113.150 52.340 113.420 52.510 ;
        RECT 113.590 52.340 113.830 52.510 ;
        RECT 114.000 52.340 114.100 52.510 ;
        RECT 112.490 52.060 114.100 52.340 ;
        RECT 105.950 50.230 106.280 51.210 ;
      LAYER li1 ;
        RECT 107.650 51.130 108.910 51.360 ;
      LAYER li1 ;
        RECT 110.950 51.350 112.190 51.480 ;
        RECT 109.090 51.310 112.190 51.350 ;
        RECT 109.090 51.180 111.120 51.310 ;
      LAYER li1 ;
        RECT 108.740 51.000 108.910 51.130 ;
        RECT 108.740 50.830 110.630 51.000 ;
      LAYER li1 ;
        RECT 103.700 49.350 106.440 50.230 ;
        RECT 103.700 49.180 103.910 49.350 ;
        RECT 104.080 49.180 104.350 49.350 ;
        RECT 104.520 49.180 104.760 49.350 ;
        RECT 104.930 49.180 105.190 49.350 ;
        RECT 105.360 49.180 105.630 49.350 ;
        RECT 105.800 49.180 106.040 49.350 ;
        RECT 106.210 49.180 106.440 49.350 ;
        RECT 103.700 49.160 106.440 49.180 ;
        RECT 107.610 49.400 108.560 50.730 ;
        RECT 107.610 49.230 107.640 49.400 ;
        RECT 107.810 49.230 108.000 49.400 ;
        RECT 108.170 49.230 108.360 49.400 ;
        RECT 108.530 49.230 108.560 49.400 ;
        RECT 107.610 49.150 108.560 49.230 ;
      LAYER li1 ;
        RECT 108.740 49.150 108.990 50.830 ;
      LAYER li1 ;
        RECT 109.170 49.400 110.120 50.650 ;
        RECT 109.170 49.230 109.200 49.400 ;
        RECT 109.370 49.230 109.560 49.400 ;
        RECT 109.730 49.230 109.920 49.400 ;
        RECT 110.090 49.230 110.120 49.400 ;
        RECT 109.170 49.150 110.120 49.230 ;
      LAYER li1 ;
        RECT 110.300 49.150 110.630 50.830 ;
        RECT 111.410 50.790 111.740 51.130 ;
      LAYER li1 ;
        RECT 110.810 49.400 111.760 50.610 ;
        RECT 110.810 49.230 110.840 49.400 ;
        RECT 111.010 49.230 111.200 49.400 ;
        RECT 111.370 49.230 111.560 49.400 ;
        RECT 111.730 49.230 111.760 49.400 ;
        RECT 110.810 49.150 111.760 49.230 ;
        RECT 111.940 49.150 112.190 51.310 ;
        RECT 112.800 51.660 114.100 52.060 ;
        RECT 114.330 52.510 115.280 52.540 ;
        RECT 114.330 52.340 114.360 52.510 ;
        RECT 114.530 52.340 114.720 52.510 ;
        RECT 114.890 52.340 115.080 52.510 ;
        RECT 115.250 52.340 115.280 52.510 ;
        RECT 115.890 52.510 116.840 52.540 ;
        RECT 112.800 50.880 113.130 51.660 ;
        RECT 114.330 51.580 115.280 52.340 ;
      LAYER li1 ;
        RECT 115.460 51.700 115.710 52.410 ;
      LAYER li1 ;
        RECT 115.890 52.340 115.920 52.510 ;
        RECT 116.090 52.340 116.280 52.510 ;
        RECT 116.450 52.340 116.640 52.510 ;
        RECT 116.810 52.340 116.840 52.510 ;
        RECT 117.450 52.510 118.400 52.540 ;
        RECT 115.890 51.880 116.840 52.340 ;
      LAYER li1 ;
        RECT 117.020 51.700 117.270 52.410 ;
        RECT 115.460 51.530 117.270 51.700 ;
      LAYER li1 ;
        RECT 117.450 52.340 117.480 52.510 ;
        RECT 117.650 52.340 117.840 52.510 ;
        RECT 118.010 52.340 118.200 52.510 ;
        RECT 118.370 52.340 118.400 52.510 ;
        RECT 119.620 52.520 122.350 52.550 ;
        RECT 117.450 51.660 118.400 52.340 ;
      LAYER li1 ;
        RECT 115.460 51.360 115.630 51.530 ;
      LAYER li1 ;
        RECT 118.580 51.480 118.910 52.410 ;
        RECT 119.620 52.350 119.790 52.520 ;
        RECT 119.960 52.350 120.230 52.520 ;
        RECT 120.400 52.350 120.640 52.520 ;
        RECT 120.810 52.350 121.070 52.520 ;
        RECT 121.240 52.350 121.510 52.520 ;
        RECT 121.680 52.350 121.920 52.520 ;
        RECT 122.090 52.350 122.350 52.520 ;
        RECT 123.970 52.510 125.770 52.540 ;
        RECT 126.460 52.510 126.990 52.540 ;
        RECT 128.810 52.510 130.420 52.540 ;
        RECT 119.620 51.550 122.350 52.350 ;
        RECT 123.470 51.680 123.800 52.410 ;
        RECT 123.970 52.340 124.160 52.510 ;
        RECT 124.330 52.340 124.520 52.510 ;
        RECT 124.690 52.340 124.880 52.510 ;
        RECT 125.050 52.340 125.240 52.510 ;
        RECT 125.410 52.340 125.600 52.510 ;
        RECT 123.970 51.860 125.770 52.340 ;
        RECT 125.950 51.800 126.280 52.410 ;
        RECT 126.630 52.340 126.820 52.510 ;
        RECT 126.460 51.980 126.990 52.340 ;
        RECT 127.330 51.800 127.660 52.370 ;
        RECT 113.340 50.220 113.670 51.210 ;
      LAYER li1 ;
        RECT 114.370 51.130 115.630 51.360 ;
      LAYER li1 ;
        RECT 117.670 51.350 118.910 51.480 ;
        RECT 115.810 51.310 118.910 51.350 ;
        RECT 115.810 51.180 117.840 51.310 ;
      LAYER li1 ;
        RECT 115.460 51.000 115.630 51.130 ;
        RECT 115.460 50.830 117.350 51.000 ;
      LAYER li1 ;
        RECT 112.570 49.350 114.020 50.220 ;
        RECT 112.570 49.180 112.820 49.350 ;
        RECT 112.990 49.180 113.180 49.350 ;
        RECT 113.350 49.180 113.620 49.350 ;
        RECT 113.790 49.180 114.020 49.350 ;
        RECT 112.570 49.150 114.020 49.180 ;
        RECT 114.330 49.400 115.280 50.730 ;
        RECT 114.330 49.230 114.360 49.400 ;
        RECT 114.530 49.230 114.720 49.400 ;
        RECT 114.890 49.230 115.080 49.400 ;
        RECT 115.250 49.230 115.280 49.400 ;
        RECT 114.330 49.150 115.280 49.230 ;
      LAYER li1 ;
        RECT 115.460 49.150 115.710 50.830 ;
      LAYER li1 ;
        RECT 115.890 49.400 116.840 50.650 ;
        RECT 115.890 49.230 115.920 49.400 ;
        RECT 116.090 49.230 116.280 49.400 ;
        RECT 116.450 49.230 116.640 49.400 ;
        RECT 116.810 49.230 116.840 49.400 ;
        RECT 115.890 49.150 116.840 49.230 ;
      LAYER li1 ;
        RECT 117.020 49.150 117.350 50.830 ;
        RECT 118.130 50.790 118.460 51.130 ;
      LAYER li1 ;
        RECT 117.530 49.400 118.480 50.610 ;
        RECT 117.530 49.230 117.560 49.400 ;
        RECT 117.730 49.230 117.920 49.400 ;
        RECT 118.090 49.230 118.280 49.400 ;
        RECT 118.450 49.230 118.480 49.400 ;
        RECT 117.530 49.150 118.480 49.230 ;
        RECT 118.660 49.150 118.910 51.310 ;
        RECT 119.780 50.880 120.110 51.550 ;
        RECT 120.510 50.230 120.840 51.210 ;
        RECT 121.060 50.880 121.390 51.550 ;
        RECT 123.470 51.510 125.770 51.680 ;
        RECT 125.950 51.620 127.660 51.800 ;
        RECT 121.790 50.230 122.120 51.210 ;
        RECT 123.470 50.630 123.720 51.510 ;
        RECT 125.600 51.450 125.770 51.510 ;
      LAYER li1 ;
        RECT 123.940 50.980 124.270 51.180 ;
        RECT 124.450 51.160 125.420 51.330 ;
      LAYER li1 ;
        RECT 125.600 51.280 127.340 51.450 ;
      LAYER li1 ;
        RECT 128.110 51.360 128.520 52.370 ;
      LAYER li1 ;
        RECT 128.810 52.340 128.860 52.510 ;
        RECT 129.030 52.340 129.300 52.510 ;
        RECT 129.470 52.340 129.740 52.510 ;
        RECT 129.910 52.340 130.150 52.510 ;
        RECT 130.320 52.340 130.420 52.510 ;
        RECT 128.810 52.060 130.420 52.340 ;
        RECT 127.010 51.180 127.340 51.280 ;
      LAYER li1 ;
        RECT 126.290 50.980 126.620 51.100 ;
        RECT 127.810 51.000 128.520 51.360 ;
        RECT 123.940 50.810 126.620 50.980 ;
        RECT 124.930 50.790 126.620 50.810 ;
        RECT 127.390 50.830 128.520 51.000 ;
      LAYER li1 ;
        RECT 129.120 51.660 130.420 52.060 ;
        RECT 130.650 52.510 131.600 52.540 ;
        RECT 130.650 52.340 130.680 52.510 ;
        RECT 130.850 52.340 131.040 52.510 ;
        RECT 131.210 52.340 131.400 52.510 ;
        RECT 131.570 52.340 131.600 52.510 ;
        RECT 132.210 52.510 133.160 52.540 ;
        RECT 129.120 50.880 129.450 51.660 ;
        RECT 130.650 51.580 131.600 52.340 ;
      LAYER li1 ;
        RECT 131.780 51.700 132.030 52.410 ;
      LAYER li1 ;
        RECT 132.210 52.340 132.240 52.510 ;
        RECT 132.410 52.340 132.600 52.510 ;
        RECT 132.770 52.340 132.960 52.510 ;
        RECT 133.130 52.340 133.160 52.510 ;
        RECT 133.770 52.510 134.720 52.540 ;
        RECT 132.210 51.880 133.160 52.340 ;
      LAYER li1 ;
        RECT 133.340 51.700 133.590 52.410 ;
        RECT 131.780 51.530 133.590 51.700 ;
      LAYER li1 ;
        RECT 133.770 52.340 133.800 52.510 ;
        RECT 133.970 52.340 134.160 52.510 ;
        RECT 134.330 52.340 134.520 52.510 ;
        RECT 134.690 52.340 134.720 52.510 ;
        RECT 135.530 52.510 137.140 52.540 ;
        RECT 133.770 51.660 134.720 52.340 ;
      LAYER li1 ;
        RECT 131.780 51.360 131.950 51.530 ;
      LAYER li1 ;
        RECT 134.900 51.480 135.230 52.410 ;
        RECT 135.530 52.340 135.580 52.510 ;
        RECT 135.750 52.340 136.020 52.510 ;
        RECT 136.190 52.340 136.460 52.510 ;
        RECT 136.630 52.340 136.870 52.510 ;
        RECT 137.040 52.340 137.140 52.510 ;
        RECT 135.530 52.060 137.140 52.340 ;
        RECT 123.470 50.460 124.700 50.630 ;
        RECT 119.540 49.350 122.280 50.230 ;
        RECT 119.540 49.180 119.750 49.350 ;
        RECT 119.920 49.180 120.190 49.350 ;
        RECT 120.360 49.180 120.600 49.350 ;
        RECT 120.770 49.180 121.030 49.350 ;
        RECT 121.200 49.180 121.470 49.350 ;
        RECT 121.640 49.180 121.880 49.350 ;
        RECT 122.050 49.180 122.280 49.350 ;
        RECT 119.540 49.160 122.280 49.180 ;
        RECT 123.450 49.400 124.350 50.280 ;
        RECT 123.450 49.230 123.460 49.400 ;
        RECT 123.630 49.230 123.820 49.400 ;
        RECT 123.990 49.230 124.180 49.400 ;
        RECT 123.450 49.150 124.350 49.230 ;
        RECT 124.530 49.150 124.700 50.460 ;
        RECT 124.880 49.400 127.210 50.610 ;
        RECT 125.050 49.230 125.240 49.400 ;
        RECT 125.410 49.230 125.600 49.400 ;
        RECT 125.770 49.230 125.960 49.400 ;
        RECT 126.130 49.230 126.320 49.400 ;
        RECT 126.490 49.230 126.680 49.400 ;
        RECT 126.850 49.230 127.040 49.400 ;
        RECT 124.880 49.150 127.210 49.230 ;
      LAYER li1 ;
        RECT 127.390 49.150 127.640 50.830 ;
      LAYER li1 ;
        RECT 127.830 49.400 128.420 50.650 ;
        RECT 129.660 50.220 129.990 51.210 ;
      LAYER li1 ;
        RECT 130.690 51.130 131.950 51.360 ;
      LAYER li1 ;
        RECT 133.990 51.350 135.230 51.480 ;
        RECT 132.130 51.310 135.230 51.350 ;
        RECT 132.130 51.180 134.160 51.310 ;
      LAYER li1 ;
        RECT 131.780 51.000 131.950 51.130 ;
        RECT 131.780 50.830 133.670 51.000 ;
      LAYER li1 ;
        RECT 127.830 49.230 127.860 49.400 ;
        RECT 128.030 49.230 128.220 49.400 ;
        RECT 128.390 49.230 128.420 49.400 ;
        RECT 127.830 49.150 128.420 49.230 ;
        RECT 128.890 49.350 130.340 50.220 ;
        RECT 128.890 49.180 129.140 49.350 ;
        RECT 129.310 49.180 129.500 49.350 ;
        RECT 129.670 49.180 129.940 49.350 ;
        RECT 130.110 49.180 130.340 49.350 ;
        RECT 128.890 49.150 130.340 49.180 ;
        RECT 130.650 49.400 131.600 50.730 ;
        RECT 130.650 49.230 130.680 49.400 ;
        RECT 130.850 49.230 131.040 49.400 ;
        RECT 131.210 49.230 131.400 49.400 ;
        RECT 131.570 49.230 131.600 49.400 ;
        RECT 130.650 49.150 131.600 49.230 ;
      LAYER li1 ;
        RECT 131.780 49.150 132.030 50.830 ;
      LAYER li1 ;
        RECT 132.210 49.400 133.160 50.650 ;
        RECT 132.210 49.230 132.240 49.400 ;
        RECT 132.410 49.230 132.600 49.400 ;
        RECT 132.770 49.230 132.960 49.400 ;
        RECT 133.130 49.230 133.160 49.400 ;
        RECT 132.210 49.150 133.160 49.230 ;
      LAYER li1 ;
        RECT 133.340 49.150 133.670 50.830 ;
        RECT 134.450 50.790 134.780 51.130 ;
      LAYER li1 ;
        RECT 133.850 49.400 134.800 50.610 ;
        RECT 133.850 49.230 133.880 49.400 ;
        RECT 134.050 49.230 134.240 49.400 ;
        RECT 134.410 49.230 134.600 49.400 ;
        RECT 134.770 49.230 134.800 49.400 ;
        RECT 133.850 49.150 134.800 49.230 ;
        RECT 134.980 49.150 135.230 51.310 ;
        RECT 135.840 51.660 137.140 52.060 ;
        RECT 137.370 52.510 138.300 52.540 ;
        RECT 137.370 52.340 137.390 52.510 ;
        RECT 137.560 52.340 137.750 52.510 ;
        RECT 137.920 52.340 138.110 52.510 ;
        RECT 138.280 52.340 138.300 52.510 ;
        RECT 139.000 52.510 139.590 52.540 ;
        RECT 135.840 50.880 136.170 51.660 ;
        RECT 137.370 51.580 138.300 52.340 ;
      LAYER li1 ;
        RECT 138.480 51.480 138.810 52.410 ;
      LAYER li1 ;
        RECT 139.000 52.340 139.030 52.510 ;
        RECT 139.200 52.340 139.390 52.510 ;
        RECT 139.560 52.340 139.590 52.510 ;
        RECT 139.000 51.660 139.590 52.340 ;
        RECT 139.850 52.510 141.460 52.540 ;
        RECT 139.850 52.340 139.900 52.510 ;
        RECT 140.070 52.340 140.340 52.510 ;
        RECT 140.510 52.340 140.780 52.510 ;
        RECT 140.950 52.340 141.190 52.510 ;
        RECT 141.360 52.340 141.460 52.510 ;
        RECT 139.850 52.060 141.460 52.340 ;
        RECT 140.160 51.660 141.460 52.060 ;
      LAYER li1 ;
        RECT 138.480 51.310 139.560 51.480 ;
      LAYER li1 ;
        RECT 136.380 50.220 136.710 51.210 ;
      LAYER li1 ;
        RECT 137.410 50.790 138.600 51.130 ;
        RECT 138.780 50.790 139.110 51.130 ;
      LAYER li1 ;
        RECT 135.610 49.350 137.060 50.220 ;
        RECT 135.610 49.180 135.860 49.350 ;
        RECT 136.030 49.180 136.220 49.350 ;
        RECT 136.390 49.180 136.660 49.350 ;
        RECT 136.830 49.180 137.060 49.350 ;
        RECT 135.610 49.150 137.060 49.180 ;
        RECT 137.370 49.400 139.040 50.610 ;
        RECT 137.370 49.230 137.400 49.400 ;
        RECT 137.570 49.230 137.760 49.400 ;
        RECT 137.930 49.230 138.120 49.400 ;
        RECT 138.290 49.230 138.480 49.400 ;
        RECT 138.650 49.230 138.840 49.400 ;
        RECT 139.010 49.230 139.040 49.400 ;
        RECT 137.370 49.150 139.040 49.230 ;
      LAYER li1 ;
        RECT 139.300 49.150 139.560 51.310 ;
      LAYER li1 ;
        RECT 140.160 50.880 140.490 51.660 ;
        RECT 140.700 50.220 141.030 51.210 ;
        RECT 139.930 49.350 141.380 50.220 ;
        RECT 139.930 49.180 140.180 49.350 ;
        RECT 140.350 49.180 140.540 49.350 ;
        RECT 140.710 49.180 140.980 49.350 ;
        RECT 141.150 49.180 141.380 49.350 ;
        RECT 139.930 49.150 141.380 49.180 ;
        RECT 5.760 48.750 5.920 48.930 ;
        RECT 6.090 48.750 6.400 48.930 ;
        RECT 6.570 48.750 6.880 48.930 ;
        RECT 7.050 48.750 7.360 48.930 ;
        RECT 7.530 48.920 7.840 48.930 ;
        RECT 8.010 48.920 8.320 48.930 ;
        RECT 7.530 48.750 7.680 48.920 ;
        RECT 8.160 48.750 8.320 48.920 ;
        RECT 8.490 48.750 8.800 48.930 ;
        RECT 8.970 48.750 9.280 48.930 ;
        RECT 9.450 48.750 9.760 48.930 ;
        RECT 9.930 48.750 10.240 48.930 ;
        RECT 10.410 48.750 10.720 48.930 ;
        RECT 10.890 48.750 11.200 48.930 ;
        RECT 11.370 48.750 11.680 48.930 ;
        RECT 11.850 48.750 12.160 48.930 ;
        RECT 12.330 48.750 12.640 48.930 ;
        RECT 12.810 48.750 13.120 48.930 ;
        RECT 13.290 48.750 13.600 48.930 ;
        RECT 13.770 48.750 14.080 48.930 ;
        RECT 14.250 48.750 14.560 48.930 ;
        RECT 14.730 48.750 15.040 48.930 ;
        RECT 15.210 48.750 15.520 48.930 ;
        RECT 15.690 48.750 16.000 48.930 ;
        RECT 16.170 48.750 16.480 48.930 ;
        RECT 16.650 48.750 16.960 48.930 ;
        RECT 17.130 48.750 17.440 48.930 ;
        RECT 17.610 48.750 17.920 48.930 ;
        RECT 18.090 48.750 18.400 48.930 ;
        RECT 18.570 48.750 18.880 48.930 ;
        RECT 19.050 48.750 19.360 48.930 ;
        RECT 19.530 48.750 19.840 48.930 ;
        RECT 20.010 48.750 20.320 48.930 ;
        RECT 20.490 48.750 20.800 48.930 ;
        RECT 20.970 48.750 21.280 48.930 ;
        RECT 21.450 48.750 21.760 48.930 ;
        RECT 21.930 48.750 22.240 48.930 ;
        RECT 22.410 48.750 22.720 48.930 ;
        RECT 22.890 48.750 23.200 48.930 ;
        RECT 23.370 48.750 23.680 48.930 ;
        RECT 23.850 48.750 24.160 48.930 ;
        RECT 24.330 48.750 24.640 48.930 ;
        RECT 24.810 48.750 25.120 48.930 ;
        RECT 25.290 48.750 25.600 48.930 ;
        RECT 25.770 48.750 26.080 48.930 ;
        RECT 26.250 48.750 26.560 48.930 ;
        RECT 26.730 48.750 27.040 48.930 ;
        RECT 27.210 48.750 27.520 48.930 ;
        RECT 27.690 48.750 28.000 48.930 ;
        RECT 28.170 48.750 28.480 48.930 ;
        RECT 28.650 48.750 28.960 48.930 ;
        RECT 29.130 48.750 29.440 48.930 ;
        RECT 29.610 48.750 29.920 48.930 ;
        RECT 30.090 48.750 30.400 48.930 ;
        RECT 30.570 48.750 30.880 48.930 ;
        RECT 31.050 48.750 31.360 48.930 ;
        RECT 31.530 48.750 31.840 48.930 ;
        RECT 32.010 48.750 32.320 48.930 ;
        RECT 32.490 48.750 32.800 48.930 ;
        RECT 32.970 48.750 33.280 48.930 ;
        RECT 33.450 48.750 33.760 48.930 ;
        RECT 33.930 48.750 34.240 48.930 ;
        RECT 34.410 48.750 34.720 48.930 ;
        RECT 34.890 48.750 35.200 48.930 ;
        RECT 35.370 48.750 35.680 48.930 ;
        RECT 35.850 48.750 36.160 48.930 ;
        RECT 36.330 48.750 36.640 48.930 ;
        RECT 36.810 48.750 37.120 48.930 ;
        RECT 37.290 48.750 37.600 48.930 ;
        RECT 37.770 48.750 38.080 48.930 ;
        RECT 38.250 48.750 38.560 48.930 ;
        RECT 38.730 48.750 39.040 48.930 ;
        RECT 39.210 48.750 39.520 48.930 ;
        RECT 39.690 48.750 40.000 48.930 ;
        RECT 40.170 48.750 40.480 48.930 ;
        RECT 40.650 48.750 40.960 48.930 ;
        RECT 41.130 48.750 41.440 48.930 ;
        RECT 41.610 48.750 41.920 48.930 ;
        RECT 42.090 48.750 42.400 48.930 ;
        RECT 42.570 48.750 42.880 48.930 ;
        RECT 43.050 48.750 43.360 48.930 ;
        RECT 43.530 48.750 43.840 48.930 ;
        RECT 44.010 48.750 44.320 48.930 ;
        RECT 44.490 48.750 44.800 48.930 ;
        RECT 44.970 48.750 45.280 48.930 ;
        RECT 45.450 48.750 45.760 48.930 ;
        RECT 45.930 48.750 46.240 48.930 ;
        RECT 46.410 48.750 46.720 48.930 ;
        RECT 46.890 48.750 47.200 48.930 ;
        RECT 47.370 48.920 47.680 48.930 ;
        RECT 47.850 48.920 48.160 48.930 ;
        RECT 47.370 48.750 47.520 48.920 ;
        RECT 48.000 48.750 48.160 48.920 ;
        RECT 48.330 48.750 48.640 48.930 ;
        RECT 48.810 48.750 49.120 48.930 ;
        RECT 49.290 48.750 49.600 48.930 ;
        RECT 49.770 48.750 50.080 48.930 ;
        RECT 50.250 48.920 50.400 48.930 ;
        RECT 50.880 48.920 51.040 48.930 ;
        RECT 50.250 48.750 50.560 48.920 ;
        RECT 50.730 48.750 51.040 48.920 ;
        RECT 51.210 48.750 51.520 48.930 ;
        RECT 51.690 48.750 52.000 48.930 ;
        RECT 52.170 48.750 52.480 48.930 ;
        RECT 52.650 48.750 52.960 48.930 ;
        RECT 53.130 48.750 53.440 48.930 ;
        RECT 53.610 48.750 53.920 48.930 ;
        RECT 54.090 48.750 54.400 48.930 ;
        RECT 54.570 48.750 54.880 48.930 ;
        RECT 55.050 48.750 55.360 48.930 ;
        RECT 55.530 48.750 55.840 48.930 ;
        RECT 56.010 48.750 56.320 48.930 ;
        RECT 56.490 48.750 56.800 48.930 ;
        RECT 56.970 48.750 57.280 48.930 ;
        RECT 57.450 48.750 57.760 48.930 ;
        RECT 57.930 48.750 58.240 48.930 ;
        RECT 58.410 48.750 58.720 48.930 ;
        RECT 58.890 48.750 59.200 48.930 ;
        RECT 59.370 48.750 59.680 48.930 ;
        RECT 59.850 48.750 60.160 48.930 ;
        RECT 60.330 48.750 60.640 48.930 ;
        RECT 60.810 48.750 61.120 48.930 ;
        RECT 61.290 48.750 61.600 48.930 ;
        RECT 61.770 48.750 62.080 48.930 ;
        RECT 62.250 48.750 62.560 48.930 ;
        RECT 62.730 48.750 63.040 48.930 ;
        RECT 63.210 48.750 63.520 48.930 ;
        RECT 63.690 48.750 64.000 48.930 ;
        RECT 64.170 48.750 64.480 48.930 ;
        RECT 64.650 48.750 64.960 48.930 ;
        RECT 65.130 48.750 65.440 48.930 ;
        RECT 65.610 48.750 65.920 48.930 ;
        RECT 66.090 48.750 66.400 48.930 ;
        RECT 66.570 48.750 66.880 48.930 ;
        RECT 67.050 48.750 67.360 48.930 ;
        RECT 67.530 48.750 67.840 48.930 ;
        RECT 68.010 48.750 68.320 48.930 ;
        RECT 68.490 48.750 68.800 48.930 ;
        RECT 68.970 48.750 69.280 48.930 ;
        RECT 69.450 48.750 69.760 48.930 ;
        RECT 69.930 48.750 70.240 48.930 ;
        RECT 70.410 48.750 70.720 48.930 ;
        RECT 70.890 48.750 71.200 48.930 ;
        RECT 71.370 48.750 71.680 48.930 ;
        RECT 71.850 48.750 72.160 48.930 ;
        RECT 72.330 48.750 72.640 48.930 ;
        RECT 72.810 48.750 73.120 48.930 ;
        RECT 73.290 48.750 73.600 48.930 ;
        RECT 73.770 48.750 74.080 48.930 ;
        RECT 74.250 48.750 74.560 48.930 ;
        RECT 74.730 48.750 75.040 48.930 ;
        RECT 75.210 48.750 75.520 48.930 ;
        RECT 75.690 48.750 76.000 48.930 ;
        RECT 76.170 48.750 76.480 48.930 ;
        RECT 76.650 48.750 76.960 48.930 ;
        RECT 77.130 48.750 77.440 48.930 ;
        RECT 77.610 48.750 77.920 48.930 ;
        RECT 78.090 48.750 78.400 48.930 ;
        RECT 78.570 48.750 78.880 48.930 ;
        RECT 79.050 48.750 79.360 48.930 ;
        RECT 79.530 48.750 79.840 48.930 ;
        RECT 80.010 48.750 80.320 48.930 ;
        RECT 80.490 48.750 80.800 48.930 ;
        RECT 80.970 48.920 81.280 48.930 ;
        RECT 81.450 48.920 81.760 48.930 ;
        RECT 80.970 48.750 81.120 48.920 ;
        RECT 81.600 48.750 81.760 48.920 ;
        RECT 81.930 48.750 82.240 48.930 ;
        RECT 82.410 48.750 82.720 48.930 ;
        RECT 82.890 48.750 83.200 48.930 ;
        RECT 83.370 48.750 83.680 48.930 ;
        RECT 83.850 48.750 84.160 48.930 ;
        RECT 84.330 48.750 84.640 48.930 ;
        RECT 84.810 48.750 85.120 48.930 ;
        RECT 85.290 48.750 85.600 48.930 ;
        RECT 85.770 48.750 86.080 48.930 ;
        RECT 86.250 48.750 86.560 48.930 ;
        RECT 86.730 48.750 87.040 48.930 ;
        RECT 87.210 48.750 87.520 48.930 ;
        RECT 87.690 48.750 88.000 48.930 ;
        RECT 88.170 48.750 88.480 48.930 ;
        RECT 88.650 48.750 88.960 48.930 ;
        RECT 89.130 48.750 89.440 48.930 ;
        RECT 89.610 48.750 89.920 48.930 ;
        RECT 90.090 48.750 90.400 48.930 ;
        RECT 90.570 48.750 90.880 48.930 ;
        RECT 91.050 48.750 91.360 48.930 ;
        RECT 91.530 48.750 91.840 48.930 ;
        RECT 92.010 48.750 92.320 48.930 ;
        RECT 92.490 48.750 92.800 48.930 ;
        RECT 92.970 48.750 93.280 48.930 ;
        RECT 93.450 48.750 93.760 48.930 ;
        RECT 93.930 48.750 94.240 48.930 ;
        RECT 94.410 48.920 94.560 48.930 ;
        RECT 95.040 48.920 95.200 48.930 ;
        RECT 94.410 48.750 94.720 48.920 ;
        RECT 94.890 48.750 95.200 48.920 ;
        RECT 95.370 48.750 95.680 48.930 ;
        RECT 95.850 48.750 96.160 48.930 ;
        RECT 96.330 48.750 96.640 48.930 ;
        RECT 96.810 48.750 97.120 48.930 ;
        RECT 97.290 48.750 97.600 48.930 ;
        RECT 97.770 48.750 98.080 48.930 ;
        RECT 98.250 48.750 98.560 48.930 ;
        RECT 98.730 48.750 99.040 48.930 ;
        RECT 99.210 48.750 99.520 48.930 ;
        RECT 99.690 48.750 100.000 48.930 ;
        RECT 100.170 48.750 100.480 48.930 ;
        RECT 100.650 48.750 100.960 48.930 ;
        RECT 101.130 48.750 101.440 48.930 ;
        RECT 101.610 48.750 101.920 48.930 ;
        RECT 102.090 48.750 102.400 48.930 ;
        RECT 102.570 48.750 102.880 48.930 ;
        RECT 103.050 48.750 103.360 48.930 ;
        RECT 103.530 48.750 103.840 48.930 ;
        RECT 104.010 48.750 104.320 48.930 ;
        RECT 104.490 48.750 104.800 48.930 ;
        RECT 104.970 48.750 105.280 48.930 ;
        RECT 105.450 48.750 105.760 48.930 ;
        RECT 105.930 48.750 106.240 48.930 ;
        RECT 106.410 48.750 106.720 48.930 ;
        RECT 106.890 48.920 107.200 48.930 ;
        RECT 107.370 48.920 107.680 48.930 ;
        RECT 106.890 48.750 107.040 48.920 ;
        RECT 107.520 48.750 107.680 48.920 ;
        RECT 107.850 48.920 108.000 48.930 ;
        RECT 108.480 48.920 108.640 48.930 ;
        RECT 107.850 48.750 108.160 48.920 ;
        RECT 108.330 48.750 108.640 48.920 ;
        RECT 108.810 48.750 109.120 48.930 ;
        RECT 109.290 48.750 109.600 48.930 ;
        RECT 109.770 48.750 110.080 48.930 ;
        RECT 110.250 48.750 110.560 48.930 ;
        RECT 110.730 48.750 111.040 48.930 ;
        RECT 111.210 48.750 111.520 48.930 ;
        RECT 111.690 48.750 112.000 48.930 ;
        RECT 112.170 48.750 112.480 48.930 ;
        RECT 112.650 48.750 112.960 48.930 ;
        RECT 113.130 48.750 113.440 48.930 ;
        RECT 113.610 48.750 113.920 48.930 ;
        RECT 114.090 48.750 114.400 48.930 ;
        RECT 114.570 48.750 114.880 48.930 ;
        RECT 115.050 48.750 115.360 48.930 ;
        RECT 115.530 48.750 115.840 48.930 ;
        RECT 116.010 48.750 116.320 48.930 ;
        RECT 116.490 48.750 116.800 48.930 ;
        RECT 116.970 48.750 117.280 48.930 ;
        RECT 117.450 48.750 117.760 48.930 ;
        RECT 117.930 48.750 118.240 48.930 ;
        RECT 118.410 48.750 118.720 48.930 ;
        RECT 118.890 48.750 119.200 48.930 ;
        RECT 119.370 48.750 119.680 48.930 ;
        RECT 119.850 48.750 120.160 48.930 ;
        RECT 120.330 48.750 120.640 48.930 ;
        RECT 120.810 48.750 121.120 48.930 ;
        RECT 121.290 48.750 121.600 48.930 ;
        RECT 121.770 48.750 122.080 48.930 ;
        RECT 122.250 48.750 122.560 48.930 ;
        RECT 122.730 48.920 123.040 48.930 ;
        RECT 123.210 48.920 123.520 48.930 ;
        RECT 122.730 48.750 122.880 48.920 ;
        RECT 123.360 48.750 123.520 48.920 ;
        RECT 123.690 48.750 124.000 48.930 ;
        RECT 124.170 48.750 124.480 48.930 ;
        RECT 124.650 48.750 124.960 48.930 ;
        RECT 125.130 48.750 125.440 48.930 ;
        RECT 125.610 48.750 125.920 48.930 ;
        RECT 126.090 48.750 126.400 48.930 ;
        RECT 126.570 48.750 126.880 48.930 ;
        RECT 127.050 48.750 127.360 48.930 ;
        RECT 127.530 48.750 127.840 48.930 ;
        RECT 128.010 48.750 128.320 48.930 ;
        RECT 128.490 48.750 128.800 48.930 ;
        RECT 128.970 48.750 129.280 48.930 ;
        RECT 129.450 48.750 129.760 48.930 ;
        RECT 129.930 48.750 130.240 48.930 ;
        RECT 130.410 48.750 130.720 48.930 ;
        RECT 130.890 48.750 131.200 48.930 ;
        RECT 131.370 48.750 131.680 48.930 ;
        RECT 131.850 48.750 132.160 48.930 ;
        RECT 132.330 48.750 132.640 48.930 ;
        RECT 132.810 48.750 133.120 48.930 ;
        RECT 133.290 48.750 133.600 48.930 ;
        RECT 133.770 48.750 134.080 48.930 ;
        RECT 134.250 48.750 134.560 48.930 ;
        RECT 134.730 48.750 135.040 48.930 ;
        RECT 135.210 48.750 135.520 48.930 ;
        RECT 135.690 48.750 136.000 48.930 ;
        RECT 136.170 48.750 136.480 48.930 ;
        RECT 136.650 48.750 136.960 48.930 ;
        RECT 137.130 48.750 137.440 48.930 ;
        RECT 137.610 48.750 137.920 48.930 ;
        RECT 138.090 48.750 138.400 48.930 ;
        RECT 138.570 48.750 138.880 48.930 ;
        RECT 139.050 48.750 139.360 48.930 ;
        RECT 139.530 48.750 139.840 48.930 ;
        RECT 140.010 48.750 140.320 48.930 ;
        RECT 140.490 48.750 140.800 48.930 ;
        RECT 140.970 48.750 141.280 48.930 ;
        RECT 141.450 48.920 141.760 48.930 ;
        RECT 141.930 48.920 142.080 48.930 ;
        RECT 141.450 48.750 141.600 48.920 ;
        RECT 6.260 48.500 9.000 48.520 ;
        RECT 6.260 48.330 6.470 48.500 ;
        RECT 6.640 48.330 6.910 48.500 ;
        RECT 7.080 48.330 7.320 48.500 ;
        RECT 7.490 48.330 7.750 48.500 ;
        RECT 7.920 48.330 8.190 48.500 ;
        RECT 8.360 48.330 8.600 48.500 ;
        RECT 8.770 48.330 9.000 48.500 ;
        RECT 6.260 47.450 9.000 48.330 ;
        RECT 10.230 48.450 10.820 48.480 ;
        RECT 10.230 48.280 10.260 48.450 ;
        RECT 10.430 48.280 10.620 48.450 ;
        RECT 10.790 48.280 10.820 48.450 ;
        RECT 6.500 46.130 6.830 46.800 ;
        RECT 7.230 46.470 7.560 47.450 ;
        RECT 7.780 46.130 8.110 46.800 ;
        RECT 8.510 46.470 8.840 47.450 ;
        RECT 9.710 47.300 10.040 48.230 ;
        RECT 10.230 47.500 10.820 48.280 ;
        RECT 11.000 48.410 12.440 48.580 ;
        RECT 11.000 47.300 11.170 48.410 ;
        RECT 9.710 47.130 11.170 47.300 ;
        RECT 6.340 45.130 9.070 46.130 ;
        RECT 9.710 45.270 9.980 47.130 ;
        RECT 10.840 46.630 11.170 47.130 ;
        RECT 11.350 46.920 11.600 48.230 ;
        RECT 11.840 47.610 12.090 48.230 ;
        RECT 12.270 47.960 12.440 48.410 ;
        RECT 12.620 48.450 12.950 48.480 ;
        RECT 12.620 48.280 12.650 48.450 ;
        RECT 12.820 48.280 12.950 48.450 ;
        RECT 12.620 48.140 12.950 48.280 ;
        RECT 13.130 48.410 14.870 48.580 ;
        RECT 13.130 47.960 13.300 48.410 ;
        RECT 12.270 47.790 13.300 47.960 ;
        RECT 13.480 47.610 13.650 48.230 ;
        RECT 14.180 47.970 14.510 48.230 ;
        RECT 11.840 47.440 13.650 47.610 ;
        RECT 13.830 47.440 14.050 47.770 ;
        RECT 13.480 47.260 13.650 47.440 ;
        RECT 11.350 46.690 11.880 46.920 ;
        RECT 11.350 45.770 11.620 46.690 ;
      LAYER li1 ;
        RECT 12.300 46.390 12.840 47.260 ;
      LAYER li1 ;
        RECT 13.480 47.090 13.700 47.260 ;
        RECT 10.160 45.140 11.110 45.770 ;
        RECT 11.290 45.270 11.620 45.770 ;
        RECT 11.800 45.140 12.390 46.020 ;
      LAYER li1 ;
        RECT 12.670 45.400 12.840 46.390 ;
        RECT 13.020 45.580 13.350 46.880 ;
      LAYER li1 ;
        RECT 13.530 46.100 13.700 47.090 ;
        RECT 13.880 46.920 14.050 47.440 ;
        RECT 14.230 47.270 14.400 47.970 ;
        RECT 14.700 47.820 14.870 48.410 ;
        RECT 15.050 48.450 16.000 48.480 ;
        RECT 15.050 48.280 15.080 48.450 ;
        RECT 15.250 48.280 15.440 48.450 ;
        RECT 15.610 48.280 15.800 48.450 ;
        RECT 15.970 48.280 16.000 48.450 ;
        RECT 15.050 48.000 16.000 48.280 ;
        RECT 16.180 48.410 17.210 48.580 ;
        RECT 16.180 47.820 16.350 48.410 ;
        RECT 14.700 47.770 16.350 47.820 ;
        RECT 14.580 47.650 16.350 47.770 ;
        RECT 14.580 47.450 14.910 47.650 ;
        RECT 16.530 47.470 16.860 48.230 ;
        RECT 17.040 48.050 17.210 48.410 ;
        RECT 17.390 48.450 18.340 48.530 ;
        RECT 17.390 48.280 17.420 48.450 ;
        RECT 17.590 48.280 17.780 48.450 ;
        RECT 17.950 48.280 18.140 48.450 ;
        RECT 18.310 48.280 18.340 48.450 ;
        RECT 17.390 48.230 18.340 48.280 ;
        RECT 17.040 47.880 18.850 48.050 ;
        RECT 15.090 47.300 16.860 47.470 ;
        RECT 15.090 47.270 15.260 47.300 ;
        RECT 14.230 47.100 15.260 47.270 ;
        RECT 18.170 47.120 18.500 47.700 ;
        RECT 13.880 46.690 14.910 46.920 ;
        RECT 14.580 46.200 14.910 46.690 ;
        RECT 15.090 46.420 15.260 47.100 ;
        RECT 15.440 46.950 18.500 47.120 ;
        RECT 15.440 46.600 15.770 46.950 ;
      LAYER li1 ;
        RECT 16.210 46.600 18.060 46.770 ;
      LAYER li1 ;
        RECT 15.090 46.250 17.710 46.420 ;
        RECT 13.530 45.600 13.800 46.100 ;
        RECT 15.090 46.020 15.260 46.250 ;
      LAYER li1 ;
        RECT 17.890 46.070 18.060 46.600 ;
      LAYER li1 ;
        RECT 14.250 45.850 15.260 46.020 ;
      LAYER li1 ;
        RECT 15.440 45.900 18.060 46.070 ;
      LAYER li1 ;
        RECT 14.250 45.600 14.580 45.850 ;
      LAYER li1 ;
        RECT 15.440 45.400 15.610 45.900 ;
        RECT 12.670 45.230 15.610 45.400 ;
      LAYER li1 ;
        RECT 16.760 45.140 17.710 45.720 ;
      LAYER li1 ;
        RECT 17.890 45.210 18.060 45.900 ;
      LAYER li1 ;
        RECT 18.240 46.100 18.500 46.950 ;
        RECT 18.680 46.530 18.850 47.880 ;
        RECT 19.030 47.620 19.280 48.530 ;
        RECT 20.090 48.450 21.040 48.480 ;
        RECT 21.870 48.450 22.770 48.480 ;
        RECT 20.090 48.280 20.120 48.450 ;
        RECT 20.290 48.280 20.480 48.450 ;
        RECT 20.650 48.280 20.840 48.450 ;
        RECT 21.010 48.280 21.040 48.450 ;
        RECT 22.040 48.280 22.230 48.450 ;
        RECT 22.400 48.280 22.590 48.450 ;
        RECT 22.760 48.280 22.770 48.450 ;
        RECT 19.030 47.450 19.910 47.620 ;
        RECT 20.090 47.450 21.040 48.280 ;
        RECT 21.440 47.480 21.690 47.950 ;
        RECT 21.870 47.660 22.770 48.280 ;
        RECT 23.380 48.450 24.320 48.510 ;
        RECT 23.380 48.280 23.400 48.450 ;
        RECT 23.570 48.280 23.760 48.450 ;
        RECT 23.930 48.280 24.120 48.450 ;
        RECT 24.290 48.280 24.320 48.450 ;
        RECT 19.230 46.710 19.560 47.210 ;
        RECT 19.740 47.130 19.910 47.450 ;
        RECT 21.440 47.310 22.450 47.480 ;
        RECT 19.740 46.960 22.100 47.130 ;
        RECT 18.680 46.360 19.850 46.530 ;
        RECT 18.240 45.390 18.570 46.100 ;
        RECT 19.030 45.560 19.360 46.100 ;
        RECT 19.570 45.860 19.850 46.360 ;
        RECT 20.030 45.560 20.200 46.960 ;
        RECT 22.280 46.780 22.450 47.310 ;
        RECT 20.410 46.610 22.450 46.780 ;
        RECT 20.410 46.220 20.740 46.610 ;
      LAYER li1 ;
        RECT 21.060 46.040 21.390 46.430 ;
      LAYER li1 ;
        RECT 19.030 45.390 20.200 45.560 ;
      LAYER li1 ;
        RECT 20.380 45.870 21.390 46.040 ;
        RECT 20.380 45.210 20.550 45.870 ;
      LAYER li1 ;
        RECT 22.220 45.770 22.450 46.610 ;
        RECT 22.950 46.780 23.200 47.780 ;
        RECT 23.380 46.970 24.320 48.280 ;
        RECT 22.950 46.450 24.320 46.780 ;
        RECT 22.950 46.270 23.160 46.450 ;
        RECT 22.830 45.770 23.160 46.270 ;
      LAYER li1 ;
        RECT 17.890 45.040 20.550 45.210 ;
      LAYER li1 ;
        RECT 20.730 45.140 21.680 45.690 ;
        RECT 22.220 45.270 22.550 45.770 ;
        RECT 23.340 45.140 24.290 46.270 ;
      LAYER li1 ;
        RECT 24.500 45.440 24.840 48.510 ;
      LAYER li1 ;
        RECT 25.210 48.500 26.660 48.530 ;
        RECT 25.210 48.330 25.460 48.500 ;
        RECT 25.630 48.330 25.820 48.500 ;
        RECT 25.990 48.330 26.260 48.500 ;
        RECT 26.430 48.330 26.660 48.500 ;
        RECT 25.210 47.460 26.660 48.330 ;
        RECT 25.440 46.020 25.770 46.800 ;
        RECT 25.980 46.470 26.310 47.460 ;
        RECT 25.440 45.620 26.740 46.020 ;
        RECT 25.130 45.140 26.740 45.620 ;
      LAYER li1 ;
        RECT 27.010 45.270 27.260 48.530 ;
      LAYER li1 ;
        RECT 27.440 48.450 30.130 48.530 ;
        RECT 27.610 48.280 27.800 48.450 ;
        RECT 27.970 48.280 28.160 48.450 ;
        RECT 28.330 48.280 28.520 48.450 ;
        RECT 28.690 48.280 28.880 48.450 ;
        RECT 29.050 48.280 29.240 48.450 ;
        RECT 29.410 48.280 29.600 48.450 ;
        RECT 29.770 48.280 29.960 48.450 ;
        RECT 27.440 47.420 30.130 48.280 ;
        RECT 30.310 47.240 30.560 48.530 ;
        RECT 27.470 47.070 30.560 47.240 ;
        RECT 27.470 46.370 27.800 47.070 ;
        RECT 30.310 46.950 30.560 47.070 ;
        RECT 30.740 48.450 32.050 48.510 ;
        RECT 30.740 48.280 30.770 48.450 ;
        RECT 30.940 48.280 31.130 48.450 ;
        RECT 31.300 48.280 31.490 48.450 ;
        RECT 31.660 48.280 31.850 48.450 ;
        RECT 32.020 48.280 32.050 48.450 ;
        RECT 30.740 46.970 32.050 48.280 ;
        RECT 32.410 48.500 33.860 48.530 ;
        RECT 32.410 48.330 32.660 48.500 ;
        RECT 32.830 48.330 33.020 48.500 ;
        RECT 33.190 48.330 33.460 48.500 ;
        RECT 33.630 48.330 33.860 48.500 ;
        RECT 32.410 47.460 33.860 48.330 ;
        RECT 34.170 48.450 35.840 48.530 ;
        RECT 34.170 48.280 34.200 48.450 ;
        RECT 34.370 48.280 34.560 48.450 ;
        RECT 34.730 48.280 34.920 48.450 ;
        RECT 35.090 48.280 35.280 48.450 ;
        RECT 35.450 48.280 35.640 48.450 ;
        RECT 35.810 48.280 35.840 48.450 ;
      LAYER li1 ;
        RECT 28.470 46.830 28.640 46.890 ;
        RECT 28.300 46.550 29.030 46.830 ;
      LAYER li1 ;
        RECT 27.470 46.200 28.680 46.370 ;
        RECT 27.440 45.140 28.330 46.020 ;
        RECT 28.510 45.990 28.680 46.200 ;
      LAYER li1 ;
        RECT 28.860 46.340 29.030 46.550 ;
        RECT 29.210 46.520 29.640 46.890 ;
        RECT 29.840 46.350 30.130 46.890 ;
        RECT 30.370 46.350 31.080 46.680 ;
        RECT 28.860 46.170 29.660 46.340 ;
        RECT 31.430 46.170 31.760 46.790 ;
        RECT 29.490 46.000 31.760 46.170 ;
      LAYER li1 ;
        RECT 32.640 46.020 32.970 46.800 ;
        RECT 33.180 46.470 33.510 47.460 ;
        RECT 34.170 47.070 35.840 48.280 ;
      LAYER li1 ;
        RECT 34.210 46.300 34.510 46.890 ;
        RECT 34.690 46.550 35.880 46.890 ;
        RECT 36.060 46.550 36.390 48.030 ;
        RECT 36.570 46.370 36.840 48.530 ;
      LAYER li1 ;
        RECT 37.690 48.500 39.140 48.530 ;
        RECT 37.690 48.330 37.940 48.500 ;
        RECT 38.110 48.330 38.300 48.500 ;
        RECT 38.470 48.330 38.740 48.500 ;
        RECT 38.910 48.330 39.140 48.500 ;
        RECT 37.690 47.460 39.140 48.330 ;
        RECT 39.450 48.450 40.400 48.530 ;
        RECT 39.450 48.280 39.480 48.450 ;
        RECT 39.650 48.280 39.840 48.450 ;
        RECT 40.010 48.280 40.200 48.450 ;
        RECT 40.370 48.280 40.400 48.450 ;
      LAYER li1 ;
        RECT 35.010 46.200 36.840 46.370 ;
      LAYER li1 ;
        RECT 28.510 45.820 29.310 45.990 ;
      LAYER li1 ;
        RECT 29.920 45.980 30.590 46.000 ;
      LAYER li1 ;
        RECT 29.140 45.650 29.740 45.820 ;
        RECT 28.630 45.210 28.960 45.640 ;
        RECT 29.410 45.390 29.740 45.650 ;
        RECT 30.230 45.210 30.560 45.800 ;
        RECT 28.630 45.040 30.560 45.210 ;
        RECT 30.770 45.140 32.070 45.820 ;
        RECT 32.640 45.620 33.940 46.020 ;
        RECT 32.330 45.140 33.940 45.620 ;
        RECT 34.170 45.140 34.760 46.100 ;
      LAYER li1 ;
        RECT 35.010 45.270 35.260 46.200 ;
      LAYER li1 ;
        RECT 35.440 45.140 36.390 46.020 ;
      LAYER li1 ;
        RECT 36.570 45.270 36.840 46.200 ;
      LAYER li1 ;
        RECT 37.920 46.020 38.250 46.800 ;
        RECT 38.460 46.470 38.790 47.460 ;
        RECT 39.450 46.950 40.400 48.280 ;
      LAYER li1 ;
        RECT 40.580 46.850 40.830 48.530 ;
      LAYER li1 ;
        RECT 41.010 48.450 41.960 48.530 ;
        RECT 41.010 48.280 41.040 48.450 ;
        RECT 41.210 48.280 41.400 48.450 ;
        RECT 41.570 48.280 41.760 48.450 ;
        RECT 41.930 48.280 41.960 48.450 ;
        RECT 41.010 47.030 41.960 48.280 ;
      LAYER li1 ;
        RECT 42.140 46.850 42.470 48.530 ;
      LAYER li1 ;
        RECT 42.650 48.450 43.600 48.530 ;
        RECT 42.650 48.280 42.680 48.450 ;
        RECT 42.850 48.280 43.040 48.450 ;
        RECT 43.210 48.280 43.400 48.450 ;
        RECT 43.570 48.280 43.600 48.450 ;
        RECT 42.650 47.070 43.600 48.280 ;
      LAYER li1 ;
        RECT 40.580 46.680 42.470 46.850 ;
        RECT 40.580 46.550 40.750 46.680 ;
        RECT 43.250 46.550 43.580 46.890 ;
        RECT 39.490 46.320 40.750 46.550 ;
      LAYER li1 ;
        RECT 40.930 46.370 42.960 46.500 ;
        RECT 43.780 46.370 44.030 48.530 ;
        RECT 44.410 48.500 45.860 48.530 ;
        RECT 44.410 48.330 44.660 48.500 ;
        RECT 44.830 48.330 45.020 48.500 ;
        RECT 45.190 48.330 45.460 48.500 ;
        RECT 45.630 48.330 45.860 48.500 ;
        RECT 44.410 47.460 45.860 48.330 ;
        RECT 46.170 48.450 47.120 48.530 ;
        RECT 46.170 48.280 46.200 48.450 ;
        RECT 46.370 48.280 46.560 48.450 ;
        RECT 46.730 48.280 46.920 48.450 ;
        RECT 47.090 48.280 47.120 48.450 ;
        RECT 40.930 46.330 44.030 46.370 ;
      LAYER li1 ;
        RECT 40.580 46.150 40.750 46.320 ;
      LAYER li1 ;
        RECT 42.790 46.200 44.030 46.330 ;
        RECT 37.920 45.620 39.220 46.020 ;
        RECT 37.610 45.140 39.220 45.620 ;
        RECT 39.450 45.140 40.400 46.100 ;
      LAYER li1 ;
        RECT 40.580 45.980 42.390 46.150 ;
        RECT 40.580 45.270 40.830 45.980 ;
      LAYER li1 ;
        RECT 41.010 45.140 41.960 45.800 ;
      LAYER li1 ;
        RECT 42.140 45.270 42.390 45.980 ;
      LAYER li1 ;
        RECT 42.570 45.140 43.520 46.020 ;
        RECT 43.700 45.270 44.030 46.200 ;
        RECT 44.640 46.020 44.970 46.800 ;
        RECT 45.180 46.470 45.510 47.460 ;
        RECT 46.170 46.950 47.120 48.280 ;
      LAYER li1 ;
        RECT 46.210 46.320 47.100 46.710 ;
        RECT 47.300 46.470 47.550 48.530 ;
      LAYER li1 ;
        RECT 47.740 48.450 48.330 48.530 ;
        RECT 47.740 48.280 47.770 48.450 ;
        RECT 47.940 48.280 48.130 48.450 ;
        RECT 48.300 48.280 48.330 48.450 ;
        RECT 47.740 46.950 48.330 48.280 ;
        RECT 48.730 48.500 50.180 48.530 ;
        RECT 48.730 48.330 48.980 48.500 ;
        RECT 49.150 48.330 49.340 48.500 ;
        RECT 49.510 48.330 49.780 48.500 ;
        RECT 49.950 48.330 50.180 48.500 ;
        RECT 48.730 47.460 50.180 48.330 ;
        RECT 50.970 48.450 51.920 48.530 ;
        RECT 50.970 48.280 51.000 48.450 ;
        RECT 51.170 48.280 51.360 48.450 ;
        RECT 51.530 48.280 51.720 48.450 ;
        RECT 51.890 48.280 51.920 48.450 ;
      LAYER li1 ;
        RECT 47.300 46.300 47.880 46.470 ;
        RECT 48.060 46.300 48.360 46.630 ;
        RECT 47.660 46.120 47.880 46.300 ;
      LAYER li1 ;
        RECT 44.640 45.620 45.940 46.020 ;
        RECT 44.330 45.140 45.940 45.620 ;
        RECT 46.170 45.140 47.480 46.120 ;
      LAYER li1 ;
        RECT 47.660 45.950 48.260 46.120 ;
        RECT 47.930 45.780 48.260 45.950 ;
      LAYER li1 ;
        RECT 48.960 46.020 49.290 46.800 ;
        RECT 49.500 46.470 49.830 47.460 ;
        RECT 50.970 46.950 51.920 48.280 ;
      LAYER li1 ;
        RECT 52.100 46.850 52.350 48.530 ;
      LAYER li1 ;
        RECT 52.530 48.450 53.480 48.530 ;
        RECT 52.530 48.280 52.560 48.450 ;
        RECT 52.730 48.280 52.920 48.450 ;
        RECT 53.090 48.280 53.280 48.450 ;
        RECT 53.450 48.280 53.480 48.450 ;
        RECT 52.530 47.030 53.480 48.280 ;
      LAYER li1 ;
        RECT 53.660 46.850 53.990 48.530 ;
      LAYER li1 ;
        RECT 54.170 48.450 55.120 48.530 ;
        RECT 54.170 48.280 54.200 48.450 ;
        RECT 54.370 48.280 54.560 48.450 ;
        RECT 54.730 48.280 54.920 48.450 ;
        RECT 55.090 48.280 55.120 48.450 ;
        RECT 54.170 47.070 55.120 48.280 ;
      LAYER li1 ;
        RECT 52.100 46.680 53.990 46.850 ;
        RECT 52.100 46.550 52.270 46.680 ;
        RECT 54.770 46.550 55.100 46.890 ;
        RECT 51.010 46.320 52.270 46.550 ;
      LAYER li1 ;
        RECT 52.450 46.370 54.480 46.500 ;
        RECT 55.300 46.370 55.550 48.530 ;
        RECT 55.930 48.500 57.380 48.530 ;
        RECT 55.930 48.330 56.180 48.500 ;
        RECT 56.350 48.330 56.540 48.500 ;
        RECT 56.710 48.330 56.980 48.500 ;
        RECT 57.150 48.330 57.380 48.500 ;
        RECT 55.930 47.460 57.380 48.330 ;
        RECT 57.690 48.450 58.640 48.530 ;
        RECT 57.690 48.280 57.720 48.450 ;
        RECT 57.890 48.280 58.080 48.450 ;
        RECT 58.250 48.280 58.440 48.450 ;
        RECT 58.610 48.280 58.640 48.450 ;
        RECT 52.450 46.330 55.550 46.370 ;
      LAYER li1 ;
        RECT 52.100 46.150 52.270 46.320 ;
      LAYER li1 ;
        RECT 54.310 46.200 55.550 46.330 ;
      LAYER li1 ;
        RECT 47.930 45.610 48.320 45.780 ;
      LAYER li1 ;
        RECT 48.960 45.620 50.260 46.020 ;
      LAYER li1 ;
        RECT 47.930 45.290 48.260 45.610 ;
      LAYER li1 ;
        RECT 48.650 45.140 50.260 45.620 ;
        RECT 50.970 45.140 51.920 46.100 ;
      LAYER li1 ;
        RECT 52.100 45.980 53.910 46.150 ;
        RECT 52.100 45.270 52.350 45.980 ;
      LAYER li1 ;
        RECT 52.530 45.140 53.480 45.800 ;
      LAYER li1 ;
        RECT 53.660 45.270 53.910 45.980 ;
      LAYER li1 ;
        RECT 54.090 45.140 55.040 46.020 ;
        RECT 55.220 45.270 55.550 46.200 ;
        RECT 56.160 46.020 56.490 46.800 ;
        RECT 56.700 46.470 57.030 47.460 ;
        RECT 57.690 46.950 58.640 48.280 ;
      LAYER li1 ;
        RECT 58.820 46.850 59.070 48.530 ;
      LAYER li1 ;
        RECT 59.250 48.450 60.200 48.530 ;
        RECT 59.250 48.280 59.280 48.450 ;
        RECT 59.450 48.280 59.640 48.450 ;
        RECT 59.810 48.280 60.000 48.450 ;
        RECT 60.170 48.280 60.200 48.450 ;
        RECT 59.250 47.030 60.200 48.280 ;
      LAYER li1 ;
        RECT 60.380 46.850 60.710 48.530 ;
      LAYER li1 ;
        RECT 60.890 48.450 61.840 48.530 ;
        RECT 60.890 48.280 60.920 48.450 ;
        RECT 61.090 48.280 61.280 48.450 ;
        RECT 61.450 48.280 61.640 48.450 ;
        RECT 61.810 48.280 61.840 48.450 ;
        RECT 60.890 47.070 61.840 48.280 ;
      LAYER li1 ;
        RECT 58.820 46.680 60.710 46.850 ;
        RECT 58.820 46.550 58.990 46.680 ;
        RECT 61.490 46.550 61.820 46.890 ;
        RECT 57.730 46.320 58.990 46.550 ;
      LAYER li1 ;
        RECT 59.170 46.370 61.200 46.500 ;
        RECT 62.020 46.370 62.270 48.530 ;
        RECT 62.650 48.500 64.100 48.530 ;
        RECT 62.650 48.330 62.900 48.500 ;
        RECT 63.070 48.330 63.260 48.500 ;
        RECT 63.430 48.330 63.700 48.500 ;
        RECT 63.870 48.330 64.100 48.500 ;
        RECT 62.650 47.460 64.100 48.330 ;
        RECT 64.410 48.450 66.080 48.530 ;
        RECT 64.410 48.280 64.440 48.450 ;
        RECT 64.610 48.280 64.800 48.450 ;
        RECT 64.970 48.280 65.160 48.450 ;
        RECT 65.330 48.280 65.520 48.450 ;
        RECT 65.690 48.280 65.880 48.450 ;
        RECT 66.050 48.280 66.080 48.450 ;
        RECT 59.170 46.330 62.270 46.370 ;
      LAYER li1 ;
        RECT 58.820 46.150 58.990 46.320 ;
      LAYER li1 ;
        RECT 61.030 46.200 62.270 46.330 ;
        RECT 56.160 45.620 57.460 46.020 ;
        RECT 55.850 45.140 57.460 45.620 ;
        RECT 57.690 45.140 58.640 46.100 ;
      LAYER li1 ;
        RECT 58.820 45.980 60.630 46.150 ;
        RECT 58.820 45.270 59.070 45.980 ;
      LAYER li1 ;
        RECT 59.250 45.140 60.200 45.800 ;
      LAYER li1 ;
        RECT 60.380 45.270 60.630 45.980 ;
      LAYER li1 ;
        RECT 60.810 45.140 61.760 46.020 ;
        RECT 61.940 45.270 62.270 46.200 ;
        RECT 62.880 46.020 63.210 46.800 ;
        RECT 63.420 46.470 63.750 47.460 ;
        RECT 64.410 47.070 66.080 48.280 ;
      LAYER li1 ;
        RECT 64.450 46.550 65.640 46.890 ;
        RECT 65.820 46.550 66.150 46.890 ;
        RECT 66.340 46.370 66.600 48.530 ;
      LAYER li1 ;
        RECT 66.970 48.500 68.420 48.530 ;
        RECT 66.970 48.330 67.220 48.500 ;
        RECT 67.390 48.330 67.580 48.500 ;
        RECT 67.750 48.330 68.020 48.500 ;
        RECT 68.190 48.330 68.420 48.500 ;
        RECT 66.970 47.460 68.420 48.330 ;
        RECT 69.270 48.450 69.860 48.480 ;
        RECT 69.270 48.280 69.300 48.450 ;
        RECT 69.470 48.280 69.660 48.450 ;
        RECT 69.830 48.280 69.860 48.450 ;
      LAYER li1 ;
        RECT 65.520 46.200 66.600 46.370 ;
      LAYER li1 ;
        RECT 62.880 45.620 64.180 46.020 ;
        RECT 62.570 45.140 64.180 45.620 ;
        RECT 64.410 45.140 65.340 46.100 ;
      LAYER li1 ;
        RECT 65.520 45.270 65.850 46.200 ;
      LAYER li1 ;
        RECT 67.200 46.020 67.530 46.800 ;
        RECT 67.740 46.470 68.070 47.460 ;
        RECT 68.750 47.300 69.080 48.230 ;
        RECT 69.270 47.500 69.860 48.280 ;
        RECT 70.040 48.410 71.480 48.580 ;
        RECT 70.040 47.300 70.210 48.410 ;
        RECT 68.750 47.130 70.210 47.300 ;
        RECT 66.040 45.140 66.630 46.020 ;
        RECT 67.200 45.620 68.500 46.020 ;
        RECT 66.890 45.140 68.500 45.620 ;
        RECT 68.750 45.270 69.020 47.130 ;
        RECT 69.880 46.630 70.210 47.130 ;
        RECT 70.390 46.920 70.640 48.230 ;
        RECT 70.880 47.610 71.130 48.230 ;
        RECT 71.310 47.960 71.480 48.410 ;
        RECT 71.660 48.450 71.990 48.480 ;
        RECT 71.660 48.280 71.690 48.450 ;
        RECT 71.860 48.280 71.990 48.450 ;
        RECT 71.660 48.140 71.990 48.280 ;
        RECT 72.170 48.410 73.910 48.580 ;
        RECT 72.170 47.960 72.340 48.410 ;
        RECT 71.310 47.790 72.340 47.960 ;
        RECT 72.520 47.610 72.690 48.230 ;
        RECT 73.220 47.970 73.550 48.230 ;
        RECT 70.880 47.440 72.690 47.610 ;
        RECT 72.870 47.440 73.090 47.770 ;
        RECT 72.520 47.260 72.690 47.440 ;
        RECT 70.390 46.690 70.920 46.920 ;
        RECT 70.390 45.770 70.660 46.690 ;
      LAYER li1 ;
        RECT 71.340 46.390 71.880 47.260 ;
      LAYER li1 ;
        RECT 72.520 47.090 72.740 47.260 ;
        RECT 69.200 45.140 70.150 45.770 ;
        RECT 70.330 45.270 70.660 45.770 ;
        RECT 70.840 45.140 71.430 46.020 ;
      LAYER li1 ;
        RECT 71.710 45.400 71.880 46.390 ;
        RECT 72.060 45.580 72.390 46.880 ;
      LAYER li1 ;
        RECT 72.570 46.100 72.740 47.090 ;
        RECT 72.920 46.920 73.090 47.440 ;
        RECT 73.270 47.270 73.440 47.970 ;
        RECT 73.740 47.820 73.910 48.410 ;
        RECT 74.090 48.450 75.040 48.480 ;
        RECT 74.090 48.280 74.120 48.450 ;
        RECT 74.290 48.280 74.480 48.450 ;
        RECT 74.650 48.280 74.840 48.450 ;
        RECT 75.010 48.280 75.040 48.450 ;
        RECT 74.090 48.000 75.040 48.280 ;
        RECT 75.220 48.410 76.250 48.580 ;
        RECT 75.220 47.820 75.390 48.410 ;
        RECT 73.740 47.770 75.390 47.820 ;
        RECT 73.620 47.650 75.390 47.770 ;
        RECT 73.620 47.450 73.950 47.650 ;
        RECT 75.570 47.470 75.900 48.230 ;
        RECT 76.080 48.050 76.250 48.410 ;
        RECT 76.430 48.450 77.380 48.530 ;
        RECT 76.430 48.280 76.460 48.450 ;
        RECT 76.630 48.280 76.820 48.450 ;
        RECT 76.990 48.280 77.180 48.450 ;
        RECT 77.350 48.280 77.380 48.450 ;
        RECT 76.430 48.230 77.380 48.280 ;
        RECT 76.080 47.880 77.890 48.050 ;
        RECT 74.130 47.300 75.900 47.470 ;
        RECT 74.130 47.270 74.300 47.300 ;
        RECT 73.270 47.100 74.300 47.270 ;
        RECT 77.210 47.120 77.540 47.700 ;
        RECT 72.920 46.690 73.950 46.920 ;
        RECT 73.620 46.200 73.950 46.690 ;
        RECT 74.130 46.420 74.300 47.100 ;
        RECT 74.480 46.950 77.540 47.120 ;
        RECT 74.480 46.600 74.810 46.950 ;
      LAYER li1 ;
        RECT 75.250 46.600 77.100 46.770 ;
      LAYER li1 ;
        RECT 74.130 46.250 76.750 46.420 ;
        RECT 72.570 45.600 72.840 46.100 ;
        RECT 74.130 46.020 74.300 46.250 ;
      LAYER li1 ;
        RECT 76.930 46.070 77.100 46.600 ;
      LAYER li1 ;
        RECT 73.290 45.850 74.300 46.020 ;
      LAYER li1 ;
        RECT 74.480 45.900 77.100 46.070 ;
      LAYER li1 ;
        RECT 73.290 45.600 73.620 45.850 ;
      LAYER li1 ;
        RECT 74.480 45.400 74.650 45.900 ;
        RECT 71.710 45.230 74.650 45.400 ;
      LAYER li1 ;
        RECT 75.800 45.140 76.750 45.720 ;
      LAYER li1 ;
        RECT 76.930 45.210 77.100 45.900 ;
      LAYER li1 ;
        RECT 77.280 46.100 77.540 46.950 ;
        RECT 77.720 46.530 77.890 47.880 ;
        RECT 78.070 47.620 78.320 48.530 ;
        RECT 79.130 48.450 80.080 48.480 ;
        RECT 80.910 48.450 81.810 48.480 ;
        RECT 79.130 48.280 79.160 48.450 ;
        RECT 79.330 48.280 79.520 48.450 ;
        RECT 79.690 48.280 79.880 48.450 ;
        RECT 80.050 48.280 80.080 48.450 ;
        RECT 81.080 48.280 81.270 48.450 ;
        RECT 81.440 48.280 81.630 48.450 ;
        RECT 81.800 48.280 81.810 48.450 ;
        RECT 78.070 47.450 78.950 47.620 ;
        RECT 79.130 47.450 80.080 48.280 ;
        RECT 80.480 47.480 80.730 47.950 ;
        RECT 80.910 47.660 81.810 48.280 ;
        RECT 82.420 48.450 83.360 48.510 ;
        RECT 82.420 48.280 82.440 48.450 ;
        RECT 82.610 48.280 82.800 48.450 ;
        RECT 82.970 48.280 83.160 48.450 ;
        RECT 83.330 48.280 83.360 48.450 ;
        RECT 78.270 46.710 78.600 47.210 ;
        RECT 78.780 47.130 78.950 47.450 ;
        RECT 80.480 47.310 81.490 47.480 ;
        RECT 78.780 46.960 81.140 47.130 ;
        RECT 77.720 46.360 78.890 46.530 ;
        RECT 77.280 45.390 77.610 46.100 ;
        RECT 78.070 45.560 78.400 46.100 ;
        RECT 78.610 45.860 78.890 46.360 ;
        RECT 79.070 45.560 79.240 46.960 ;
        RECT 81.320 46.780 81.490 47.310 ;
        RECT 79.450 46.610 81.490 46.780 ;
        RECT 79.450 46.220 79.780 46.610 ;
      LAYER li1 ;
        RECT 80.100 46.040 80.430 46.430 ;
      LAYER li1 ;
        RECT 78.070 45.390 79.240 45.560 ;
      LAYER li1 ;
        RECT 79.420 45.870 80.430 46.040 ;
        RECT 79.420 45.210 79.590 45.870 ;
      LAYER li1 ;
        RECT 81.260 45.770 81.490 46.610 ;
        RECT 81.990 46.780 82.240 47.780 ;
        RECT 82.420 46.970 83.360 48.280 ;
        RECT 81.990 46.450 83.360 46.780 ;
        RECT 81.990 46.270 82.200 46.450 ;
        RECT 81.870 45.770 82.200 46.270 ;
      LAYER li1 ;
        RECT 76.930 45.040 79.590 45.210 ;
      LAYER li1 ;
        RECT 79.770 45.140 80.720 45.690 ;
        RECT 81.260 45.270 81.590 45.770 ;
        RECT 82.380 45.140 83.330 46.270 ;
      LAYER li1 ;
        RECT 83.540 45.440 83.880 48.510 ;
      LAYER li1 ;
        RECT 84.250 48.500 85.700 48.530 ;
        RECT 84.250 48.330 84.500 48.500 ;
        RECT 84.670 48.330 84.860 48.500 ;
        RECT 85.030 48.330 85.300 48.500 ;
        RECT 85.470 48.330 85.700 48.500 ;
        RECT 84.250 47.460 85.700 48.330 ;
        RECT 86.010 48.450 86.960 48.530 ;
        RECT 86.010 48.280 86.040 48.450 ;
        RECT 86.210 48.280 86.400 48.450 ;
        RECT 86.570 48.280 86.760 48.450 ;
        RECT 86.930 48.280 86.960 48.450 ;
        RECT 84.480 46.020 84.810 46.800 ;
        RECT 85.020 46.470 85.350 47.460 ;
        RECT 86.010 46.950 86.960 48.280 ;
      LAYER li1 ;
        RECT 87.140 46.850 87.390 48.530 ;
      LAYER li1 ;
        RECT 87.570 48.450 88.520 48.530 ;
        RECT 87.570 48.280 87.600 48.450 ;
        RECT 87.770 48.280 87.960 48.450 ;
        RECT 88.130 48.280 88.320 48.450 ;
        RECT 88.490 48.280 88.520 48.450 ;
        RECT 87.570 47.030 88.520 48.280 ;
      LAYER li1 ;
        RECT 88.700 46.850 89.030 48.530 ;
      LAYER li1 ;
        RECT 89.210 48.450 90.160 48.530 ;
        RECT 89.210 48.280 89.240 48.450 ;
        RECT 89.410 48.280 89.600 48.450 ;
        RECT 89.770 48.280 89.960 48.450 ;
        RECT 90.130 48.280 90.160 48.450 ;
        RECT 89.210 47.070 90.160 48.280 ;
      LAYER li1 ;
        RECT 87.140 46.680 89.030 46.850 ;
        RECT 87.140 46.550 87.310 46.680 ;
        RECT 89.810 46.550 90.140 46.890 ;
        RECT 86.050 46.320 87.310 46.550 ;
      LAYER li1 ;
        RECT 87.490 46.370 89.520 46.500 ;
        RECT 90.340 46.370 90.590 48.530 ;
        RECT 91.220 48.500 93.960 48.520 ;
        RECT 91.220 48.330 91.430 48.500 ;
        RECT 91.600 48.330 91.870 48.500 ;
        RECT 92.040 48.330 92.280 48.500 ;
        RECT 92.450 48.330 92.710 48.500 ;
        RECT 92.880 48.330 93.150 48.500 ;
        RECT 93.320 48.330 93.560 48.500 ;
        RECT 93.730 48.330 93.960 48.500 ;
        RECT 91.220 47.450 93.960 48.330 ;
        RECT 87.490 46.330 90.590 46.370 ;
      LAYER li1 ;
        RECT 87.140 46.150 87.310 46.320 ;
      LAYER li1 ;
        RECT 89.350 46.200 90.590 46.330 ;
        RECT 84.480 45.620 85.780 46.020 ;
        RECT 84.170 45.140 85.780 45.620 ;
        RECT 86.010 45.140 86.960 46.100 ;
      LAYER li1 ;
        RECT 87.140 45.980 88.950 46.150 ;
        RECT 87.140 45.270 87.390 45.980 ;
      LAYER li1 ;
        RECT 87.570 45.140 88.520 45.800 ;
      LAYER li1 ;
        RECT 88.700 45.270 88.950 45.980 ;
      LAYER li1 ;
        RECT 89.130 45.140 90.080 46.020 ;
        RECT 90.260 45.270 90.590 46.200 ;
        RECT 91.460 46.130 91.790 46.800 ;
        RECT 92.190 46.470 92.520 47.450 ;
        RECT 92.740 46.130 93.070 46.800 ;
        RECT 93.470 46.470 93.800 47.450 ;
        RECT 91.300 45.130 94.030 46.130 ;
      LAYER li1 ;
        RECT 95.170 45.270 95.420 48.530 ;
      LAYER li1 ;
        RECT 95.600 48.450 98.290 48.530 ;
        RECT 95.770 48.280 95.960 48.450 ;
        RECT 96.130 48.280 96.320 48.450 ;
        RECT 96.490 48.280 96.680 48.450 ;
        RECT 96.850 48.280 97.040 48.450 ;
        RECT 97.210 48.280 97.400 48.450 ;
        RECT 97.570 48.280 97.760 48.450 ;
        RECT 97.930 48.280 98.120 48.450 ;
        RECT 95.600 47.420 98.290 48.280 ;
        RECT 98.470 47.240 98.720 48.530 ;
        RECT 95.630 47.070 98.720 47.240 ;
        RECT 95.630 46.370 95.960 47.070 ;
        RECT 98.470 46.950 98.720 47.070 ;
        RECT 98.900 48.450 100.210 48.510 ;
        RECT 98.900 48.280 98.930 48.450 ;
        RECT 99.100 48.280 99.290 48.450 ;
        RECT 99.460 48.280 99.650 48.450 ;
        RECT 99.820 48.280 100.010 48.450 ;
        RECT 100.180 48.280 100.210 48.450 ;
        RECT 98.900 46.970 100.210 48.280 ;
        RECT 100.570 48.500 102.020 48.530 ;
        RECT 100.570 48.330 100.820 48.500 ;
        RECT 100.990 48.330 101.180 48.500 ;
        RECT 101.350 48.330 101.620 48.500 ;
        RECT 101.790 48.330 102.020 48.500 ;
        RECT 100.570 47.460 102.020 48.330 ;
        RECT 102.330 48.450 103.590 48.530 ;
        RECT 102.330 48.280 102.340 48.450 ;
        RECT 102.510 48.280 102.700 48.450 ;
        RECT 102.870 48.280 103.060 48.450 ;
        RECT 103.230 48.280 103.420 48.450 ;
      LAYER li1 ;
        RECT 96.630 46.830 96.800 46.890 ;
        RECT 96.460 46.550 97.190 46.830 ;
      LAYER li1 ;
        RECT 95.630 46.200 96.840 46.370 ;
        RECT 95.600 45.140 96.490 46.020 ;
        RECT 96.670 45.990 96.840 46.200 ;
      LAYER li1 ;
        RECT 97.020 46.340 97.190 46.550 ;
        RECT 97.370 46.520 97.800 46.890 ;
        RECT 98.000 46.350 98.290 46.890 ;
        RECT 98.530 46.350 99.240 46.680 ;
        RECT 97.020 46.170 97.820 46.340 ;
        RECT 99.590 46.170 99.920 46.790 ;
        RECT 97.650 46.000 99.920 46.170 ;
      LAYER li1 ;
        RECT 100.800 46.020 101.130 46.800 ;
        RECT 101.340 46.470 101.670 47.460 ;
        RECT 102.330 47.050 103.590 48.280 ;
      LAYER li1 ;
        RECT 104.120 48.030 104.290 48.530 ;
        RECT 103.770 46.950 104.290 48.030 ;
      LAYER li1 ;
        RECT 104.550 48.450 105.860 48.530 ;
        RECT 104.550 48.280 104.580 48.450 ;
        RECT 104.750 48.280 104.940 48.450 ;
        RECT 105.110 48.280 105.300 48.450 ;
        RECT 105.470 48.280 105.660 48.450 ;
        RECT 105.830 48.280 105.860 48.450 ;
        RECT 104.550 47.070 105.860 48.280 ;
        RECT 106.330 48.500 107.780 48.530 ;
        RECT 106.330 48.330 106.580 48.500 ;
        RECT 106.750 48.330 106.940 48.500 ;
        RECT 107.110 48.330 107.380 48.500 ;
        RECT 107.550 48.330 107.780 48.500 ;
        RECT 106.330 47.460 107.780 48.330 ;
        RECT 108.570 48.450 109.520 48.530 ;
        RECT 108.570 48.280 108.600 48.450 ;
        RECT 108.770 48.280 108.960 48.450 ;
        RECT 109.130 48.280 109.320 48.450 ;
        RECT 109.490 48.280 109.520 48.450 ;
      LAYER li1 ;
        RECT 103.770 46.870 104.040 46.950 ;
        RECT 102.980 46.700 104.040 46.870 ;
        RECT 102.370 46.310 102.790 46.640 ;
        RECT 102.980 46.130 103.150 46.700 ;
        RECT 104.490 46.580 105.000 46.890 ;
        RECT 105.250 46.580 105.960 46.890 ;
        RECT 103.330 46.310 103.840 46.520 ;
      LAYER li1 ;
        RECT 104.040 46.230 105.910 46.400 ;
        RECT 96.670 45.820 97.470 45.990 ;
      LAYER li1 ;
        RECT 98.080 45.980 98.750 46.000 ;
      LAYER li1 ;
        RECT 97.300 45.650 97.900 45.820 ;
        RECT 96.790 45.210 97.120 45.640 ;
        RECT 97.570 45.390 97.900 45.650 ;
        RECT 98.390 45.210 98.720 45.800 ;
        RECT 96.790 45.040 98.720 45.210 ;
        RECT 98.930 45.140 100.230 45.820 ;
        RECT 100.800 45.620 102.100 46.020 ;
        RECT 100.490 45.140 102.100 45.620 ;
        RECT 102.400 45.210 102.730 46.130 ;
      LAYER li1 ;
        RECT 102.980 45.780 103.510 46.130 ;
        RECT 102.980 45.610 103.520 45.780 ;
        RECT 102.980 45.390 103.510 45.610 ;
      LAYER li1 ;
        RECT 104.040 45.210 104.210 46.230 ;
        RECT 102.400 45.040 104.210 45.210 ;
        RECT 104.390 45.140 105.490 46.050 ;
        RECT 105.660 45.300 105.910 46.230 ;
        RECT 106.560 46.020 106.890 46.800 ;
        RECT 107.100 46.470 107.430 47.460 ;
        RECT 108.570 46.950 109.520 48.280 ;
      LAYER li1 ;
        RECT 109.700 46.850 109.950 48.530 ;
      LAYER li1 ;
        RECT 110.130 48.450 111.080 48.530 ;
        RECT 110.130 48.280 110.160 48.450 ;
        RECT 110.330 48.280 110.520 48.450 ;
        RECT 110.690 48.280 110.880 48.450 ;
        RECT 111.050 48.280 111.080 48.450 ;
        RECT 110.130 47.030 111.080 48.280 ;
      LAYER li1 ;
        RECT 111.260 46.850 111.590 48.530 ;
      LAYER li1 ;
        RECT 111.770 48.450 112.720 48.530 ;
        RECT 111.770 48.280 111.800 48.450 ;
        RECT 111.970 48.280 112.160 48.450 ;
        RECT 112.330 48.280 112.520 48.450 ;
        RECT 112.690 48.280 112.720 48.450 ;
        RECT 111.770 47.070 112.720 48.280 ;
      LAYER li1 ;
        RECT 109.700 46.680 111.590 46.850 ;
        RECT 109.700 46.550 109.870 46.680 ;
        RECT 112.370 46.550 112.700 46.890 ;
        RECT 108.610 46.320 109.870 46.550 ;
      LAYER li1 ;
        RECT 110.050 46.370 112.080 46.500 ;
        RECT 112.900 46.370 113.150 48.530 ;
        RECT 113.530 48.500 114.980 48.530 ;
        RECT 113.530 48.330 113.780 48.500 ;
        RECT 113.950 48.330 114.140 48.500 ;
        RECT 114.310 48.330 114.580 48.500 ;
        RECT 114.750 48.330 114.980 48.500 ;
        RECT 113.530 47.460 114.980 48.330 ;
        RECT 116.250 48.450 117.200 48.530 ;
        RECT 116.250 48.280 116.280 48.450 ;
        RECT 116.450 48.280 116.640 48.450 ;
        RECT 116.810 48.280 117.000 48.450 ;
        RECT 117.170 48.280 117.200 48.450 ;
        RECT 110.050 46.330 113.150 46.370 ;
      LAYER li1 ;
        RECT 109.700 46.150 109.870 46.320 ;
      LAYER li1 ;
        RECT 111.910 46.200 113.150 46.330 ;
        RECT 106.560 45.620 107.860 46.020 ;
        RECT 106.250 45.140 107.860 45.620 ;
        RECT 108.570 45.140 109.520 46.100 ;
      LAYER li1 ;
        RECT 109.700 45.980 111.510 46.150 ;
        RECT 109.700 45.270 109.950 45.980 ;
      LAYER li1 ;
        RECT 110.130 45.140 111.080 45.800 ;
      LAYER li1 ;
        RECT 111.260 45.270 111.510 45.980 ;
      LAYER li1 ;
        RECT 111.690 45.140 112.640 46.020 ;
        RECT 112.820 45.270 113.150 46.200 ;
        RECT 113.760 46.020 114.090 46.800 ;
        RECT 114.300 46.470 114.630 47.460 ;
        RECT 116.250 46.950 117.200 48.280 ;
      LAYER li1 ;
        RECT 117.380 46.850 117.630 48.530 ;
      LAYER li1 ;
        RECT 117.810 48.450 118.760 48.530 ;
        RECT 117.810 48.280 117.840 48.450 ;
        RECT 118.010 48.280 118.200 48.450 ;
        RECT 118.370 48.280 118.560 48.450 ;
        RECT 118.730 48.280 118.760 48.450 ;
        RECT 117.810 47.030 118.760 48.280 ;
      LAYER li1 ;
        RECT 118.940 46.850 119.270 48.530 ;
      LAYER li1 ;
        RECT 119.450 48.450 120.400 48.530 ;
        RECT 119.450 48.280 119.480 48.450 ;
        RECT 119.650 48.280 119.840 48.450 ;
        RECT 120.010 48.280 120.200 48.450 ;
        RECT 120.370 48.280 120.400 48.450 ;
        RECT 119.450 47.070 120.400 48.280 ;
      LAYER li1 ;
        RECT 117.380 46.680 119.270 46.850 ;
        RECT 117.380 46.550 117.550 46.680 ;
        RECT 120.050 46.550 120.380 46.890 ;
        RECT 116.290 46.320 117.550 46.550 ;
      LAYER li1 ;
        RECT 117.730 46.370 119.760 46.500 ;
        RECT 120.580 46.370 120.830 48.530 ;
        RECT 121.460 48.500 124.200 48.520 ;
        RECT 121.460 48.330 121.670 48.500 ;
        RECT 121.840 48.330 122.110 48.500 ;
        RECT 122.280 48.330 122.520 48.500 ;
        RECT 122.690 48.330 122.950 48.500 ;
        RECT 123.120 48.330 123.390 48.500 ;
        RECT 123.560 48.330 123.800 48.500 ;
        RECT 123.970 48.330 124.200 48.500 ;
        RECT 121.460 47.450 124.200 48.330 ;
        RECT 125.430 48.450 126.020 48.480 ;
        RECT 125.430 48.280 125.460 48.450 ;
        RECT 125.630 48.280 125.820 48.450 ;
        RECT 125.990 48.280 126.020 48.450 ;
        RECT 117.730 46.330 120.830 46.370 ;
      LAYER li1 ;
        RECT 117.380 46.150 117.550 46.320 ;
      LAYER li1 ;
        RECT 119.590 46.200 120.830 46.330 ;
        RECT 113.760 45.620 115.060 46.020 ;
        RECT 113.450 45.140 115.060 45.620 ;
        RECT 116.250 45.140 117.200 46.100 ;
      LAYER li1 ;
        RECT 117.380 45.980 119.190 46.150 ;
        RECT 117.380 45.270 117.630 45.980 ;
      LAYER li1 ;
        RECT 117.810 45.140 118.760 45.800 ;
      LAYER li1 ;
        RECT 118.940 45.270 119.190 45.980 ;
      LAYER li1 ;
        RECT 119.370 45.140 120.320 46.020 ;
        RECT 120.500 45.270 120.830 46.200 ;
        RECT 121.700 46.130 122.030 46.800 ;
        RECT 122.430 46.470 122.760 47.450 ;
        RECT 122.980 46.130 123.310 46.800 ;
        RECT 123.710 46.470 124.040 47.450 ;
        RECT 124.910 47.300 125.240 48.230 ;
        RECT 125.430 47.500 126.020 48.280 ;
        RECT 126.200 48.410 127.640 48.580 ;
        RECT 126.200 47.300 126.370 48.410 ;
        RECT 124.910 47.130 126.370 47.300 ;
        RECT 121.540 45.130 124.270 46.130 ;
        RECT 124.910 45.270 125.180 47.130 ;
        RECT 126.040 46.630 126.370 47.130 ;
        RECT 126.550 46.920 126.800 48.230 ;
        RECT 127.040 47.610 127.290 48.230 ;
        RECT 127.470 47.960 127.640 48.410 ;
        RECT 127.820 48.450 128.150 48.480 ;
        RECT 127.820 48.280 127.850 48.450 ;
        RECT 128.020 48.280 128.150 48.450 ;
        RECT 127.820 48.140 128.150 48.280 ;
        RECT 128.330 48.410 130.070 48.580 ;
        RECT 128.330 47.960 128.500 48.410 ;
        RECT 127.470 47.790 128.500 47.960 ;
        RECT 128.680 47.610 128.850 48.230 ;
        RECT 129.380 47.970 129.710 48.230 ;
        RECT 127.040 47.440 128.850 47.610 ;
        RECT 129.030 47.440 129.250 47.770 ;
        RECT 128.680 47.260 128.850 47.440 ;
        RECT 126.550 46.690 127.080 46.920 ;
        RECT 126.550 45.770 126.820 46.690 ;
      LAYER li1 ;
        RECT 127.500 46.390 128.040 47.260 ;
      LAYER li1 ;
        RECT 128.680 47.090 128.900 47.260 ;
        RECT 125.360 45.140 126.310 45.770 ;
        RECT 126.490 45.270 126.820 45.770 ;
        RECT 127.000 45.140 127.590 46.020 ;
      LAYER li1 ;
        RECT 127.870 45.400 128.040 46.390 ;
        RECT 128.220 45.580 128.550 46.880 ;
      LAYER li1 ;
        RECT 128.730 46.100 128.900 47.090 ;
        RECT 129.080 46.920 129.250 47.440 ;
        RECT 129.430 47.270 129.600 47.970 ;
        RECT 129.900 47.820 130.070 48.410 ;
        RECT 130.250 48.450 131.200 48.480 ;
        RECT 130.250 48.280 130.280 48.450 ;
        RECT 130.450 48.280 130.640 48.450 ;
        RECT 130.810 48.280 131.000 48.450 ;
        RECT 131.170 48.280 131.200 48.450 ;
        RECT 130.250 48.000 131.200 48.280 ;
        RECT 131.380 48.410 132.410 48.580 ;
        RECT 131.380 47.820 131.550 48.410 ;
        RECT 129.900 47.770 131.550 47.820 ;
        RECT 129.780 47.650 131.550 47.770 ;
        RECT 129.780 47.450 130.110 47.650 ;
        RECT 131.730 47.470 132.060 48.230 ;
        RECT 132.240 48.050 132.410 48.410 ;
        RECT 132.590 48.450 133.540 48.530 ;
        RECT 132.590 48.280 132.620 48.450 ;
        RECT 132.790 48.280 132.980 48.450 ;
        RECT 133.150 48.280 133.340 48.450 ;
        RECT 133.510 48.280 133.540 48.450 ;
        RECT 132.590 48.230 133.540 48.280 ;
        RECT 132.240 47.880 134.050 48.050 ;
        RECT 130.290 47.300 132.060 47.470 ;
        RECT 130.290 47.270 130.460 47.300 ;
        RECT 129.430 47.100 130.460 47.270 ;
        RECT 133.370 47.120 133.700 47.700 ;
        RECT 129.080 46.690 130.110 46.920 ;
        RECT 129.780 46.200 130.110 46.690 ;
        RECT 130.290 46.420 130.460 47.100 ;
        RECT 130.640 46.950 133.700 47.120 ;
        RECT 130.640 46.600 130.970 46.950 ;
      LAYER li1 ;
        RECT 131.410 46.600 133.260 46.770 ;
      LAYER li1 ;
        RECT 130.290 46.250 132.910 46.420 ;
        RECT 128.730 45.600 129.000 46.100 ;
        RECT 130.290 46.020 130.460 46.250 ;
      LAYER li1 ;
        RECT 133.090 46.070 133.260 46.600 ;
      LAYER li1 ;
        RECT 129.450 45.850 130.460 46.020 ;
      LAYER li1 ;
        RECT 130.640 45.900 133.260 46.070 ;
      LAYER li1 ;
        RECT 129.450 45.600 129.780 45.850 ;
      LAYER li1 ;
        RECT 130.640 45.400 130.810 45.900 ;
        RECT 127.870 45.230 130.810 45.400 ;
      LAYER li1 ;
        RECT 131.960 45.140 132.910 45.720 ;
      LAYER li1 ;
        RECT 133.090 45.210 133.260 45.900 ;
      LAYER li1 ;
        RECT 133.440 46.100 133.700 46.950 ;
        RECT 133.880 46.530 134.050 47.880 ;
        RECT 134.230 47.620 134.480 48.530 ;
        RECT 135.290 48.450 136.240 48.480 ;
        RECT 137.070 48.450 137.970 48.480 ;
        RECT 135.290 48.280 135.320 48.450 ;
        RECT 135.490 48.280 135.680 48.450 ;
        RECT 135.850 48.280 136.040 48.450 ;
        RECT 136.210 48.280 136.240 48.450 ;
        RECT 137.240 48.280 137.430 48.450 ;
        RECT 137.600 48.280 137.790 48.450 ;
        RECT 137.960 48.280 137.970 48.450 ;
        RECT 134.230 47.450 135.110 47.620 ;
        RECT 135.290 47.450 136.240 48.280 ;
        RECT 136.640 47.480 136.890 47.950 ;
        RECT 137.070 47.660 137.970 48.280 ;
        RECT 138.580 48.450 139.520 48.510 ;
        RECT 138.580 48.280 138.600 48.450 ;
        RECT 138.770 48.280 138.960 48.450 ;
        RECT 139.130 48.280 139.320 48.450 ;
        RECT 139.490 48.280 139.520 48.450 ;
        RECT 134.430 46.710 134.760 47.210 ;
        RECT 134.940 47.130 135.110 47.450 ;
        RECT 136.640 47.310 137.650 47.480 ;
        RECT 134.940 46.960 137.300 47.130 ;
        RECT 133.880 46.360 135.050 46.530 ;
        RECT 133.440 45.390 133.770 46.100 ;
        RECT 134.230 45.560 134.560 46.100 ;
        RECT 134.770 45.860 135.050 46.360 ;
        RECT 135.230 45.560 135.400 46.960 ;
        RECT 137.480 46.780 137.650 47.310 ;
        RECT 135.610 46.610 137.650 46.780 ;
        RECT 135.610 46.220 135.940 46.610 ;
      LAYER li1 ;
        RECT 136.260 46.150 136.590 46.430 ;
        RECT 136.260 46.040 136.640 46.150 ;
      LAYER li1 ;
        RECT 134.230 45.390 135.400 45.560 ;
      LAYER li1 ;
        RECT 135.580 45.980 136.640 46.040 ;
        RECT 135.580 45.870 136.590 45.980 ;
        RECT 135.580 45.210 135.750 45.870 ;
      LAYER li1 ;
        RECT 137.420 45.770 137.650 46.610 ;
        RECT 138.150 46.780 138.400 47.780 ;
        RECT 138.580 46.970 139.520 48.280 ;
        RECT 138.150 46.450 139.520 46.780 ;
        RECT 138.150 46.270 138.360 46.450 ;
        RECT 138.030 45.770 138.360 46.270 ;
      LAYER li1 ;
        RECT 133.090 45.040 135.750 45.210 ;
      LAYER li1 ;
        RECT 135.930 45.140 136.880 45.690 ;
        RECT 137.420 45.270 137.750 45.770 ;
        RECT 138.540 45.140 139.490 46.270 ;
      LAYER li1 ;
        RECT 139.700 45.440 140.040 48.510 ;
      LAYER li1 ;
        RECT 140.410 48.500 141.860 48.530 ;
        RECT 140.410 48.330 140.660 48.500 ;
        RECT 140.830 48.330 141.020 48.500 ;
        RECT 141.190 48.330 141.460 48.500 ;
        RECT 141.630 48.330 141.860 48.500 ;
        RECT 140.410 47.460 141.860 48.330 ;
        RECT 140.640 46.020 140.970 46.800 ;
        RECT 141.180 46.470 141.510 47.460 ;
        RECT 140.640 45.620 141.940 46.020 ;
        RECT 140.330 45.140 141.940 45.620 ;
        RECT 5.760 44.680 5.920 44.860 ;
        RECT 6.090 44.680 6.400 44.860 ;
        RECT 6.570 44.680 6.880 44.860 ;
        RECT 7.050 44.680 7.360 44.860 ;
        RECT 7.530 44.680 7.840 44.860 ;
        RECT 8.010 44.680 8.320 44.860 ;
        RECT 8.490 44.680 8.800 44.860 ;
        RECT 8.970 44.680 9.280 44.860 ;
        RECT 9.450 44.680 9.760 44.860 ;
        RECT 9.930 44.680 10.240 44.860 ;
        RECT 10.410 44.680 10.720 44.860 ;
        RECT 10.890 44.680 11.200 44.860 ;
        RECT 11.370 44.680 11.680 44.860 ;
        RECT 11.850 44.680 12.160 44.860 ;
        RECT 12.330 44.680 12.640 44.860 ;
        RECT 12.810 44.680 13.120 44.860 ;
        RECT 13.290 44.680 13.600 44.860 ;
        RECT 13.770 44.680 14.080 44.860 ;
        RECT 14.250 44.680 14.560 44.860 ;
        RECT 14.730 44.680 15.040 44.860 ;
        RECT 15.210 44.680 15.520 44.860 ;
        RECT 15.690 44.680 16.000 44.860 ;
        RECT 16.170 44.680 16.480 44.860 ;
        RECT 16.650 44.680 16.960 44.860 ;
        RECT 17.130 44.680 17.440 44.860 ;
        RECT 17.610 44.680 17.920 44.860 ;
        RECT 18.090 44.680 18.400 44.860 ;
        RECT 18.570 44.680 18.880 44.860 ;
        RECT 19.050 44.680 19.360 44.860 ;
        RECT 19.530 44.680 19.840 44.860 ;
        RECT 20.010 44.680 20.320 44.860 ;
        RECT 20.490 44.680 20.800 44.860 ;
        RECT 20.970 44.680 21.280 44.860 ;
        RECT 21.450 44.680 21.760 44.860 ;
        RECT 21.930 44.680 22.240 44.860 ;
        RECT 22.410 44.680 22.720 44.860 ;
        RECT 22.890 44.680 23.200 44.860 ;
        RECT 23.370 44.680 23.680 44.860 ;
        RECT 23.850 44.680 24.160 44.860 ;
        RECT 24.330 44.680 24.640 44.860 ;
        RECT 24.810 44.680 25.120 44.860 ;
        RECT 25.290 44.680 25.600 44.860 ;
        RECT 25.770 44.680 26.080 44.860 ;
        RECT 26.250 44.680 26.560 44.860 ;
        RECT 26.730 44.680 27.040 44.860 ;
        RECT 27.210 44.680 27.520 44.860 ;
        RECT 27.690 44.680 28.000 44.860 ;
        RECT 28.170 44.680 28.480 44.860 ;
        RECT 28.650 44.680 28.960 44.860 ;
        RECT 29.130 44.680 29.440 44.860 ;
        RECT 29.610 44.680 29.920 44.860 ;
        RECT 30.090 44.680 30.400 44.860 ;
        RECT 30.570 44.680 30.880 44.860 ;
        RECT 31.050 44.680 31.360 44.860 ;
        RECT 31.530 44.680 31.840 44.860 ;
        RECT 32.010 44.680 32.320 44.860 ;
        RECT 32.490 44.680 32.800 44.860 ;
        RECT 32.970 44.680 33.280 44.860 ;
        RECT 33.450 44.680 33.760 44.860 ;
        RECT 33.930 44.680 34.240 44.860 ;
        RECT 34.410 44.680 34.720 44.860 ;
        RECT 34.890 44.680 35.200 44.860 ;
        RECT 35.370 44.680 35.680 44.860 ;
        RECT 35.850 44.680 36.160 44.860 ;
        RECT 36.330 44.680 36.640 44.860 ;
        RECT 36.810 44.680 37.120 44.860 ;
        RECT 37.290 44.680 37.600 44.860 ;
        RECT 37.770 44.680 38.080 44.860 ;
        RECT 38.250 44.680 38.560 44.860 ;
        RECT 38.730 44.680 39.040 44.860 ;
        RECT 39.210 44.680 39.520 44.860 ;
        RECT 39.690 44.680 40.000 44.860 ;
        RECT 40.170 44.680 40.480 44.860 ;
        RECT 40.650 44.680 40.960 44.860 ;
        RECT 41.130 44.680 41.440 44.860 ;
        RECT 41.610 44.680 41.920 44.860 ;
        RECT 42.090 44.680 42.400 44.860 ;
        RECT 42.570 44.680 42.880 44.860 ;
        RECT 43.050 44.680 43.360 44.860 ;
        RECT 43.530 44.680 43.840 44.860 ;
        RECT 44.010 44.680 44.320 44.860 ;
        RECT 44.490 44.680 44.800 44.860 ;
        RECT 44.970 44.680 45.280 44.860 ;
        RECT 45.450 44.680 45.760 44.860 ;
        RECT 45.930 44.680 46.240 44.860 ;
        RECT 46.410 44.680 46.720 44.860 ;
        RECT 46.890 44.680 47.200 44.860 ;
        RECT 47.370 44.680 47.680 44.860 ;
        RECT 47.850 44.680 48.160 44.860 ;
        RECT 48.330 44.680 48.640 44.860 ;
        RECT 48.810 44.680 49.120 44.860 ;
        RECT 49.290 44.680 49.600 44.860 ;
        RECT 49.770 44.680 50.080 44.860 ;
        RECT 50.250 44.680 50.400 44.860 ;
        RECT 50.880 44.680 51.040 44.860 ;
        RECT 51.210 44.680 51.520 44.860 ;
        RECT 51.690 44.680 52.000 44.860 ;
        RECT 52.170 44.680 52.480 44.860 ;
        RECT 52.650 44.680 52.960 44.860 ;
        RECT 53.130 44.680 53.440 44.860 ;
        RECT 53.610 44.680 53.920 44.860 ;
        RECT 54.090 44.680 54.400 44.860 ;
        RECT 54.570 44.680 54.880 44.860 ;
        RECT 55.050 44.680 55.360 44.860 ;
        RECT 55.530 44.680 55.840 44.860 ;
        RECT 56.010 44.680 56.320 44.860 ;
        RECT 56.490 44.680 56.800 44.860 ;
        RECT 56.970 44.680 57.280 44.860 ;
        RECT 57.450 44.680 57.760 44.860 ;
        RECT 57.930 44.680 58.240 44.860 ;
        RECT 58.410 44.680 58.720 44.860 ;
        RECT 58.890 44.680 59.200 44.860 ;
        RECT 59.370 44.680 59.680 44.860 ;
        RECT 59.850 44.680 60.160 44.860 ;
        RECT 60.330 44.680 60.640 44.860 ;
        RECT 60.810 44.680 61.120 44.860 ;
        RECT 61.290 44.680 61.600 44.860 ;
        RECT 61.770 44.680 62.080 44.860 ;
        RECT 62.250 44.680 62.560 44.860 ;
        RECT 62.730 44.680 63.040 44.860 ;
        RECT 63.210 44.680 63.520 44.860 ;
        RECT 63.690 44.680 64.000 44.860 ;
        RECT 64.170 44.680 64.480 44.860 ;
        RECT 64.650 44.680 64.960 44.860 ;
        RECT 65.130 44.680 65.440 44.860 ;
        RECT 65.610 44.680 65.920 44.860 ;
        RECT 66.090 44.680 66.400 44.860 ;
        RECT 66.570 44.680 66.880 44.860 ;
        RECT 67.050 44.680 67.360 44.860 ;
        RECT 67.530 44.680 67.840 44.860 ;
        RECT 68.010 44.680 68.320 44.860 ;
        RECT 68.490 44.680 68.800 44.860 ;
        RECT 68.970 44.680 69.280 44.860 ;
        RECT 69.450 44.680 69.760 44.860 ;
        RECT 69.930 44.680 70.240 44.860 ;
        RECT 70.410 44.680 70.720 44.860 ;
        RECT 70.890 44.680 71.200 44.860 ;
        RECT 71.370 44.680 71.680 44.860 ;
        RECT 71.850 44.680 72.160 44.860 ;
        RECT 72.330 44.680 72.640 44.860 ;
        RECT 72.810 44.680 73.120 44.860 ;
        RECT 73.290 44.680 73.600 44.860 ;
        RECT 73.770 44.680 74.080 44.860 ;
        RECT 74.250 44.680 74.560 44.860 ;
        RECT 74.730 44.680 75.040 44.860 ;
        RECT 75.210 44.680 75.520 44.860 ;
        RECT 75.690 44.680 76.000 44.860 ;
        RECT 76.170 44.680 76.480 44.860 ;
        RECT 76.650 44.680 76.960 44.860 ;
        RECT 77.130 44.680 77.440 44.860 ;
        RECT 77.610 44.680 77.920 44.860 ;
        RECT 78.090 44.680 78.400 44.860 ;
        RECT 78.570 44.680 78.880 44.860 ;
        RECT 79.050 44.680 79.360 44.860 ;
        RECT 79.530 44.680 79.840 44.860 ;
        RECT 80.010 44.680 80.320 44.860 ;
        RECT 80.490 44.680 80.800 44.860 ;
        RECT 80.970 44.680 81.280 44.860 ;
        RECT 81.450 44.680 81.760 44.860 ;
        RECT 81.930 44.680 82.240 44.860 ;
        RECT 82.410 44.680 82.720 44.860 ;
        RECT 82.890 44.680 83.200 44.860 ;
        RECT 83.370 44.680 83.680 44.860 ;
        RECT 83.850 44.680 84.160 44.860 ;
        RECT 84.330 44.680 84.640 44.860 ;
        RECT 84.810 44.680 85.120 44.860 ;
        RECT 85.290 44.680 85.600 44.860 ;
        RECT 85.770 44.680 86.080 44.860 ;
        RECT 86.250 44.680 86.560 44.860 ;
        RECT 86.730 44.680 87.040 44.860 ;
        RECT 87.210 44.680 87.520 44.860 ;
        RECT 87.690 44.680 88.000 44.860 ;
        RECT 88.170 44.680 88.480 44.860 ;
        RECT 88.650 44.680 88.960 44.860 ;
        RECT 89.130 44.680 89.440 44.860 ;
        RECT 89.610 44.680 89.920 44.860 ;
        RECT 90.090 44.680 90.400 44.860 ;
        RECT 90.570 44.680 90.880 44.860 ;
        RECT 91.050 44.680 91.360 44.860 ;
        RECT 91.530 44.680 91.840 44.860 ;
        RECT 92.010 44.680 92.320 44.860 ;
        RECT 92.490 44.680 92.800 44.860 ;
        RECT 92.970 44.680 93.280 44.860 ;
        RECT 93.450 44.680 93.760 44.860 ;
        RECT 93.930 44.680 94.240 44.860 ;
        RECT 94.410 44.680 94.560 44.860 ;
        RECT 95.040 44.680 95.200 44.860 ;
        RECT 95.370 44.680 95.680 44.860 ;
        RECT 95.850 44.680 96.160 44.860 ;
        RECT 96.330 44.680 96.640 44.860 ;
        RECT 96.810 44.680 97.120 44.860 ;
        RECT 97.290 44.680 97.600 44.860 ;
        RECT 97.770 44.680 98.080 44.860 ;
        RECT 98.250 44.680 98.560 44.860 ;
        RECT 98.730 44.680 99.040 44.860 ;
        RECT 99.210 44.680 99.520 44.860 ;
        RECT 99.690 44.680 100.000 44.860 ;
        RECT 100.170 44.680 100.480 44.860 ;
        RECT 100.650 44.680 100.960 44.860 ;
        RECT 101.130 44.680 101.440 44.860 ;
        RECT 101.610 44.680 101.920 44.860 ;
        RECT 102.090 44.680 102.400 44.860 ;
        RECT 102.570 44.680 102.880 44.860 ;
        RECT 103.050 44.680 103.360 44.860 ;
        RECT 103.530 44.680 103.840 44.860 ;
        RECT 104.010 44.680 104.320 44.860 ;
        RECT 104.490 44.680 104.800 44.860 ;
        RECT 104.970 44.680 105.280 44.860 ;
        RECT 105.450 44.680 105.760 44.860 ;
        RECT 105.930 44.680 106.240 44.860 ;
        RECT 106.410 44.680 106.720 44.860 ;
        RECT 106.890 44.680 107.200 44.860 ;
        RECT 107.370 44.680 107.680 44.860 ;
        RECT 107.850 44.680 108.000 44.860 ;
        RECT 108.480 44.680 108.640 44.860 ;
        RECT 108.810 44.680 109.120 44.860 ;
        RECT 109.290 44.680 109.600 44.860 ;
        RECT 109.770 44.680 110.080 44.860 ;
        RECT 110.250 44.680 110.560 44.860 ;
        RECT 110.730 44.680 111.040 44.860 ;
        RECT 111.210 44.680 111.520 44.860 ;
        RECT 111.690 44.680 112.000 44.860 ;
        RECT 112.170 44.680 112.480 44.860 ;
        RECT 112.650 44.680 112.960 44.860 ;
        RECT 113.130 44.680 113.440 44.860 ;
        RECT 113.610 44.680 113.920 44.860 ;
        RECT 114.090 44.680 114.400 44.860 ;
        RECT 114.570 44.680 114.880 44.860 ;
        RECT 115.050 44.680 115.360 44.860 ;
        RECT 115.530 44.680 115.840 44.860 ;
        RECT 116.010 44.680 116.320 44.860 ;
        RECT 116.490 44.680 116.800 44.860 ;
        RECT 116.970 44.680 117.280 44.860 ;
        RECT 117.450 44.680 117.760 44.860 ;
        RECT 117.930 44.680 118.240 44.860 ;
        RECT 118.410 44.680 118.720 44.860 ;
        RECT 118.890 44.680 119.200 44.860 ;
        RECT 119.370 44.680 119.680 44.860 ;
        RECT 119.850 44.680 120.160 44.860 ;
        RECT 120.330 44.680 120.640 44.860 ;
        RECT 120.810 44.680 121.120 44.860 ;
        RECT 121.290 44.680 121.600 44.860 ;
        RECT 121.770 44.680 122.080 44.860 ;
        RECT 122.250 44.680 122.560 44.860 ;
        RECT 122.730 44.680 123.040 44.860 ;
        RECT 123.210 44.680 123.520 44.860 ;
        RECT 123.690 44.680 124.000 44.860 ;
        RECT 124.170 44.680 124.480 44.860 ;
        RECT 124.650 44.680 124.960 44.860 ;
        RECT 125.130 44.680 125.440 44.860 ;
        RECT 125.610 44.680 125.920 44.860 ;
        RECT 126.090 44.680 126.400 44.860 ;
        RECT 126.570 44.680 126.880 44.860 ;
        RECT 127.050 44.680 127.360 44.860 ;
        RECT 127.530 44.680 127.840 44.860 ;
        RECT 128.010 44.680 128.320 44.860 ;
        RECT 128.490 44.680 128.800 44.860 ;
        RECT 128.970 44.680 129.280 44.860 ;
        RECT 129.450 44.680 129.760 44.860 ;
        RECT 129.930 44.680 130.240 44.860 ;
        RECT 130.410 44.680 130.720 44.860 ;
        RECT 130.890 44.680 131.200 44.860 ;
        RECT 131.370 44.680 131.680 44.860 ;
        RECT 131.850 44.680 132.160 44.860 ;
        RECT 132.330 44.680 132.640 44.860 ;
        RECT 132.810 44.680 133.120 44.860 ;
        RECT 133.290 44.680 133.600 44.860 ;
        RECT 133.770 44.680 134.080 44.860 ;
        RECT 134.250 44.680 134.560 44.860 ;
        RECT 134.730 44.680 135.040 44.860 ;
        RECT 135.210 44.680 135.520 44.860 ;
        RECT 135.690 44.680 136.000 44.860 ;
        RECT 136.170 44.680 136.480 44.860 ;
        RECT 136.650 44.680 136.960 44.860 ;
        RECT 137.130 44.680 137.440 44.860 ;
        RECT 137.610 44.680 137.920 44.860 ;
        RECT 138.090 44.680 138.400 44.860 ;
        RECT 138.570 44.680 138.880 44.860 ;
        RECT 139.050 44.680 139.360 44.860 ;
        RECT 139.530 44.680 139.840 44.860 ;
        RECT 140.010 44.680 140.320 44.860 ;
        RECT 140.490 44.680 140.800 44.860 ;
        RECT 140.970 44.680 141.280 44.860 ;
        RECT 141.450 44.680 141.760 44.860 ;
        RECT 141.930 44.680 142.080 44.860 ;
        RECT 6.340 44.380 9.070 44.410 ;
        RECT 6.340 44.210 6.510 44.380 ;
        RECT 6.680 44.210 6.950 44.380 ;
        RECT 7.120 44.210 7.360 44.380 ;
        RECT 7.530 44.210 7.790 44.380 ;
        RECT 7.960 44.210 8.230 44.380 ;
        RECT 8.400 44.210 8.640 44.380 ;
        RECT 8.810 44.210 9.070 44.380 ;
        RECT 6.340 43.410 9.070 44.210 ;
        RECT 9.770 44.370 11.380 44.400 ;
        RECT 9.770 44.200 9.820 44.370 ;
        RECT 9.990 44.200 10.260 44.370 ;
        RECT 10.430 44.200 10.700 44.370 ;
        RECT 10.870 44.200 11.110 44.370 ;
        RECT 11.280 44.200 11.380 44.370 ;
        RECT 9.770 43.920 11.380 44.200 ;
        RECT 10.080 43.520 11.380 43.920 ;
        RECT 12.570 44.370 13.160 44.400 ;
        RECT 12.570 44.200 12.600 44.370 ;
        RECT 12.770 44.200 12.960 44.370 ;
        RECT 13.130 44.200 13.160 44.370 ;
        RECT 14.090 44.370 15.700 44.400 ;
        RECT 16.390 44.370 17.640 44.400 ;
        RECT 18.410 44.370 20.020 44.400 ;
        RECT 20.800 44.370 21.690 44.400 ;
        RECT 23.690 44.370 25.300 44.400 ;
        RECT 26.080 44.370 26.970 44.400 ;
        RECT 28.970 44.370 30.580 44.400 ;
        RECT 6.500 42.740 6.830 43.410 ;
        RECT 7.230 42.090 7.560 43.070 ;
        RECT 7.780 42.740 8.110 43.410 ;
        RECT 8.510 42.090 8.840 43.070 ;
        RECT 10.080 42.740 10.410 43.520 ;
        RECT 12.570 43.440 13.160 44.200 ;
        RECT 6.260 41.210 9.000 42.090 ;
        RECT 10.620 42.080 10.950 43.070 ;
      LAYER li1 ;
        RECT 12.610 42.830 13.320 43.220 ;
        RECT 13.500 42.590 13.830 44.270 ;
      LAYER li1 ;
        RECT 14.090 44.200 14.140 44.370 ;
        RECT 14.310 44.200 14.580 44.370 ;
        RECT 14.750 44.200 15.020 44.370 ;
        RECT 15.190 44.200 15.430 44.370 ;
        RECT 15.600 44.200 15.700 44.370 ;
        RECT 14.090 43.920 15.700 44.200 ;
        RECT 14.400 43.520 15.700 43.920 ;
        RECT 14.400 42.740 14.730 43.520 ;
        RECT 6.260 41.040 6.470 41.210 ;
        RECT 6.640 41.040 6.910 41.210 ;
        RECT 7.080 41.040 7.320 41.210 ;
        RECT 7.490 41.040 7.750 41.210 ;
        RECT 7.920 41.040 8.190 41.210 ;
        RECT 8.360 41.040 8.600 41.210 ;
        RECT 8.770 41.040 9.000 41.210 ;
        RECT 6.260 41.020 9.000 41.040 ;
        RECT 9.850 41.210 11.300 42.080 ;
        RECT 9.850 41.040 10.100 41.210 ;
        RECT 10.270 41.040 10.460 41.210 ;
        RECT 10.630 41.040 10.900 41.210 ;
        RECT 11.070 41.040 11.300 41.210 ;
        RECT 9.850 41.010 11.300 41.040 ;
        RECT 12.570 41.260 13.160 42.590 ;
        RECT 12.570 41.090 12.600 41.260 ;
        RECT 12.770 41.090 12.960 41.260 ;
        RECT 13.130 41.090 13.160 41.260 ;
        RECT 12.570 41.010 13.160 41.090 ;
      LAYER li1 ;
        RECT 13.440 41.010 13.830 42.590 ;
      LAYER li1 ;
        RECT 14.940 42.080 15.270 43.070 ;
      LAYER li1 ;
        RECT 15.960 42.590 16.210 44.270 ;
      LAYER li1 ;
        RECT 16.560 44.200 16.750 44.370 ;
        RECT 16.920 44.200 17.110 44.370 ;
        RECT 17.280 44.200 17.470 44.370 ;
        RECT 16.390 43.830 17.640 44.200 ;
        RECT 17.820 43.650 18.070 44.270 ;
        RECT 18.410 44.200 18.460 44.370 ;
        RECT 18.630 44.200 18.900 44.370 ;
        RECT 19.070 44.200 19.340 44.370 ;
        RECT 19.510 44.200 19.750 44.370 ;
        RECT 19.920 44.200 20.020 44.370 ;
        RECT 18.410 43.920 20.020 44.200 ;
        RECT 16.520 43.480 18.070 43.650 ;
        RECT 16.520 43.020 16.850 43.480 ;
        RECT 14.170 41.210 15.620 42.080 ;
        RECT 14.170 41.040 14.420 41.210 ;
        RECT 14.590 41.040 14.780 41.210 ;
        RECT 14.950 41.040 15.220 41.210 ;
        RECT 15.390 41.040 15.620 41.210 ;
        RECT 14.170 41.010 15.620 41.040 ;
      LAYER li1 ;
        RECT 15.960 41.010 16.390 42.590 ;
      LAYER li1 ;
        RECT 16.570 41.260 17.130 42.590 ;
      LAYER li1 ;
        RECT 17.310 41.510 17.640 43.300 ;
      LAYER li1 ;
        RECT 17.820 41.760 18.070 43.480 ;
        RECT 18.720 43.520 20.020 43.920 ;
        RECT 20.290 43.660 20.620 44.270 ;
        RECT 20.970 44.200 21.160 44.370 ;
        RECT 21.330 44.200 21.520 44.370 ;
        RECT 20.800 43.840 21.690 44.200 ;
        RECT 21.870 43.660 22.200 44.270 ;
        RECT 18.720 42.740 19.050 43.520 ;
        RECT 20.290 43.490 22.200 43.660 ;
        RECT 20.290 43.440 20.620 43.490 ;
      LAYER li1 ;
        RECT 22.650 43.310 22.980 44.270 ;
      LAYER li1 ;
        RECT 23.690 44.200 23.740 44.370 ;
        RECT 23.910 44.200 24.180 44.370 ;
        RECT 24.350 44.200 24.620 44.370 ;
        RECT 24.790 44.200 25.030 44.370 ;
        RECT 25.200 44.200 25.300 44.370 ;
        RECT 23.690 43.920 25.300 44.200 ;
        RECT 19.260 42.080 19.590 43.070 ;
      LAYER li1 ;
        RECT 20.290 42.930 21.020 43.260 ;
        RECT 21.230 43.010 21.960 43.260 ;
        RECT 22.140 43.140 22.980 43.310 ;
      LAYER li1 ;
        RECT 24.000 43.520 25.300 43.920 ;
        RECT 25.570 43.660 25.900 44.270 ;
        RECT 26.250 44.200 26.440 44.370 ;
        RECT 26.610 44.200 26.800 44.370 ;
        RECT 26.080 43.840 26.970 44.200 ;
        RECT 27.150 43.660 27.480 44.270 ;
      LAYER li1 ;
        RECT 22.140 42.830 22.310 43.140 ;
        RECT 21.730 42.660 22.310 42.830 ;
      LAYER li1 ;
        RECT 16.570 41.090 16.580 41.260 ;
        RECT 16.750 41.090 16.940 41.260 ;
        RECT 17.110 41.090 17.130 41.260 ;
        RECT 16.570 41.010 17.130 41.090 ;
        RECT 18.490 41.210 19.940 42.080 ;
        RECT 18.490 41.040 18.740 41.210 ;
        RECT 18.910 41.040 19.100 41.210 ;
        RECT 19.270 41.040 19.540 41.210 ;
        RECT 19.710 41.040 19.940 41.210 ;
        RECT 18.490 41.010 19.940 41.040 ;
        RECT 20.250 41.260 21.200 42.590 ;
        RECT 20.250 41.090 20.280 41.260 ;
        RECT 20.450 41.090 20.640 41.260 ;
        RECT 20.810 41.090 21.000 41.260 ;
        RECT 21.170 41.090 21.200 41.260 ;
        RECT 20.250 41.010 21.200 41.090 ;
      LAYER li1 ;
        RECT 21.730 41.010 22.200 42.660 ;
        RECT 22.490 42.650 23.400 42.960 ;
      LAYER li1 ;
        RECT 24.000 42.740 24.330 43.520 ;
        RECT 25.570 43.490 27.480 43.660 ;
        RECT 25.570 43.440 25.900 43.490 ;
      LAYER li1 ;
        RECT 27.930 43.310 28.260 44.270 ;
      LAYER li1 ;
        RECT 28.970 44.200 29.020 44.370 ;
        RECT 29.190 44.200 29.460 44.370 ;
        RECT 29.630 44.200 29.900 44.370 ;
        RECT 30.070 44.200 30.310 44.370 ;
        RECT 30.480 44.200 30.580 44.370 ;
        RECT 28.970 43.920 30.580 44.200 ;
        RECT 22.380 41.260 23.330 42.470 ;
        RECT 24.540 42.080 24.870 43.070 ;
      LAYER li1 ;
        RECT 25.570 42.930 26.300 43.260 ;
        RECT 26.510 43.010 27.240 43.260 ;
        RECT 27.420 43.140 28.260 43.310 ;
      LAYER li1 ;
        RECT 29.280 43.520 30.580 43.920 ;
        RECT 30.810 44.370 31.760 44.400 ;
        RECT 30.810 44.200 30.840 44.370 ;
        RECT 31.010 44.200 31.200 44.370 ;
        RECT 31.370 44.200 31.560 44.370 ;
        RECT 31.730 44.200 31.760 44.370 ;
        RECT 32.370 44.370 33.320 44.400 ;
      LAYER li1 ;
        RECT 27.420 42.830 27.590 43.140 ;
        RECT 27.010 42.660 27.590 42.830 ;
      LAYER li1 ;
        RECT 22.380 41.090 22.410 41.260 ;
        RECT 22.580 41.090 22.770 41.260 ;
        RECT 22.940 41.090 23.130 41.260 ;
        RECT 23.300 41.090 23.330 41.260 ;
        RECT 22.380 41.010 23.330 41.090 ;
        RECT 23.770 41.210 25.220 42.080 ;
        RECT 23.770 41.040 24.020 41.210 ;
        RECT 24.190 41.040 24.380 41.210 ;
        RECT 24.550 41.040 24.820 41.210 ;
        RECT 24.990 41.040 25.220 41.210 ;
        RECT 23.770 41.010 25.220 41.040 ;
        RECT 25.530 41.260 26.480 42.590 ;
        RECT 25.530 41.090 25.560 41.260 ;
        RECT 25.730 41.090 25.920 41.260 ;
        RECT 26.090 41.090 26.280 41.260 ;
        RECT 26.450 41.090 26.480 41.260 ;
        RECT 25.530 41.010 26.480 41.090 ;
      LAYER li1 ;
        RECT 27.010 41.010 27.480 42.660 ;
        RECT 27.770 42.650 28.680 42.960 ;
      LAYER li1 ;
        RECT 29.280 42.740 29.610 43.520 ;
        RECT 30.810 43.440 31.760 44.200 ;
      LAYER li1 ;
        RECT 31.940 43.560 32.190 44.270 ;
      LAYER li1 ;
        RECT 32.370 44.200 32.400 44.370 ;
        RECT 32.570 44.200 32.760 44.370 ;
        RECT 32.930 44.200 33.120 44.370 ;
        RECT 33.290 44.200 33.320 44.370 ;
        RECT 33.930 44.370 34.880 44.400 ;
        RECT 32.370 43.740 33.320 44.200 ;
      LAYER li1 ;
        RECT 33.500 43.560 33.750 44.270 ;
        RECT 31.940 43.390 33.750 43.560 ;
      LAYER li1 ;
        RECT 33.930 44.200 33.960 44.370 ;
        RECT 34.130 44.200 34.320 44.370 ;
        RECT 34.490 44.200 34.680 44.370 ;
        RECT 34.850 44.200 34.880 44.370 ;
        RECT 35.690 44.370 37.300 44.400 ;
        RECT 33.930 43.520 34.880 44.200 ;
      LAYER li1 ;
        RECT 31.940 43.220 32.110 43.390 ;
      LAYER li1 ;
        RECT 35.060 43.340 35.390 44.270 ;
        RECT 35.690 44.200 35.740 44.370 ;
        RECT 35.910 44.200 36.180 44.370 ;
        RECT 36.350 44.200 36.620 44.370 ;
        RECT 36.790 44.200 37.030 44.370 ;
        RECT 37.200 44.200 37.300 44.370 ;
        RECT 35.690 43.920 37.300 44.200 ;
        RECT 27.660 41.260 28.610 42.470 ;
        RECT 29.820 42.080 30.150 43.070 ;
      LAYER li1 ;
        RECT 30.850 42.990 32.110 43.220 ;
      LAYER li1 ;
        RECT 34.150 43.210 35.390 43.340 ;
        RECT 32.290 43.170 35.390 43.210 ;
        RECT 32.290 43.040 34.320 43.170 ;
      LAYER li1 ;
        RECT 31.940 42.860 32.110 42.990 ;
        RECT 31.940 42.690 33.830 42.860 ;
      LAYER li1 ;
        RECT 27.660 41.090 27.690 41.260 ;
        RECT 27.860 41.090 28.050 41.260 ;
        RECT 28.220 41.090 28.410 41.260 ;
        RECT 28.580 41.090 28.610 41.260 ;
        RECT 27.660 41.010 28.610 41.090 ;
        RECT 29.050 41.210 30.500 42.080 ;
        RECT 29.050 41.040 29.300 41.210 ;
        RECT 29.470 41.040 29.660 41.210 ;
        RECT 29.830 41.040 30.100 41.210 ;
        RECT 30.270 41.040 30.500 41.210 ;
        RECT 29.050 41.010 30.500 41.040 ;
        RECT 30.810 41.260 31.760 42.590 ;
        RECT 30.810 41.090 30.840 41.260 ;
        RECT 31.010 41.090 31.200 41.260 ;
        RECT 31.370 41.090 31.560 41.260 ;
        RECT 31.730 41.090 31.760 41.260 ;
        RECT 30.810 41.010 31.760 41.090 ;
      LAYER li1 ;
        RECT 31.940 41.010 32.190 42.690 ;
      LAYER li1 ;
        RECT 32.370 41.260 33.320 42.510 ;
        RECT 32.370 41.090 32.400 41.260 ;
        RECT 32.570 41.090 32.760 41.260 ;
        RECT 32.930 41.090 33.120 41.260 ;
        RECT 33.290 41.090 33.320 41.260 ;
        RECT 32.370 41.010 33.320 41.090 ;
      LAYER li1 ;
        RECT 33.500 41.010 33.830 42.690 ;
        RECT 34.610 42.650 34.940 42.990 ;
      LAYER li1 ;
        RECT 34.010 41.260 34.960 42.470 ;
        RECT 34.010 41.090 34.040 41.260 ;
        RECT 34.210 41.090 34.400 41.260 ;
        RECT 34.570 41.090 34.760 41.260 ;
        RECT 34.930 41.090 34.960 41.260 ;
        RECT 34.010 41.010 34.960 41.090 ;
        RECT 35.140 41.010 35.390 43.170 ;
        RECT 36.000 43.520 37.300 43.920 ;
        RECT 37.530 44.370 38.120 44.400 ;
        RECT 37.530 44.200 37.560 44.370 ;
        RECT 37.730 44.200 37.920 44.370 ;
        RECT 38.090 44.200 38.120 44.370 ;
        RECT 39.050 44.370 40.660 44.400 ;
        RECT 36.000 42.740 36.330 43.520 ;
        RECT 37.530 43.440 38.120 44.200 ;
        RECT 36.540 42.080 36.870 43.070 ;
      LAYER li1 ;
        RECT 37.570 42.830 38.280 43.220 ;
        RECT 38.460 42.590 38.790 44.270 ;
      LAYER li1 ;
        RECT 39.050 44.200 39.100 44.370 ;
        RECT 39.270 44.200 39.540 44.370 ;
        RECT 39.710 44.200 39.980 44.370 ;
        RECT 40.150 44.200 40.390 44.370 ;
        RECT 40.560 44.200 40.660 44.370 ;
        RECT 39.050 43.920 40.660 44.200 ;
        RECT 39.360 43.520 40.660 43.920 ;
        RECT 40.890 44.370 41.840 44.400 ;
        RECT 40.890 44.200 40.920 44.370 ;
        RECT 41.090 44.200 41.280 44.370 ;
        RECT 41.450 44.200 41.640 44.370 ;
        RECT 41.810 44.200 41.840 44.370 ;
        RECT 42.450 44.370 43.400 44.400 ;
        RECT 39.360 42.740 39.690 43.520 ;
        RECT 40.890 43.440 41.840 44.200 ;
      LAYER li1 ;
        RECT 42.020 43.560 42.270 44.270 ;
      LAYER li1 ;
        RECT 42.450 44.200 42.480 44.370 ;
        RECT 42.650 44.200 42.840 44.370 ;
        RECT 43.010 44.200 43.200 44.370 ;
        RECT 43.370 44.200 43.400 44.370 ;
        RECT 44.010 44.370 44.960 44.400 ;
        RECT 42.450 43.740 43.400 44.200 ;
      LAYER li1 ;
        RECT 43.580 43.560 43.830 44.270 ;
        RECT 42.020 43.390 43.830 43.560 ;
      LAYER li1 ;
        RECT 44.010 44.200 44.040 44.370 ;
        RECT 44.210 44.200 44.400 44.370 ;
        RECT 44.570 44.200 44.760 44.370 ;
        RECT 44.930 44.200 44.960 44.370 ;
        RECT 45.770 44.370 47.380 44.400 ;
        RECT 44.010 43.520 44.960 44.200 ;
      LAYER li1 ;
        RECT 42.020 43.220 42.190 43.390 ;
      LAYER li1 ;
        RECT 45.140 43.340 45.470 44.270 ;
        RECT 45.770 44.200 45.820 44.370 ;
        RECT 45.990 44.200 46.260 44.370 ;
        RECT 46.430 44.200 46.700 44.370 ;
        RECT 46.870 44.200 47.110 44.370 ;
        RECT 47.280 44.200 47.380 44.370 ;
        RECT 45.770 43.920 47.380 44.200 ;
        RECT 35.770 41.210 37.220 42.080 ;
        RECT 35.770 41.040 36.020 41.210 ;
        RECT 36.190 41.040 36.380 41.210 ;
        RECT 36.550 41.040 36.820 41.210 ;
        RECT 36.990 41.040 37.220 41.210 ;
        RECT 35.770 41.010 37.220 41.040 ;
        RECT 37.530 41.260 38.120 42.590 ;
        RECT 37.530 41.090 37.560 41.260 ;
        RECT 37.730 41.090 37.920 41.260 ;
        RECT 38.090 41.090 38.120 41.260 ;
        RECT 37.530 41.010 38.120 41.090 ;
      LAYER li1 ;
        RECT 38.400 41.010 38.790 42.590 ;
      LAYER li1 ;
        RECT 39.900 42.080 40.230 43.070 ;
      LAYER li1 ;
        RECT 40.930 42.990 42.190 43.220 ;
      LAYER li1 ;
        RECT 44.230 43.210 45.470 43.340 ;
        RECT 42.370 43.170 45.470 43.210 ;
        RECT 42.370 43.040 44.400 43.170 ;
      LAYER li1 ;
        RECT 42.020 42.860 42.190 42.990 ;
        RECT 42.020 42.690 43.910 42.860 ;
      LAYER li1 ;
        RECT 39.130 41.210 40.580 42.080 ;
        RECT 39.130 41.040 39.380 41.210 ;
        RECT 39.550 41.040 39.740 41.210 ;
        RECT 39.910 41.040 40.180 41.210 ;
        RECT 40.350 41.040 40.580 41.210 ;
        RECT 39.130 41.010 40.580 41.040 ;
        RECT 40.890 41.260 41.840 42.590 ;
        RECT 40.890 41.090 40.920 41.260 ;
        RECT 41.090 41.090 41.280 41.260 ;
        RECT 41.450 41.090 41.640 41.260 ;
        RECT 41.810 41.090 41.840 41.260 ;
        RECT 40.890 41.010 41.840 41.090 ;
      LAYER li1 ;
        RECT 42.020 41.010 42.270 42.690 ;
      LAYER li1 ;
        RECT 42.450 41.260 43.400 42.510 ;
        RECT 42.450 41.090 42.480 41.260 ;
        RECT 42.650 41.090 42.840 41.260 ;
        RECT 43.010 41.090 43.200 41.260 ;
        RECT 43.370 41.090 43.400 41.260 ;
        RECT 42.450 41.010 43.400 41.090 ;
      LAYER li1 ;
        RECT 43.580 41.010 43.910 42.690 ;
        RECT 44.690 42.650 45.020 42.990 ;
      LAYER li1 ;
        RECT 44.090 41.260 45.040 42.470 ;
        RECT 44.090 41.090 44.120 41.260 ;
        RECT 44.290 41.090 44.480 41.260 ;
        RECT 44.650 41.090 44.840 41.260 ;
        RECT 45.010 41.090 45.040 41.260 ;
        RECT 44.090 41.010 45.040 41.090 ;
        RECT 45.220 41.010 45.470 43.170 ;
        RECT 46.080 43.520 47.380 43.920 ;
        RECT 47.610 44.370 48.560 44.400 ;
        RECT 47.610 44.200 47.640 44.370 ;
        RECT 47.810 44.200 48.000 44.370 ;
        RECT 48.170 44.200 48.360 44.370 ;
        RECT 48.530 44.200 48.560 44.370 ;
        RECT 49.170 44.370 50.120 44.400 ;
        RECT 46.080 42.740 46.410 43.520 ;
        RECT 47.610 43.440 48.560 44.200 ;
      LAYER li1 ;
        RECT 48.740 43.560 48.990 44.270 ;
      LAYER li1 ;
        RECT 49.170 44.200 49.200 44.370 ;
        RECT 49.370 44.200 49.560 44.370 ;
        RECT 49.730 44.200 49.920 44.370 ;
        RECT 50.090 44.200 50.120 44.370 ;
        RECT 50.730 44.370 51.680 44.400 ;
        RECT 49.170 43.740 50.120 44.200 ;
      LAYER li1 ;
        RECT 50.300 43.560 50.550 44.270 ;
        RECT 48.740 43.390 50.550 43.560 ;
      LAYER li1 ;
        RECT 50.730 44.200 50.760 44.370 ;
        RECT 50.930 44.200 51.120 44.370 ;
        RECT 51.290 44.200 51.480 44.370 ;
        RECT 51.650 44.200 51.680 44.370 ;
        RECT 52.490 44.370 54.100 44.400 ;
        RECT 50.730 43.520 51.680 44.200 ;
      LAYER li1 ;
        RECT 48.740 43.220 48.910 43.390 ;
      LAYER li1 ;
        RECT 51.860 43.340 52.190 44.270 ;
        RECT 52.490 44.200 52.540 44.370 ;
        RECT 52.710 44.200 52.980 44.370 ;
        RECT 53.150 44.200 53.420 44.370 ;
        RECT 53.590 44.200 53.830 44.370 ;
        RECT 54.000 44.200 54.100 44.370 ;
        RECT 52.490 43.920 54.100 44.200 ;
        RECT 46.620 42.080 46.950 43.070 ;
      LAYER li1 ;
        RECT 47.650 42.990 48.910 43.220 ;
      LAYER li1 ;
        RECT 50.950 43.210 52.190 43.340 ;
        RECT 49.090 43.170 52.190 43.210 ;
        RECT 49.090 43.040 51.120 43.170 ;
      LAYER li1 ;
        RECT 48.740 42.860 48.910 42.990 ;
        RECT 48.740 42.690 50.630 42.860 ;
      LAYER li1 ;
        RECT 45.850 41.210 47.300 42.080 ;
        RECT 45.850 41.040 46.100 41.210 ;
        RECT 46.270 41.040 46.460 41.210 ;
        RECT 46.630 41.040 46.900 41.210 ;
        RECT 47.070 41.040 47.300 41.210 ;
        RECT 45.850 41.010 47.300 41.040 ;
        RECT 47.610 41.260 48.560 42.590 ;
        RECT 47.610 41.090 47.640 41.260 ;
        RECT 47.810 41.090 48.000 41.260 ;
        RECT 48.170 41.090 48.360 41.260 ;
        RECT 48.530 41.090 48.560 41.260 ;
        RECT 47.610 41.010 48.560 41.090 ;
      LAYER li1 ;
        RECT 48.740 41.010 48.990 42.690 ;
      LAYER li1 ;
        RECT 49.170 41.260 50.120 42.510 ;
        RECT 49.170 41.090 49.200 41.260 ;
        RECT 49.370 41.090 49.560 41.260 ;
        RECT 49.730 41.090 49.920 41.260 ;
        RECT 50.090 41.090 50.120 41.260 ;
        RECT 49.170 41.010 50.120 41.090 ;
      LAYER li1 ;
        RECT 50.300 41.010 50.630 42.690 ;
        RECT 51.410 42.650 51.740 42.990 ;
      LAYER li1 ;
        RECT 50.810 41.260 51.760 42.470 ;
        RECT 50.810 41.090 50.840 41.260 ;
        RECT 51.010 41.090 51.200 41.260 ;
        RECT 51.370 41.090 51.560 41.260 ;
        RECT 51.730 41.090 51.760 41.260 ;
        RECT 50.810 41.010 51.760 41.090 ;
        RECT 51.940 41.010 52.190 43.170 ;
        RECT 52.800 43.520 54.100 43.920 ;
        RECT 54.330 44.370 55.280 44.400 ;
        RECT 54.330 44.200 54.360 44.370 ;
        RECT 54.530 44.200 54.720 44.370 ;
        RECT 54.890 44.200 55.080 44.370 ;
        RECT 55.250 44.200 55.280 44.370 ;
        RECT 55.890 44.370 56.840 44.400 ;
        RECT 52.800 42.740 53.130 43.520 ;
        RECT 54.330 43.440 55.280 44.200 ;
      LAYER li1 ;
        RECT 55.460 43.560 55.710 44.270 ;
      LAYER li1 ;
        RECT 55.890 44.200 55.920 44.370 ;
        RECT 56.090 44.200 56.280 44.370 ;
        RECT 56.450 44.200 56.640 44.370 ;
        RECT 56.810 44.200 56.840 44.370 ;
        RECT 57.450 44.370 58.400 44.400 ;
        RECT 55.890 43.740 56.840 44.200 ;
      LAYER li1 ;
        RECT 57.020 43.560 57.270 44.270 ;
        RECT 55.460 43.390 57.270 43.560 ;
      LAYER li1 ;
        RECT 57.450 44.200 57.480 44.370 ;
        RECT 57.650 44.200 57.840 44.370 ;
        RECT 58.010 44.200 58.200 44.370 ;
        RECT 58.370 44.200 58.400 44.370 ;
        RECT 59.210 44.370 60.820 44.400 ;
        RECT 57.450 43.520 58.400 44.200 ;
      LAYER li1 ;
        RECT 55.460 43.220 55.630 43.390 ;
      LAYER li1 ;
        RECT 58.580 43.340 58.910 44.270 ;
        RECT 59.210 44.200 59.260 44.370 ;
        RECT 59.430 44.200 59.700 44.370 ;
        RECT 59.870 44.200 60.140 44.370 ;
        RECT 60.310 44.200 60.550 44.370 ;
        RECT 60.720 44.200 60.820 44.370 ;
        RECT 59.210 43.920 60.820 44.200 ;
        RECT 53.340 42.080 53.670 43.070 ;
      LAYER li1 ;
        RECT 54.370 42.990 55.630 43.220 ;
      LAYER li1 ;
        RECT 57.670 43.210 58.910 43.340 ;
        RECT 55.810 43.170 58.910 43.210 ;
        RECT 55.810 43.040 57.840 43.170 ;
      LAYER li1 ;
        RECT 55.460 42.860 55.630 42.990 ;
        RECT 55.460 42.690 57.350 42.860 ;
      LAYER li1 ;
        RECT 52.570 41.210 54.020 42.080 ;
        RECT 52.570 41.040 52.820 41.210 ;
        RECT 52.990 41.040 53.180 41.210 ;
        RECT 53.350 41.040 53.620 41.210 ;
        RECT 53.790 41.040 54.020 41.210 ;
        RECT 52.570 41.010 54.020 41.040 ;
        RECT 54.330 41.260 55.280 42.590 ;
        RECT 54.330 41.090 54.360 41.260 ;
        RECT 54.530 41.090 54.720 41.260 ;
        RECT 54.890 41.090 55.080 41.260 ;
        RECT 55.250 41.090 55.280 41.260 ;
        RECT 54.330 41.010 55.280 41.090 ;
      LAYER li1 ;
        RECT 55.460 41.010 55.710 42.690 ;
      LAYER li1 ;
        RECT 55.890 41.260 56.840 42.510 ;
        RECT 55.890 41.090 55.920 41.260 ;
        RECT 56.090 41.090 56.280 41.260 ;
        RECT 56.450 41.090 56.640 41.260 ;
        RECT 56.810 41.090 56.840 41.260 ;
        RECT 55.890 41.010 56.840 41.090 ;
      LAYER li1 ;
        RECT 57.020 41.010 57.350 42.690 ;
        RECT 58.130 42.650 58.460 42.990 ;
      LAYER li1 ;
        RECT 57.530 41.260 58.480 42.470 ;
        RECT 57.530 41.090 57.560 41.260 ;
        RECT 57.730 41.090 57.920 41.260 ;
        RECT 58.090 41.090 58.280 41.260 ;
        RECT 58.450 41.090 58.480 41.260 ;
        RECT 57.530 41.010 58.480 41.090 ;
        RECT 58.660 41.010 58.910 43.170 ;
        RECT 59.520 43.520 60.820 43.920 ;
        RECT 61.050 44.370 62.000 44.400 ;
        RECT 61.050 44.200 61.080 44.370 ;
        RECT 61.250 44.200 61.440 44.370 ;
        RECT 61.610 44.200 61.800 44.370 ;
        RECT 61.970 44.200 62.000 44.370 ;
        RECT 62.610 44.370 63.560 44.400 ;
        RECT 59.520 42.740 59.850 43.520 ;
        RECT 61.050 43.440 62.000 44.200 ;
      LAYER li1 ;
        RECT 62.180 43.560 62.430 44.270 ;
      LAYER li1 ;
        RECT 62.610 44.200 62.640 44.370 ;
        RECT 62.810 44.200 63.000 44.370 ;
        RECT 63.170 44.200 63.360 44.370 ;
        RECT 63.530 44.200 63.560 44.370 ;
        RECT 64.170 44.370 65.120 44.400 ;
        RECT 62.610 43.740 63.560 44.200 ;
      LAYER li1 ;
        RECT 63.740 43.560 63.990 44.270 ;
        RECT 62.180 43.390 63.990 43.560 ;
      LAYER li1 ;
        RECT 64.170 44.200 64.200 44.370 ;
        RECT 64.370 44.200 64.560 44.370 ;
        RECT 64.730 44.200 64.920 44.370 ;
        RECT 65.090 44.200 65.120 44.370 ;
        RECT 65.930 44.370 67.540 44.400 ;
        RECT 64.170 43.520 65.120 44.200 ;
      LAYER li1 ;
        RECT 62.180 43.220 62.350 43.390 ;
      LAYER li1 ;
        RECT 65.300 43.340 65.630 44.270 ;
        RECT 65.930 44.200 65.980 44.370 ;
        RECT 66.150 44.200 66.420 44.370 ;
        RECT 66.590 44.200 66.860 44.370 ;
        RECT 67.030 44.200 67.270 44.370 ;
        RECT 67.440 44.200 67.540 44.370 ;
        RECT 65.930 43.920 67.540 44.200 ;
        RECT 60.060 42.080 60.390 43.070 ;
      LAYER li1 ;
        RECT 61.090 42.990 62.350 43.220 ;
      LAYER li1 ;
        RECT 64.390 43.210 65.630 43.340 ;
        RECT 62.530 43.170 65.630 43.210 ;
        RECT 62.530 43.040 64.560 43.170 ;
      LAYER li1 ;
        RECT 62.180 42.860 62.350 42.990 ;
        RECT 62.180 42.690 64.070 42.860 ;
      LAYER li1 ;
        RECT 59.290 41.210 60.740 42.080 ;
        RECT 59.290 41.040 59.540 41.210 ;
        RECT 59.710 41.040 59.900 41.210 ;
        RECT 60.070 41.040 60.340 41.210 ;
        RECT 60.510 41.040 60.740 41.210 ;
        RECT 59.290 41.010 60.740 41.040 ;
        RECT 61.050 41.260 62.000 42.590 ;
        RECT 61.050 41.090 61.080 41.260 ;
        RECT 61.250 41.090 61.440 41.260 ;
        RECT 61.610 41.090 61.800 41.260 ;
        RECT 61.970 41.090 62.000 41.260 ;
        RECT 61.050 41.010 62.000 41.090 ;
      LAYER li1 ;
        RECT 62.180 41.010 62.430 42.690 ;
      LAYER li1 ;
        RECT 62.610 41.260 63.560 42.510 ;
        RECT 62.610 41.090 62.640 41.260 ;
        RECT 62.810 41.090 63.000 41.260 ;
        RECT 63.170 41.090 63.360 41.260 ;
        RECT 63.530 41.090 63.560 41.260 ;
        RECT 62.610 41.010 63.560 41.090 ;
      LAYER li1 ;
        RECT 63.740 41.010 64.070 42.690 ;
        RECT 64.850 42.650 65.180 42.990 ;
      LAYER li1 ;
        RECT 64.250 41.260 65.200 42.470 ;
        RECT 64.250 41.090 64.280 41.260 ;
        RECT 64.450 41.090 64.640 41.260 ;
        RECT 64.810 41.090 65.000 41.260 ;
        RECT 65.170 41.090 65.200 41.260 ;
        RECT 64.250 41.010 65.200 41.090 ;
        RECT 65.380 41.010 65.630 43.170 ;
        RECT 66.240 43.520 67.540 43.920 ;
        RECT 67.770 44.370 68.720 44.400 ;
        RECT 67.770 44.200 67.800 44.370 ;
        RECT 67.970 44.200 68.160 44.370 ;
        RECT 68.330 44.200 68.520 44.370 ;
        RECT 68.690 44.200 68.720 44.370 ;
        RECT 69.330 44.370 70.280 44.400 ;
        RECT 66.240 42.740 66.570 43.520 ;
        RECT 67.770 43.440 68.720 44.200 ;
      LAYER li1 ;
        RECT 68.900 43.560 69.150 44.270 ;
      LAYER li1 ;
        RECT 69.330 44.200 69.360 44.370 ;
        RECT 69.530 44.200 69.720 44.370 ;
        RECT 69.890 44.200 70.080 44.370 ;
        RECT 70.250 44.200 70.280 44.370 ;
        RECT 70.890 44.370 71.840 44.400 ;
        RECT 69.330 43.740 70.280 44.200 ;
      LAYER li1 ;
        RECT 70.460 43.560 70.710 44.270 ;
        RECT 68.900 43.390 70.710 43.560 ;
      LAYER li1 ;
        RECT 70.890 44.200 70.920 44.370 ;
        RECT 71.090 44.200 71.280 44.370 ;
        RECT 71.450 44.200 71.640 44.370 ;
        RECT 71.810 44.200 71.840 44.370 ;
        RECT 72.650 44.370 74.260 44.400 ;
        RECT 70.890 43.520 71.840 44.200 ;
      LAYER li1 ;
        RECT 68.900 43.220 69.070 43.390 ;
      LAYER li1 ;
        RECT 72.020 43.340 72.350 44.270 ;
        RECT 72.650 44.200 72.700 44.370 ;
        RECT 72.870 44.200 73.140 44.370 ;
        RECT 73.310 44.200 73.580 44.370 ;
        RECT 73.750 44.200 73.990 44.370 ;
        RECT 74.160 44.200 74.260 44.370 ;
        RECT 72.650 43.920 74.260 44.200 ;
        RECT 66.780 42.080 67.110 43.070 ;
      LAYER li1 ;
        RECT 67.810 42.990 69.070 43.220 ;
      LAYER li1 ;
        RECT 71.110 43.210 72.350 43.340 ;
        RECT 69.250 43.170 72.350 43.210 ;
        RECT 69.250 43.040 71.280 43.170 ;
      LAYER li1 ;
        RECT 68.900 42.860 69.070 42.990 ;
        RECT 68.900 42.690 70.790 42.860 ;
      LAYER li1 ;
        RECT 66.010 41.210 67.460 42.080 ;
        RECT 66.010 41.040 66.260 41.210 ;
        RECT 66.430 41.040 66.620 41.210 ;
        RECT 66.790 41.040 67.060 41.210 ;
        RECT 67.230 41.040 67.460 41.210 ;
        RECT 66.010 41.010 67.460 41.040 ;
        RECT 67.770 41.260 68.720 42.590 ;
        RECT 67.770 41.090 67.800 41.260 ;
        RECT 67.970 41.090 68.160 41.260 ;
        RECT 68.330 41.090 68.520 41.260 ;
        RECT 68.690 41.090 68.720 41.260 ;
        RECT 67.770 41.010 68.720 41.090 ;
      LAYER li1 ;
        RECT 68.900 41.010 69.150 42.690 ;
      LAYER li1 ;
        RECT 69.330 41.260 70.280 42.510 ;
        RECT 69.330 41.090 69.360 41.260 ;
        RECT 69.530 41.090 69.720 41.260 ;
        RECT 69.890 41.090 70.080 41.260 ;
        RECT 70.250 41.090 70.280 41.260 ;
        RECT 69.330 41.010 70.280 41.090 ;
      LAYER li1 ;
        RECT 70.460 41.010 70.790 42.690 ;
        RECT 71.570 42.650 71.900 42.990 ;
      LAYER li1 ;
        RECT 70.970 41.260 71.920 42.470 ;
        RECT 70.970 41.090 71.000 41.260 ;
        RECT 71.170 41.090 71.360 41.260 ;
        RECT 71.530 41.090 71.720 41.260 ;
        RECT 71.890 41.090 71.920 41.260 ;
        RECT 70.970 41.010 71.920 41.090 ;
        RECT 72.100 41.010 72.350 43.170 ;
        RECT 72.960 43.520 74.260 43.920 ;
        RECT 74.490 44.370 75.440 44.400 ;
        RECT 74.490 44.200 74.520 44.370 ;
        RECT 74.690 44.200 74.880 44.370 ;
        RECT 75.050 44.200 75.240 44.370 ;
        RECT 75.410 44.200 75.440 44.370 ;
        RECT 76.050 44.370 77.000 44.400 ;
        RECT 72.960 42.740 73.290 43.520 ;
        RECT 74.490 43.440 75.440 44.200 ;
      LAYER li1 ;
        RECT 75.620 43.560 75.870 44.270 ;
      LAYER li1 ;
        RECT 76.050 44.200 76.080 44.370 ;
        RECT 76.250 44.200 76.440 44.370 ;
        RECT 76.610 44.200 76.800 44.370 ;
        RECT 76.970 44.200 77.000 44.370 ;
        RECT 77.610 44.370 78.560 44.400 ;
        RECT 76.050 43.740 77.000 44.200 ;
      LAYER li1 ;
        RECT 77.180 43.560 77.430 44.270 ;
        RECT 75.620 43.390 77.430 43.560 ;
      LAYER li1 ;
        RECT 77.610 44.200 77.640 44.370 ;
        RECT 77.810 44.200 78.000 44.370 ;
        RECT 78.170 44.200 78.360 44.370 ;
        RECT 78.530 44.200 78.560 44.370 ;
        RECT 79.370 44.370 80.980 44.400 ;
        RECT 77.610 43.520 78.560 44.200 ;
      LAYER li1 ;
        RECT 75.620 43.220 75.790 43.390 ;
      LAYER li1 ;
        RECT 78.740 43.340 79.070 44.270 ;
        RECT 79.370 44.200 79.420 44.370 ;
        RECT 79.590 44.200 79.860 44.370 ;
        RECT 80.030 44.200 80.300 44.370 ;
        RECT 80.470 44.200 80.710 44.370 ;
        RECT 80.880 44.200 80.980 44.370 ;
        RECT 79.370 43.920 80.980 44.200 ;
        RECT 73.500 42.080 73.830 43.070 ;
      LAYER li1 ;
        RECT 74.530 42.990 75.790 43.220 ;
      LAYER li1 ;
        RECT 77.830 43.210 79.070 43.340 ;
        RECT 75.970 43.170 79.070 43.210 ;
        RECT 75.970 43.040 78.000 43.170 ;
      LAYER li1 ;
        RECT 75.620 42.860 75.790 42.990 ;
        RECT 75.620 42.690 77.510 42.860 ;
      LAYER li1 ;
        RECT 72.730 41.210 74.180 42.080 ;
        RECT 72.730 41.040 72.980 41.210 ;
        RECT 73.150 41.040 73.340 41.210 ;
        RECT 73.510 41.040 73.780 41.210 ;
        RECT 73.950 41.040 74.180 41.210 ;
        RECT 72.730 41.010 74.180 41.040 ;
        RECT 74.490 41.260 75.440 42.590 ;
        RECT 74.490 41.090 74.520 41.260 ;
        RECT 74.690 41.090 74.880 41.260 ;
        RECT 75.050 41.090 75.240 41.260 ;
        RECT 75.410 41.090 75.440 41.260 ;
        RECT 74.490 41.010 75.440 41.090 ;
      LAYER li1 ;
        RECT 75.620 41.010 75.870 42.690 ;
      LAYER li1 ;
        RECT 76.050 41.260 77.000 42.510 ;
        RECT 76.050 41.090 76.080 41.260 ;
        RECT 76.250 41.090 76.440 41.260 ;
        RECT 76.610 41.090 76.800 41.260 ;
        RECT 76.970 41.090 77.000 41.260 ;
        RECT 76.050 41.010 77.000 41.090 ;
      LAYER li1 ;
        RECT 77.180 41.010 77.510 42.690 ;
        RECT 78.290 42.650 78.620 42.990 ;
      LAYER li1 ;
        RECT 77.690 41.260 78.640 42.470 ;
        RECT 77.690 41.090 77.720 41.260 ;
        RECT 77.890 41.090 78.080 41.260 ;
        RECT 78.250 41.090 78.440 41.260 ;
        RECT 78.610 41.090 78.640 41.260 ;
        RECT 77.690 41.010 78.640 41.090 ;
        RECT 78.820 41.010 79.070 43.170 ;
        RECT 79.680 43.520 80.980 43.920 ;
        RECT 81.210 44.370 82.160 44.400 ;
        RECT 81.210 44.200 81.240 44.370 ;
        RECT 81.410 44.200 81.600 44.370 ;
        RECT 81.770 44.200 81.960 44.370 ;
        RECT 82.130 44.200 82.160 44.370 ;
        RECT 82.770 44.370 83.720 44.400 ;
        RECT 79.680 42.740 80.010 43.520 ;
        RECT 81.210 43.440 82.160 44.200 ;
      LAYER li1 ;
        RECT 82.340 43.560 82.590 44.270 ;
      LAYER li1 ;
        RECT 82.770 44.200 82.800 44.370 ;
        RECT 82.970 44.200 83.160 44.370 ;
        RECT 83.330 44.200 83.520 44.370 ;
        RECT 83.690 44.200 83.720 44.370 ;
        RECT 84.330 44.370 85.280 44.400 ;
        RECT 82.770 43.740 83.720 44.200 ;
      LAYER li1 ;
        RECT 83.900 43.560 84.150 44.270 ;
        RECT 82.340 43.390 84.150 43.560 ;
      LAYER li1 ;
        RECT 84.330 44.200 84.360 44.370 ;
        RECT 84.530 44.200 84.720 44.370 ;
        RECT 84.890 44.200 85.080 44.370 ;
        RECT 85.250 44.200 85.280 44.370 ;
        RECT 86.090 44.370 87.700 44.400 ;
        RECT 84.330 43.520 85.280 44.200 ;
      LAYER li1 ;
        RECT 82.340 43.220 82.510 43.390 ;
      LAYER li1 ;
        RECT 85.460 43.340 85.790 44.270 ;
        RECT 86.090 44.200 86.140 44.370 ;
        RECT 86.310 44.200 86.580 44.370 ;
        RECT 86.750 44.200 87.020 44.370 ;
        RECT 87.190 44.200 87.430 44.370 ;
        RECT 87.600 44.200 87.700 44.370 ;
        RECT 86.090 43.920 87.700 44.200 ;
        RECT 80.220 42.080 80.550 43.070 ;
      LAYER li1 ;
        RECT 81.250 42.990 82.510 43.220 ;
      LAYER li1 ;
        RECT 84.550 43.210 85.790 43.340 ;
        RECT 82.690 43.170 85.790 43.210 ;
        RECT 82.690 43.040 84.720 43.170 ;
      LAYER li1 ;
        RECT 82.340 42.860 82.510 42.990 ;
        RECT 82.340 42.690 84.230 42.860 ;
      LAYER li1 ;
        RECT 79.450 41.210 80.900 42.080 ;
        RECT 79.450 41.040 79.700 41.210 ;
        RECT 79.870 41.040 80.060 41.210 ;
        RECT 80.230 41.040 80.500 41.210 ;
        RECT 80.670 41.040 80.900 41.210 ;
        RECT 79.450 41.010 80.900 41.040 ;
        RECT 81.210 41.260 82.160 42.590 ;
        RECT 81.210 41.090 81.240 41.260 ;
        RECT 81.410 41.090 81.600 41.260 ;
        RECT 81.770 41.090 81.960 41.260 ;
        RECT 82.130 41.090 82.160 41.260 ;
        RECT 81.210 41.010 82.160 41.090 ;
      LAYER li1 ;
        RECT 82.340 41.010 82.590 42.690 ;
      LAYER li1 ;
        RECT 82.770 41.260 83.720 42.510 ;
        RECT 82.770 41.090 82.800 41.260 ;
        RECT 82.970 41.090 83.160 41.260 ;
        RECT 83.330 41.090 83.520 41.260 ;
        RECT 83.690 41.090 83.720 41.260 ;
        RECT 82.770 41.010 83.720 41.090 ;
      LAYER li1 ;
        RECT 83.900 41.010 84.230 42.690 ;
        RECT 85.010 42.650 85.340 42.990 ;
      LAYER li1 ;
        RECT 84.410 41.260 85.360 42.470 ;
        RECT 84.410 41.090 84.440 41.260 ;
        RECT 84.610 41.090 84.800 41.260 ;
        RECT 84.970 41.090 85.160 41.260 ;
        RECT 85.330 41.090 85.360 41.260 ;
        RECT 84.410 41.010 85.360 41.090 ;
        RECT 85.540 41.010 85.790 43.170 ;
        RECT 86.400 43.520 87.700 43.920 ;
        RECT 87.930 44.370 88.880 44.400 ;
        RECT 87.930 44.200 87.960 44.370 ;
        RECT 88.130 44.200 88.320 44.370 ;
        RECT 88.490 44.200 88.680 44.370 ;
        RECT 88.850 44.200 88.880 44.370 ;
        RECT 89.490 44.370 90.440 44.400 ;
        RECT 86.400 42.740 86.730 43.520 ;
        RECT 87.930 43.440 88.880 44.200 ;
      LAYER li1 ;
        RECT 89.060 43.560 89.310 44.270 ;
      LAYER li1 ;
        RECT 89.490 44.200 89.520 44.370 ;
        RECT 89.690 44.200 89.880 44.370 ;
        RECT 90.050 44.200 90.240 44.370 ;
        RECT 90.410 44.200 90.440 44.370 ;
        RECT 91.050 44.370 92.000 44.400 ;
        RECT 89.490 43.740 90.440 44.200 ;
      LAYER li1 ;
        RECT 90.620 43.560 90.870 44.270 ;
        RECT 89.060 43.390 90.870 43.560 ;
      LAYER li1 ;
        RECT 91.050 44.200 91.080 44.370 ;
        RECT 91.250 44.200 91.440 44.370 ;
        RECT 91.610 44.200 91.800 44.370 ;
        RECT 91.970 44.200 92.000 44.370 ;
        RECT 92.810 44.370 94.420 44.400 ;
        RECT 91.050 43.520 92.000 44.200 ;
      LAYER li1 ;
        RECT 89.060 43.220 89.230 43.390 ;
      LAYER li1 ;
        RECT 92.180 43.340 92.510 44.270 ;
        RECT 92.810 44.200 92.860 44.370 ;
        RECT 93.030 44.200 93.300 44.370 ;
        RECT 93.470 44.200 93.740 44.370 ;
        RECT 93.910 44.200 94.150 44.370 ;
        RECT 94.320 44.200 94.420 44.370 ;
        RECT 92.810 43.920 94.420 44.200 ;
        RECT 86.940 42.080 87.270 43.070 ;
      LAYER li1 ;
        RECT 87.970 42.990 89.230 43.220 ;
      LAYER li1 ;
        RECT 91.270 43.210 92.510 43.340 ;
        RECT 89.410 43.170 92.510 43.210 ;
        RECT 89.410 43.040 91.440 43.170 ;
      LAYER li1 ;
        RECT 89.060 42.860 89.230 42.990 ;
        RECT 89.060 42.690 90.950 42.860 ;
      LAYER li1 ;
        RECT 86.170 41.210 87.620 42.080 ;
        RECT 86.170 41.040 86.420 41.210 ;
        RECT 86.590 41.040 86.780 41.210 ;
        RECT 86.950 41.040 87.220 41.210 ;
        RECT 87.390 41.040 87.620 41.210 ;
        RECT 86.170 41.010 87.620 41.040 ;
        RECT 87.930 41.260 88.880 42.590 ;
        RECT 87.930 41.090 87.960 41.260 ;
        RECT 88.130 41.090 88.320 41.260 ;
        RECT 88.490 41.090 88.680 41.260 ;
        RECT 88.850 41.090 88.880 41.260 ;
        RECT 87.930 41.010 88.880 41.090 ;
      LAYER li1 ;
        RECT 89.060 41.010 89.310 42.690 ;
      LAYER li1 ;
        RECT 89.490 41.260 90.440 42.510 ;
        RECT 89.490 41.090 89.520 41.260 ;
        RECT 89.690 41.090 89.880 41.260 ;
        RECT 90.050 41.090 90.240 41.260 ;
        RECT 90.410 41.090 90.440 41.260 ;
        RECT 89.490 41.010 90.440 41.090 ;
      LAYER li1 ;
        RECT 90.620 41.010 90.950 42.690 ;
        RECT 91.730 42.650 92.060 42.990 ;
      LAYER li1 ;
        RECT 91.130 41.260 92.080 42.470 ;
        RECT 91.130 41.090 91.160 41.260 ;
        RECT 91.330 41.090 91.520 41.260 ;
        RECT 91.690 41.090 91.880 41.260 ;
        RECT 92.050 41.090 92.080 41.260 ;
        RECT 91.130 41.010 92.080 41.090 ;
        RECT 92.260 41.010 92.510 43.170 ;
        RECT 93.120 43.520 94.420 43.920 ;
        RECT 94.720 44.330 96.530 44.500 ;
        RECT 93.120 42.740 93.450 43.520 ;
        RECT 94.720 43.410 95.050 44.330 ;
      LAYER li1 ;
        RECT 95.300 43.410 95.830 44.150 ;
      LAYER li1 ;
        RECT 93.660 42.080 93.990 43.070 ;
      LAYER li1 ;
        RECT 94.690 42.900 95.110 43.230 ;
        RECT 95.300 42.840 95.470 43.410 ;
      LAYER li1 ;
        RECT 96.360 43.310 96.530 44.330 ;
        RECT 96.710 44.370 97.810 44.400 ;
        RECT 96.710 44.200 96.760 44.370 ;
        RECT 96.930 44.200 97.120 44.370 ;
        RECT 97.290 44.200 97.480 44.370 ;
        RECT 97.650 44.200 97.810 44.370 ;
        RECT 98.570 44.370 100.180 44.400 ;
        RECT 96.710 43.490 97.810 44.200 ;
        RECT 97.980 43.310 98.230 44.240 ;
        RECT 98.570 44.200 98.620 44.370 ;
        RECT 98.790 44.200 99.060 44.370 ;
        RECT 99.230 44.200 99.500 44.370 ;
        RECT 99.670 44.200 99.910 44.370 ;
        RECT 100.080 44.200 100.180 44.370 ;
        RECT 98.570 43.920 100.180 44.200 ;
      LAYER li1 ;
        RECT 95.650 43.020 96.160 43.230 ;
      LAYER li1 ;
        RECT 96.360 43.140 98.230 43.310 ;
        RECT 98.880 43.520 100.180 43.920 ;
        RECT 101.370 44.370 102.320 44.400 ;
        RECT 101.370 44.200 101.400 44.370 ;
        RECT 101.570 44.200 101.760 44.370 ;
        RECT 101.930 44.200 102.120 44.370 ;
        RECT 102.290 44.200 102.320 44.370 ;
        RECT 102.930 44.370 103.880 44.400 ;
      LAYER li1 ;
        RECT 95.300 42.670 96.360 42.840 ;
        RECT 96.090 42.590 96.360 42.670 ;
        RECT 96.810 42.650 97.320 42.960 ;
        RECT 97.570 42.650 98.280 42.960 ;
      LAYER li1 ;
        RECT 98.880 42.740 99.210 43.520 ;
        RECT 101.370 43.440 102.320 44.200 ;
      LAYER li1 ;
        RECT 102.500 43.560 102.750 44.270 ;
      LAYER li1 ;
        RECT 102.930 44.200 102.960 44.370 ;
        RECT 103.130 44.200 103.320 44.370 ;
        RECT 103.490 44.200 103.680 44.370 ;
        RECT 103.850 44.200 103.880 44.370 ;
        RECT 104.490 44.370 105.440 44.400 ;
        RECT 102.930 43.740 103.880 44.200 ;
      LAYER li1 ;
        RECT 104.060 43.560 104.310 44.270 ;
        RECT 102.500 43.390 104.310 43.560 ;
      LAYER li1 ;
        RECT 104.490 44.200 104.520 44.370 ;
        RECT 104.690 44.200 104.880 44.370 ;
        RECT 105.050 44.200 105.240 44.370 ;
        RECT 105.410 44.200 105.440 44.370 ;
        RECT 106.250 44.370 107.860 44.400 ;
        RECT 104.490 43.520 105.440 44.200 ;
      LAYER li1 ;
        RECT 102.500 43.220 102.670 43.390 ;
      LAYER li1 ;
        RECT 105.620 43.340 105.950 44.270 ;
        RECT 106.250 44.200 106.300 44.370 ;
        RECT 106.470 44.200 106.740 44.370 ;
        RECT 106.910 44.200 107.180 44.370 ;
        RECT 107.350 44.200 107.590 44.370 ;
        RECT 107.760 44.200 107.860 44.370 ;
        RECT 106.250 43.920 107.860 44.200 ;
        RECT 92.890 41.210 94.340 42.080 ;
        RECT 92.890 41.040 93.140 41.210 ;
        RECT 93.310 41.040 93.500 41.210 ;
        RECT 93.670 41.040 93.940 41.210 ;
        RECT 94.110 41.040 94.340 41.210 ;
        RECT 92.890 41.010 94.340 41.040 ;
        RECT 94.650 41.260 95.910 42.490 ;
      LAYER li1 ;
        RECT 96.090 41.510 96.610 42.590 ;
      LAYER li1 ;
        RECT 94.650 41.090 94.660 41.260 ;
        RECT 94.830 41.090 95.020 41.260 ;
        RECT 95.190 41.090 95.380 41.260 ;
        RECT 95.550 41.090 95.740 41.260 ;
        RECT 94.650 41.010 95.910 41.090 ;
      LAYER li1 ;
        RECT 96.440 41.010 96.610 41.510 ;
      LAYER li1 ;
        RECT 96.870 41.260 98.180 42.470 ;
        RECT 99.420 42.080 99.750 43.070 ;
      LAYER li1 ;
        RECT 101.410 42.990 102.670 43.220 ;
      LAYER li1 ;
        RECT 104.710 43.210 105.950 43.340 ;
        RECT 102.850 43.170 105.950 43.210 ;
        RECT 102.850 43.040 104.880 43.170 ;
      LAYER li1 ;
        RECT 102.500 42.860 102.670 42.990 ;
        RECT 102.500 42.690 104.390 42.860 ;
      LAYER li1 ;
        RECT 96.870 41.090 96.900 41.260 ;
        RECT 97.070 41.090 97.260 41.260 ;
        RECT 97.430 41.090 97.620 41.260 ;
        RECT 97.790 41.090 97.980 41.260 ;
        RECT 98.150 41.090 98.180 41.260 ;
        RECT 96.870 41.010 98.180 41.090 ;
        RECT 98.650 41.210 100.100 42.080 ;
      LAYER li1 ;
        RECT 100.470 41.540 100.640 42.450 ;
      LAYER li1 ;
        RECT 98.650 41.040 98.900 41.210 ;
        RECT 99.070 41.040 99.260 41.210 ;
        RECT 99.430 41.040 99.700 41.210 ;
        RECT 99.870 41.040 100.100 41.210 ;
        RECT 98.650 41.010 100.100 41.040 ;
        RECT 101.370 41.260 102.320 42.590 ;
        RECT 101.370 41.090 101.400 41.260 ;
        RECT 101.570 41.090 101.760 41.260 ;
        RECT 101.930 41.090 102.120 41.260 ;
        RECT 102.290 41.090 102.320 41.260 ;
        RECT 101.370 41.010 102.320 41.090 ;
      LAYER li1 ;
        RECT 102.500 41.010 102.750 42.690 ;
      LAYER li1 ;
        RECT 102.930 41.260 103.880 42.510 ;
        RECT 102.930 41.090 102.960 41.260 ;
        RECT 103.130 41.090 103.320 41.260 ;
        RECT 103.490 41.090 103.680 41.260 ;
        RECT 103.850 41.090 103.880 41.260 ;
        RECT 102.930 41.010 103.880 41.090 ;
      LAYER li1 ;
        RECT 104.060 41.010 104.390 42.690 ;
        RECT 105.170 42.650 105.500 42.990 ;
      LAYER li1 ;
        RECT 104.570 41.260 105.520 42.470 ;
        RECT 104.570 41.090 104.600 41.260 ;
        RECT 104.770 41.090 104.960 41.260 ;
        RECT 105.130 41.090 105.320 41.260 ;
        RECT 105.490 41.090 105.520 41.260 ;
        RECT 104.570 41.010 105.520 41.090 ;
        RECT 105.700 41.010 105.950 43.170 ;
        RECT 106.560 43.520 107.860 43.920 ;
        RECT 108.090 44.370 109.040 44.400 ;
        RECT 108.090 44.200 108.120 44.370 ;
        RECT 108.290 44.200 108.480 44.370 ;
        RECT 108.650 44.200 108.840 44.370 ;
        RECT 109.010 44.200 109.040 44.370 ;
        RECT 109.650 44.370 110.600 44.400 ;
        RECT 106.560 42.740 106.890 43.520 ;
        RECT 108.090 43.440 109.040 44.200 ;
      LAYER li1 ;
        RECT 109.220 43.560 109.470 44.270 ;
      LAYER li1 ;
        RECT 109.650 44.200 109.680 44.370 ;
        RECT 109.850 44.200 110.040 44.370 ;
        RECT 110.210 44.200 110.400 44.370 ;
        RECT 110.570 44.200 110.600 44.370 ;
        RECT 111.210 44.370 112.160 44.400 ;
        RECT 109.650 43.740 110.600 44.200 ;
      LAYER li1 ;
        RECT 110.780 43.560 111.030 44.270 ;
        RECT 109.220 43.390 111.030 43.560 ;
      LAYER li1 ;
        RECT 111.210 44.200 111.240 44.370 ;
        RECT 111.410 44.200 111.600 44.370 ;
        RECT 111.770 44.200 111.960 44.370 ;
        RECT 112.130 44.200 112.160 44.370 ;
        RECT 112.970 44.370 114.580 44.400 ;
        RECT 111.210 43.520 112.160 44.200 ;
      LAYER li1 ;
        RECT 109.220 43.220 109.390 43.390 ;
      LAYER li1 ;
        RECT 112.340 43.340 112.670 44.270 ;
        RECT 112.970 44.200 113.020 44.370 ;
        RECT 113.190 44.200 113.460 44.370 ;
        RECT 113.630 44.200 113.900 44.370 ;
        RECT 114.070 44.200 114.310 44.370 ;
        RECT 114.480 44.200 114.580 44.370 ;
        RECT 112.970 43.920 114.580 44.200 ;
        RECT 107.100 42.080 107.430 43.070 ;
      LAYER li1 ;
        RECT 108.130 42.990 109.390 43.220 ;
      LAYER li1 ;
        RECT 111.430 43.210 112.670 43.340 ;
        RECT 109.570 43.170 112.670 43.210 ;
        RECT 109.570 43.040 111.600 43.170 ;
      LAYER li1 ;
        RECT 109.220 42.860 109.390 42.990 ;
        RECT 109.220 42.690 111.110 42.860 ;
      LAYER li1 ;
        RECT 106.330 41.210 107.780 42.080 ;
        RECT 106.330 41.040 106.580 41.210 ;
        RECT 106.750 41.040 106.940 41.210 ;
        RECT 107.110 41.040 107.380 41.210 ;
        RECT 107.550 41.040 107.780 41.210 ;
        RECT 106.330 41.010 107.780 41.040 ;
        RECT 108.090 41.260 109.040 42.590 ;
        RECT 108.090 41.090 108.120 41.260 ;
        RECT 108.290 41.090 108.480 41.260 ;
        RECT 108.650 41.090 108.840 41.260 ;
        RECT 109.010 41.090 109.040 41.260 ;
        RECT 108.090 41.010 109.040 41.090 ;
      LAYER li1 ;
        RECT 109.220 41.010 109.470 42.690 ;
      LAYER li1 ;
        RECT 109.650 41.260 110.600 42.510 ;
        RECT 109.650 41.090 109.680 41.260 ;
        RECT 109.850 41.090 110.040 41.260 ;
        RECT 110.210 41.090 110.400 41.260 ;
        RECT 110.570 41.090 110.600 41.260 ;
        RECT 109.650 41.010 110.600 41.090 ;
      LAYER li1 ;
        RECT 110.780 41.010 111.110 42.690 ;
        RECT 111.890 42.650 112.220 42.990 ;
      LAYER li1 ;
        RECT 111.290 41.260 112.240 42.470 ;
        RECT 111.290 41.090 111.320 41.260 ;
        RECT 111.490 41.090 111.680 41.260 ;
        RECT 111.850 41.090 112.040 41.260 ;
        RECT 112.210 41.090 112.240 41.260 ;
        RECT 111.290 41.010 112.240 41.090 ;
        RECT 112.420 41.010 112.670 43.170 ;
        RECT 113.280 43.520 114.580 43.920 ;
        RECT 116.250 44.370 117.200 44.400 ;
        RECT 116.250 44.200 116.280 44.370 ;
        RECT 116.450 44.200 116.640 44.370 ;
        RECT 116.810 44.200 117.000 44.370 ;
        RECT 117.170 44.200 117.200 44.370 ;
        RECT 117.810 44.370 118.760 44.400 ;
        RECT 113.280 42.740 113.610 43.520 ;
        RECT 116.250 43.440 117.200 44.200 ;
      LAYER li1 ;
        RECT 117.380 43.560 117.630 44.270 ;
      LAYER li1 ;
        RECT 117.810 44.200 117.840 44.370 ;
        RECT 118.010 44.200 118.200 44.370 ;
        RECT 118.370 44.200 118.560 44.370 ;
        RECT 118.730 44.200 118.760 44.370 ;
        RECT 119.370 44.370 120.320 44.400 ;
        RECT 117.810 43.740 118.760 44.200 ;
      LAYER li1 ;
        RECT 118.940 43.560 119.190 44.270 ;
        RECT 117.380 43.390 119.190 43.560 ;
      LAYER li1 ;
        RECT 119.370 44.200 119.400 44.370 ;
        RECT 119.570 44.200 119.760 44.370 ;
        RECT 119.930 44.200 120.120 44.370 ;
        RECT 120.290 44.200 120.320 44.370 ;
        RECT 121.130 44.370 122.740 44.400 ;
        RECT 119.370 43.520 120.320 44.200 ;
      LAYER li1 ;
        RECT 117.380 43.220 117.550 43.390 ;
      LAYER li1 ;
        RECT 120.500 43.340 120.830 44.270 ;
        RECT 121.130 44.200 121.180 44.370 ;
        RECT 121.350 44.200 121.620 44.370 ;
        RECT 121.790 44.200 122.060 44.370 ;
        RECT 122.230 44.200 122.470 44.370 ;
        RECT 122.640 44.200 122.740 44.370 ;
        RECT 121.130 43.920 122.740 44.200 ;
        RECT 113.820 42.080 114.150 43.070 ;
      LAYER li1 ;
        RECT 116.290 42.990 117.550 43.220 ;
      LAYER li1 ;
        RECT 119.590 43.210 120.830 43.340 ;
        RECT 117.730 43.170 120.830 43.210 ;
        RECT 117.730 43.040 119.760 43.170 ;
      LAYER li1 ;
        RECT 117.380 42.860 117.550 42.990 ;
        RECT 117.380 42.690 119.270 42.860 ;
      LAYER li1 ;
        RECT 113.050 41.210 114.500 42.080 ;
        RECT 113.050 41.040 113.300 41.210 ;
        RECT 113.470 41.040 113.660 41.210 ;
        RECT 113.830 41.040 114.100 41.210 ;
        RECT 114.270 41.040 114.500 41.210 ;
        RECT 113.050 41.010 114.500 41.040 ;
        RECT 116.250 41.260 117.200 42.590 ;
        RECT 116.250 41.090 116.280 41.260 ;
        RECT 116.450 41.090 116.640 41.260 ;
        RECT 116.810 41.090 117.000 41.260 ;
        RECT 117.170 41.090 117.200 41.260 ;
        RECT 116.250 41.010 117.200 41.090 ;
      LAYER li1 ;
        RECT 117.380 41.010 117.630 42.690 ;
      LAYER li1 ;
        RECT 117.810 41.260 118.760 42.510 ;
        RECT 117.810 41.090 117.840 41.260 ;
        RECT 118.010 41.090 118.200 41.260 ;
        RECT 118.370 41.090 118.560 41.260 ;
        RECT 118.730 41.090 118.760 41.260 ;
        RECT 117.810 41.010 118.760 41.090 ;
      LAYER li1 ;
        RECT 118.940 41.010 119.270 42.690 ;
        RECT 120.050 42.650 120.380 42.990 ;
      LAYER li1 ;
        RECT 119.450 41.260 120.400 42.470 ;
        RECT 119.450 41.090 119.480 41.260 ;
        RECT 119.650 41.090 119.840 41.260 ;
        RECT 120.010 41.090 120.200 41.260 ;
        RECT 120.370 41.090 120.400 41.260 ;
        RECT 119.450 41.010 120.400 41.090 ;
        RECT 120.580 41.010 120.830 43.170 ;
        RECT 121.440 43.520 122.740 43.920 ;
        RECT 122.970 44.370 123.920 44.400 ;
        RECT 122.970 44.200 123.000 44.370 ;
        RECT 123.170 44.200 123.360 44.370 ;
        RECT 123.530 44.200 123.720 44.370 ;
        RECT 123.890 44.200 123.920 44.370 ;
        RECT 124.530 44.370 125.480 44.400 ;
        RECT 121.440 42.740 121.770 43.520 ;
        RECT 122.970 43.440 123.920 44.200 ;
      LAYER li1 ;
        RECT 124.100 43.560 124.350 44.270 ;
      LAYER li1 ;
        RECT 124.530 44.200 124.560 44.370 ;
        RECT 124.730 44.200 124.920 44.370 ;
        RECT 125.090 44.200 125.280 44.370 ;
        RECT 125.450 44.200 125.480 44.370 ;
        RECT 126.090 44.370 127.040 44.400 ;
        RECT 124.530 43.740 125.480 44.200 ;
      LAYER li1 ;
        RECT 125.660 43.560 125.910 44.270 ;
        RECT 124.100 43.390 125.910 43.560 ;
      LAYER li1 ;
        RECT 126.090 44.200 126.120 44.370 ;
        RECT 126.290 44.200 126.480 44.370 ;
        RECT 126.650 44.200 126.840 44.370 ;
        RECT 127.010 44.200 127.040 44.370 ;
        RECT 127.850 44.370 129.460 44.400 ;
        RECT 126.090 43.520 127.040 44.200 ;
      LAYER li1 ;
        RECT 124.100 43.220 124.270 43.390 ;
      LAYER li1 ;
        RECT 127.220 43.340 127.550 44.270 ;
        RECT 127.850 44.200 127.900 44.370 ;
        RECT 128.070 44.200 128.340 44.370 ;
        RECT 128.510 44.200 128.780 44.370 ;
        RECT 128.950 44.200 129.190 44.370 ;
        RECT 129.360 44.200 129.460 44.370 ;
        RECT 127.850 43.920 129.460 44.200 ;
        RECT 121.980 42.080 122.310 43.070 ;
      LAYER li1 ;
        RECT 123.010 42.990 124.270 43.220 ;
      LAYER li1 ;
        RECT 126.310 43.210 127.550 43.340 ;
        RECT 124.450 43.170 127.550 43.210 ;
        RECT 124.450 43.040 126.480 43.170 ;
      LAYER li1 ;
        RECT 124.100 42.860 124.270 42.990 ;
        RECT 124.100 42.690 125.990 42.860 ;
      LAYER li1 ;
        RECT 121.210 41.210 122.660 42.080 ;
        RECT 121.210 41.040 121.460 41.210 ;
        RECT 121.630 41.040 121.820 41.210 ;
        RECT 121.990 41.040 122.260 41.210 ;
        RECT 122.430 41.040 122.660 41.210 ;
        RECT 121.210 41.010 122.660 41.040 ;
        RECT 122.970 41.260 123.920 42.590 ;
        RECT 122.970 41.090 123.000 41.260 ;
        RECT 123.170 41.090 123.360 41.260 ;
        RECT 123.530 41.090 123.720 41.260 ;
        RECT 123.890 41.090 123.920 41.260 ;
        RECT 122.970 41.010 123.920 41.090 ;
      LAYER li1 ;
        RECT 124.100 41.010 124.350 42.690 ;
      LAYER li1 ;
        RECT 124.530 41.260 125.480 42.510 ;
        RECT 124.530 41.090 124.560 41.260 ;
        RECT 124.730 41.090 124.920 41.260 ;
        RECT 125.090 41.090 125.280 41.260 ;
        RECT 125.450 41.090 125.480 41.260 ;
        RECT 124.530 41.010 125.480 41.090 ;
      LAYER li1 ;
        RECT 125.660 41.010 125.990 42.690 ;
        RECT 126.770 42.650 127.100 42.990 ;
      LAYER li1 ;
        RECT 126.170 41.260 127.120 42.470 ;
        RECT 126.170 41.090 126.200 41.260 ;
        RECT 126.370 41.090 126.560 41.260 ;
        RECT 126.730 41.090 126.920 41.260 ;
        RECT 127.090 41.090 127.120 41.260 ;
        RECT 126.170 41.010 127.120 41.090 ;
        RECT 127.300 41.010 127.550 43.170 ;
        RECT 128.160 43.520 129.460 43.920 ;
        RECT 129.690 44.370 130.640 44.400 ;
        RECT 129.690 44.200 129.720 44.370 ;
        RECT 129.890 44.200 130.080 44.370 ;
        RECT 130.250 44.200 130.440 44.370 ;
        RECT 130.610 44.200 130.640 44.370 ;
        RECT 131.250 44.370 132.200 44.400 ;
        RECT 128.160 42.740 128.490 43.520 ;
        RECT 129.690 43.440 130.640 44.200 ;
      LAYER li1 ;
        RECT 130.820 43.560 131.070 44.270 ;
      LAYER li1 ;
        RECT 131.250 44.200 131.280 44.370 ;
        RECT 131.450 44.200 131.640 44.370 ;
        RECT 131.810 44.200 132.000 44.370 ;
        RECT 132.170 44.200 132.200 44.370 ;
        RECT 132.810 44.370 133.760 44.400 ;
        RECT 131.250 43.740 132.200 44.200 ;
      LAYER li1 ;
        RECT 132.380 43.560 132.630 44.270 ;
        RECT 130.820 43.390 132.630 43.560 ;
      LAYER li1 ;
        RECT 132.810 44.200 132.840 44.370 ;
        RECT 133.010 44.200 133.200 44.370 ;
        RECT 133.370 44.200 133.560 44.370 ;
        RECT 133.730 44.200 133.760 44.370 ;
        RECT 134.570 44.370 136.180 44.400 ;
        RECT 132.810 43.520 133.760 44.200 ;
      LAYER li1 ;
        RECT 130.820 43.220 130.990 43.390 ;
      LAYER li1 ;
        RECT 133.940 43.340 134.270 44.270 ;
        RECT 134.570 44.200 134.620 44.370 ;
        RECT 134.790 44.200 135.060 44.370 ;
        RECT 135.230 44.200 135.500 44.370 ;
        RECT 135.670 44.200 135.910 44.370 ;
        RECT 136.080 44.200 136.180 44.370 ;
        RECT 134.570 43.920 136.180 44.200 ;
        RECT 128.700 42.080 129.030 43.070 ;
      LAYER li1 ;
        RECT 129.730 42.990 130.990 43.220 ;
      LAYER li1 ;
        RECT 133.030 43.210 134.270 43.340 ;
        RECT 131.170 43.170 134.270 43.210 ;
        RECT 131.170 43.040 133.200 43.170 ;
      LAYER li1 ;
        RECT 130.820 42.860 130.990 42.990 ;
        RECT 130.820 42.690 132.710 42.860 ;
      LAYER li1 ;
        RECT 127.930 41.210 129.380 42.080 ;
        RECT 127.930 41.040 128.180 41.210 ;
        RECT 128.350 41.040 128.540 41.210 ;
        RECT 128.710 41.040 128.980 41.210 ;
        RECT 129.150 41.040 129.380 41.210 ;
        RECT 127.930 41.010 129.380 41.040 ;
        RECT 129.690 41.260 130.640 42.590 ;
        RECT 129.690 41.090 129.720 41.260 ;
        RECT 129.890 41.090 130.080 41.260 ;
        RECT 130.250 41.090 130.440 41.260 ;
        RECT 130.610 41.090 130.640 41.260 ;
        RECT 129.690 41.010 130.640 41.090 ;
      LAYER li1 ;
        RECT 130.820 41.010 131.070 42.690 ;
      LAYER li1 ;
        RECT 131.250 41.260 132.200 42.510 ;
        RECT 131.250 41.090 131.280 41.260 ;
        RECT 131.450 41.090 131.640 41.260 ;
        RECT 131.810 41.090 132.000 41.260 ;
        RECT 132.170 41.090 132.200 41.260 ;
        RECT 131.250 41.010 132.200 41.090 ;
      LAYER li1 ;
        RECT 132.380 41.010 132.710 42.690 ;
        RECT 133.490 42.650 133.820 42.990 ;
      LAYER li1 ;
        RECT 132.890 41.260 133.840 42.470 ;
        RECT 132.890 41.090 132.920 41.260 ;
        RECT 133.090 41.090 133.280 41.260 ;
        RECT 133.450 41.090 133.640 41.260 ;
        RECT 133.810 41.090 133.840 41.260 ;
        RECT 132.890 41.010 133.840 41.090 ;
        RECT 134.020 41.010 134.270 43.170 ;
        RECT 134.880 43.520 136.180 43.920 ;
        RECT 136.650 44.370 138.360 44.400 ;
        RECT 136.650 44.200 136.700 44.370 ;
        RECT 136.870 44.200 137.060 44.370 ;
        RECT 137.230 44.200 137.420 44.370 ;
        RECT 137.590 44.200 137.780 44.370 ;
        RECT 137.950 44.200 138.140 44.370 ;
        RECT 138.310 44.200 138.360 44.370 ;
        RECT 139.000 44.370 139.590 44.400 ;
        RECT 134.880 42.740 135.210 43.520 ;
        RECT 136.650 43.440 138.360 44.200 ;
      LAYER li1 ;
        RECT 138.540 43.310 138.790 44.270 ;
      LAYER li1 ;
        RECT 139.000 44.200 139.030 44.370 ;
        RECT 139.200 44.200 139.390 44.370 ;
        RECT 139.560 44.200 139.590 44.370 ;
        RECT 139.000 43.490 139.590 44.200 ;
        RECT 139.850 44.370 141.460 44.400 ;
        RECT 139.850 44.200 139.900 44.370 ;
        RECT 140.070 44.200 140.340 44.370 ;
        RECT 140.510 44.200 140.780 44.370 ;
        RECT 140.950 44.200 141.190 44.370 ;
        RECT 141.360 44.200 141.460 44.370 ;
        RECT 139.850 43.920 141.460 44.200 ;
        RECT 140.160 43.520 141.460 43.920 ;
        RECT 135.420 42.080 135.750 43.070 ;
      LAYER li1 ;
        RECT 136.450 43.020 137.640 43.260 ;
        RECT 137.890 43.020 138.240 43.260 ;
        RECT 138.540 43.140 139.560 43.310 ;
      LAYER li1 ;
        RECT 136.580 42.670 138.610 42.840 ;
        RECT 134.650 41.210 136.100 42.080 ;
        RECT 134.650 41.040 134.900 41.210 ;
        RECT 135.070 41.040 135.260 41.210 ;
        RECT 135.430 41.040 135.700 41.210 ;
        RECT 135.870 41.040 136.100 41.210 ;
        RECT 134.650 41.010 136.100 41.040 ;
        RECT 136.580 41.010 136.830 42.670 ;
        RECT 137.010 41.260 138.260 42.490 ;
        RECT 137.180 41.090 137.370 41.260 ;
        RECT 137.540 41.090 137.730 41.260 ;
        RECT 137.900 41.090 138.090 41.260 ;
        RECT 137.010 41.010 138.260 41.090 ;
        RECT 138.440 41.010 138.610 42.670 ;
      LAYER li1 ;
        RECT 138.790 41.510 139.120 42.960 ;
        RECT 139.300 41.010 139.560 43.140 ;
      LAYER li1 ;
        RECT 140.160 42.740 140.490 43.520 ;
        RECT 140.700 42.080 141.030 43.070 ;
        RECT 139.930 41.210 141.380 42.080 ;
        RECT 139.930 41.040 140.180 41.210 ;
        RECT 140.350 41.040 140.540 41.210 ;
        RECT 140.710 41.040 140.980 41.210 ;
        RECT 141.150 41.040 141.380 41.210 ;
        RECT 139.930 41.010 141.380 41.040 ;
        RECT 5.760 40.610 5.920 40.790 ;
        RECT 6.090 40.610 6.400 40.790 ;
        RECT 6.570 40.610 6.880 40.790 ;
        RECT 7.050 40.610 7.360 40.790 ;
        RECT 7.530 40.610 7.840 40.790 ;
        RECT 8.010 40.610 8.320 40.790 ;
        RECT 8.490 40.610 8.800 40.790 ;
        RECT 8.970 40.610 9.280 40.790 ;
        RECT 9.450 40.610 9.760 40.790 ;
        RECT 9.930 40.610 10.240 40.790 ;
        RECT 10.410 40.610 10.720 40.790 ;
        RECT 10.890 40.610 11.200 40.790 ;
        RECT 11.370 40.610 11.680 40.790 ;
        RECT 11.850 40.610 12.160 40.790 ;
        RECT 12.330 40.610 12.640 40.790 ;
        RECT 12.810 40.610 13.120 40.790 ;
        RECT 13.290 40.610 13.600 40.790 ;
        RECT 13.770 40.610 14.080 40.790 ;
        RECT 14.250 40.780 14.400 40.790 ;
        RECT 14.880 40.780 15.040 40.790 ;
        RECT 14.250 40.610 14.560 40.780 ;
        RECT 14.730 40.610 15.040 40.780 ;
        RECT 15.210 40.610 15.520 40.790 ;
        RECT 15.690 40.610 16.000 40.790 ;
        RECT 16.170 40.610 16.480 40.790 ;
        RECT 16.650 40.610 16.960 40.790 ;
        RECT 17.130 40.610 17.440 40.790 ;
        RECT 17.610 40.610 17.920 40.790 ;
        RECT 18.090 40.610 18.400 40.790 ;
        RECT 18.570 40.610 18.880 40.790 ;
        RECT 19.050 40.610 19.360 40.790 ;
        RECT 19.530 40.610 19.840 40.790 ;
        RECT 20.010 40.610 20.320 40.790 ;
        RECT 20.490 40.610 20.800 40.790 ;
        RECT 20.970 40.610 21.280 40.790 ;
        RECT 21.450 40.610 21.760 40.790 ;
        RECT 21.930 40.610 22.240 40.790 ;
        RECT 22.410 40.610 22.720 40.790 ;
        RECT 22.890 40.610 23.200 40.790 ;
        RECT 23.370 40.610 23.680 40.790 ;
        RECT 23.850 40.610 24.160 40.790 ;
        RECT 24.330 40.610 24.640 40.790 ;
        RECT 24.810 40.610 25.120 40.790 ;
        RECT 25.290 40.610 25.600 40.790 ;
        RECT 25.770 40.610 26.080 40.790 ;
        RECT 26.250 40.610 26.560 40.790 ;
        RECT 26.730 40.610 27.040 40.790 ;
        RECT 27.210 40.610 27.520 40.790 ;
        RECT 27.690 40.610 28.000 40.790 ;
        RECT 28.170 40.610 28.480 40.790 ;
        RECT 28.650 40.610 28.960 40.790 ;
        RECT 29.130 40.610 29.440 40.790 ;
        RECT 29.610 40.610 29.920 40.790 ;
        RECT 30.090 40.610 30.400 40.790 ;
        RECT 30.570 40.610 30.880 40.790 ;
        RECT 31.050 40.610 31.360 40.790 ;
        RECT 31.530 40.610 31.840 40.790 ;
        RECT 32.010 40.610 32.320 40.790 ;
        RECT 32.490 40.610 32.800 40.790 ;
        RECT 32.970 40.610 33.280 40.790 ;
        RECT 33.450 40.610 33.760 40.790 ;
        RECT 33.930 40.610 34.240 40.790 ;
        RECT 34.410 40.610 34.720 40.790 ;
        RECT 34.890 40.610 35.200 40.790 ;
        RECT 35.370 40.610 35.680 40.790 ;
        RECT 35.850 40.610 36.160 40.790 ;
        RECT 36.330 40.610 36.640 40.790 ;
        RECT 36.810 40.610 37.120 40.790 ;
        RECT 37.290 40.610 37.600 40.790 ;
        RECT 37.770 40.610 38.080 40.790 ;
        RECT 38.250 40.610 38.560 40.790 ;
        RECT 38.730 40.610 39.040 40.790 ;
        RECT 39.210 40.610 39.520 40.790 ;
        RECT 39.690 40.610 40.000 40.790 ;
        RECT 40.170 40.610 40.480 40.790 ;
        RECT 40.650 40.610 40.960 40.790 ;
        RECT 41.130 40.610 41.440 40.790 ;
        RECT 41.610 40.610 41.920 40.790 ;
        RECT 42.090 40.610 42.400 40.790 ;
        RECT 42.570 40.610 42.880 40.790 ;
        RECT 43.050 40.610 43.360 40.790 ;
        RECT 43.530 40.610 43.840 40.790 ;
        RECT 44.010 40.610 44.320 40.790 ;
        RECT 44.490 40.610 44.800 40.790 ;
        RECT 44.970 40.610 45.280 40.790 ;
        RECT 45.450 40.610 45.760 40.790 ;
        RECT 45.930 40.610 46.240 40.790 ;
        RECT 46.410 40.610 46.720 40.790 ;
        RECT 46.890 40.610 47.200 40.790 ;
        RECT 47.370 40.610 47.680 40.790 ;
        RECT 47.850 40.610 48.160 40.790 ;
        RECT 48.330 40.610 48.640 40.790 ;
        RECT 48.810 40.610 49.120 40.790 ;
        RECT 49.290 40.610 49.600 40.790 ;
        RECT 49.770 40.610 50.080 40.790 ;
        RECT 50.250 40.610 50.560 40.790 ;
        RECT 50.730 40.610 51.040 40.790 ;
        RECT 51.210 40.610 51.520 40.790 ;
        RECT 51.690 40.610 52.000 40.790 ;
        RECT 52.170 40.610 52.480 40.790 ;
        RECT 52.650 40.610 52.960 40.790 ;
        RECT 53.130 40.610 53.440 40.790 ;
        RECT 53.610 40.610 53.920 40.790 ;
        RECT 54.090 40.610 54.400 40.790 ;
        RECT 54.570 40.610 54.880 40.790 ;
        RECT 55.050 40.610 55.360 40.790 ;
        RECT 55.530 40.610 55.840 40.790 ;
        RECT 56.010 40.610 56.320 40.790 ;
        RECT 56.490 40.610 56.800 40.790 ;
        RECT 56.970 40.610 57.280 40.790 ;
        RECT 57.450 40.610 57.760 40.790 ;
        RECT 57.930 40.610 58.240 40.790 ;
        RECT 58.410 40.610 58.720 40.790 ;
        RECT 58.890 40.610 59.200 40.790 ;
        RECT 59.370 40.610 59.680 40.790 ;
        RECT 59.850 40.610 60.160 40.790 ;
        RECT 60.330 40.610 60.640 40.790 ;
        RECT 60.810 40.610 61.120 40.790 ;
        RECT 61.290 40.610 61.600 40.790 ;
        RECT 61.770 40.610 62.080 40.790 ;
        RECT 62.250 40.610 62.560 40.790 ;
        RECT 62.730 40.610 63.040 40.790 ;
        RECT 63.210 40.610 63.520 40.790 ;
        RECT 63.690 40.610 64.000 40.790 ;
        RECT 64.170 40.610 64.480 40.790 ;
        RECT 64.650 40.610 64.960 40.790 ;
        RECT 65.130 40.610 65.440 40.790 ;
        RECT 65.610 40.610 65.920 40.790 ;
        RECT 66.090 40.610 66.400 40.790 ;
        RECT 66.570 40.610 66.880 40.790 ;
        RECT 67.050 40.610 67.360 40.790 ;
        RECT 67.530 40.610 67.840 40.790 ;
        RECT 68.010 40.610 68.320 40.790 ;
        RECT 68.490 40.610 68.800 40.790 ;
        RECT 68.970 40.610 69.280 40.790 ;
        RECT 69.450 40.610 69.760 40.790 ;
        RECT 69.930 40.610 70.240 40.790 ;
        RECT 70.410 40.610 70.720 40.790 ;
        RECT 70.890 40.610 71.200 40.790 ;
        RECT 71.370 40.610 71.680 40.790 ;
        RECT 71.850 40.610 72.160 40.790 ;
        RECT 72.330 40.610 72.640 40.790 ;
        RECT 72.810 40.610 73.120 40.790 ;
        RECT 73.290 40.610 73.600 40.790 ;
        RECT 73.770 40.610 74.080 40.790 ;
        RECT 74.250 40.610 74.560 40.790 ;
        RECT 74.730 40.610 75.040 40.790 ;
        RECT 75.210 40.610 75.520 40.790 ;
        RECT 75.690 40.610 76.000 40.790 ;
        RECT 76.170 40.610 76.480 40.790 ;
        RECT 76.650 40.610 76.960 40.790 ;
        RECT 77.130 40.610 77.440 40.790 ;
        RECT 77.610 40.780 77.760 40.790 ;
        RECT 78.240 40.780 78.400 40.790 ;
        RECT 77.610 40.610 77.920 40.780 ;
        RECT 78.090 40.610 78.400 40.780 ;
        RECT 78.570 40.610 78.880 40.790 ;
        RECT 79.050 40.610 79.360 40.790 ;
        RECT 79.530 40.610 79.840 40.790 ;
        RECT 80.010 40.610 80.320 40.790 ;
        RECT 80.490 40.610 80.800 40.790 ;
        RECT 80.970 40.610 81.280 40.790 ;
        RECT 81.450 40.610 81.760 40.790 ;
        RECT 81.930 40.610 82.240 40.790 ;
        RECT 82.410 40.610 82.720 40.790 ;
        RECT 82.890 40.610 83.200 40.790 ;
        RECT 83.370 40.610 83.680 40.790 ;
        RECT 83.850 40.610 84.160 40.790 ;
        RECT 84.330 40.610 84.640 40.790 ;
        RECT 84.810 40.610 85.120 40.790 ;
        RECT 85.290 40.610 85.600 40.790 ;
        RECT 85.770 40.610 86.080 40.790 ;
        RECT 86.250 40.610 86.560 40.790 ;
        RECT 86.730 40.610 87.040 40.790 ;
        RECT 87.210 40.610 87.520 40.790 ;
        RECT 87.690 40.610 88.000 40.790 ;
        RECT 88.170 40.610 88.480 40.790 ;
        RECT 88.650 40.610 88.960 40.790 ;
        RECT 89.130 40.610 89.440 40.790 ;
        RECT 89.610 40.610 89.920 40.790 ;
        RECT 90.090 40.610 90.400 40.790 ;
        RECT 90.570 40.610 90.880 40.790 ;
        RECT 91.050 40.610 91.360 40.790 ;
        RECT 91.530 40.610 91.840 40.790 ;
        RECT 92.010 40.610 92.320 40.790 ;
        RECT 92.490 40.610 92.800 40.790 ;
        RECT 92.970 40.610 93.280 40.790 ;
        RECT 93.450 40.610 93.760 40.790 ;
        RECT 93.930 40.610 94.240 40.790 ;
        RECT 94.410 40.610 94.720 40.790 ;
        RECT 94.890 40.610 95.200 40.790 ;
        RECT 95.370 40.610 95.680 40.790 ;
        RECT 95.850 40.610 96.160 40.790 ;
        RECT 96.330 40.610 96.640 40.790 ;
        RECT 96.810 40.610 97.120 40.790 ;
        RECT 97.290 40.610 97.600 40.790 ;
        RECT 97.770 40.610 98.080 40.790 ;
        RECT 98.250 40.610 98.560 40.790 ;
        RECT 98.730 40.610 99.040 40.790 ;
        RECT 99.210 40.610 99.520 40.790 ;
        RECT 99.690 40.610 100.000 40.790 ;
        RECT 100.170 40.610 100.480 40.790 ;
        RECT 100.650 40.610 100.960 40.790 ;
        RECT 101.130 40.610 101.440 40.790 ;
        RECT 101.610 40.610 101.920 40.790 ;
        RECT 102.090 40.610 102.400 40.790 ;
        RECT 102.570 40.610 102.880 40.790 ;
        RECT 103.050 40.610 103.360 40.790 ;
        RECT 103.530 40.610 103.840 40.790 ;
        RECT 104.010 40.610 104.320 40.790 ;
        RECT 104.490 40.610 104.800 40.790 ;
        RECT 104.970 40.610 105.280 40.790 ;
        RECT 105.450 40.610 105.760 40.790 ;
        RECT 105.930 40.610 106.240 40.790 ;
        RECT 106.410 40.610 106.720 40.790 ;
        RECT 106.890 40.610 107.200 40.790 ;
        RECT 107.370 40.610 107.680 40.790 ;
        RECT 107.850 40.610 108.160 40.790 ;
        RECT 108.330 40.610 108.640 40.790 ;
        RECT 108.810 40.610 109.120 40.790 ;
        RECT 109.290 40.610 109.600 40.790 ;
        RECT 109.770 40.610 110.080 40.790 ;
        RECT 110.250 40.780 110.400 40.790 ;
        RECT 110.880 40.780 111.040 40.790 ;
        RECT 110.250 40.610 110.560 40.780 ;
        RECT 110.730 40.610 111.040 40.780 ;
        RECT 111.210 40.610 111.520 40.790 ;
        RECT 111.690 40.610 112.000 40.790 ;
        RECT 112.170 40.610 112.480 40.790 ;
        RECT 112.650 40.610 112.960 40.790 ;
        RECT 113.130 40.610 113.440 40.790 ;
        RECT 113.610 40.610 113.920 40.790 ;
        RECT 114.090 40.610 114.400 40.790 ;
        RECT 114.570 40.610 114.880 40.790 ;
        RECT 115.050 40.610 115.360 40.790 ;
        RECT 115.530 40.780 115.840 40.790 ;
        RECT 116.010 40.780 116.320 40.790 ;
        RECT 115.530 40.610 115.680 40.780 ;
        RECT 116.160 40.610 116.320 40.780 ;
        RECT 116.490 40.610 116.800 40.790 ;
        RECT 116.970 40.610 117.280 40.790 ;
        RECT 117.450 40.610 117.760 40.790 ;
        RECT 117.930 40.610 118.240 40.790 ;
        RECT 118.410 40.610 118.720 40.790 ;
        RECT 118.890 40.610 119.200 40.790 ;
        RECT 119.370 40.610 119.680 40.790 ;
        RECT 119.850 40.610 120.160 40.790 ;
        RECT 120.330 40.610 120.640 40.790 ;
        RECT 120.810 40.610 121.120 40.790 ;
        RECT 121.290 40.610 121.600 40.790 ;
        RECT 121.770 40.610 122.080 40.790 ;
        RECT 122.250 40.610 122.560 40.790 ;
        RECT 122.730 40.610 123.040 40.790 ;
        RECT 123.210 40.610 123.520 40.790 ;
        RECT 123.690 40.610 124.000 40.790 ;
        RECT 124.170 40.610 124.480 40.790 ;
        RECT 124.650 40.610 124.960 40.790 ;
        RECT 125.130 40.610 125.440 40.790 ;
        RECT 125.610 40.610 125.920 40.790 ;
        RECT 126.090 40.610 126.400 40.790 ;
        RECT 126.570 40.610 126.880 40.790 ;
        RECT 127.050 40.610 127.360 40.790 ;
        RECT 127.530 40.610 127.840 40.790 ;
        RECT 128.010 40.610 128.320 40.790 ;
        RECT 128.490 40.610 128.800 40.790 ;
        RECT 128.970 40.610 129.280 40.790 ;
        RECT 129.450 40.610 129.760 40.790 ;
        RECT 129.930 40.610 130.240 40.790 ;
        RECT 130.410 40.610 130.720 40.790 ;
        RECT 130.890 40.610 131.200 40.790 ;
        RECT 131.370 40.610 131.680 40.790 ;
        RECT 131.850 40.610 132.160 40.790 ;
        RECT 132.330 40.610 132.640 40.790 ;
        RECT 132.810 40.610 133.120 40.790 ;
        RECT 133.290 40.610 133.600 40.790 ;
        RECT 133.770 40.610 134.080 40.790 ;
        RECT 134.250 40.610 134.560 40.790 ;
        RECT 134.730 40.610 135.040 40.790 ;
        RECT 135.210 40.610 135.520 40.790 ;
        RECT 135.690 40.610 136.000 40.790 ;
        RECT 136.170 40.610 136.480 40.790 ;
        RECT 136.650 40.610 136.960 40.790 ;
        RECT 137.130 40.610 137.440 40.790 ;
        RECT 137.610 40.610 137.920 40.790 ;
        RECT 138.090 40.610 138.400 40.790 ;
        RECT 138.570 40.610 138.880 40.790 ;
        RECT 139.050 40.610 139.360 40.790 ;
        RECT 139.530 40.610 139.840 40.790 ;
        RECT 140.010 40.610 140.320 40.790 ;
        RECT 140.490 40.610 140.800 40.790 ;
        RECT 140.970 40.610 141.280 40.790 ;
        RECT 141.450 40.780 141.760 40.790 ;
        RECT 141.930 40.780 142.080 40.790 ;
        RECT 141.450 40.610 141.600 40.780 ;
        RECT 6.260 40.360 9.000 40.380 ;
        RECT 6.260 40.190 6.470 40.360 ;
        RECT 6.640 40.190 6.910 40.360 ;
        RECT 7.080 40.190 7.320 40.360 ;
        RECT 7.490 40.190 7.750 40.360 ;
        RECT 7.920 40.190 8.190 40.360 ;
        RECT 8.360 40.190 8.600 40.360 ;
        RECT 8.770 40.190 9.000 40.360 ;
        RECT 6.260 39.310 9.000 40.190 ;
        RECT 10.100 40.360 12.840 40.380 ;
        RECT 10.100 40.190 10.310 40.360 ;
        RECT 10.480 40.190 10.750 40.360 ;
        RECT 10.920 40.190 11.160 40.360 ;
        RECT 11.330 40.190 11.590 40.360 ;
        RECT 11.760 40.190 12.030 40.360 ;
        RECT 12.200 40.190 12.440 40.360 ;
        RECT 12.610 40.190 12.840 40.360 ;
        RECT 10.100 39.310 12.840 40.190 ;
        RECT 14.970 40.310 15.560 40.390 ;
        RECT 14.970 40.140 15.000 40.310 ;
        RECT 15.170 40.140 15.360 40.310 ;
        RECT 15.530 40.140 15.560 40.310 ;
        RECT 6.500 37.990 6.830 38.660 ;
        RECT 7.230 38.330 7.560 39.310 ;
        RECT 7.780 37.990 8.110 38.660 ;
        RECT 8.510 38.330 8.840 39.310 ;
        RECT 10.340 37.990 10.670 38.660 ;
        RECT 11.070 38.330 11.400 39.310 ;
        RECT 11.620 37.990 11.950 38.660 ;
        RECT 12.350 38.330 12.680 39.310 ;
        RECT 14.970 38.810 15.560 40.140 ;
      LAYER li1 ;
        RECT 15.840 38.810 16.230 40.390 ;
      LAYER li1 ;
        RECT 16.570 40.360 18.020 40.390 ;
        RECT 16.570 40.190 16.820 40.360 ;
        RECT 16.990 40.190 17.180 40.360 ;
        RECT 17.350 40.190 17.620 40.360 ;
        RECT 17.790 40.190 18.020 40.360 ;
        RECT 16.570 39.320 18.020 40.190 ;
        RECT 18.330 40.310 20.000 40.390 ;
        RECT 18.330 40.140 18.360 40.310 ;
        RECT 18.530 40.140 18.720 40.310 ;
        RECT 18.890 40.140 19.080 40.310 ;
        RECT 19.250 40.140 19.440 40.310 ;
        RECT 19.610 40.140 19.800 40.310 ;
        RECT 19.970 40.140 20.000 40.310 ;
      LAYER li1 ;
        RECT 15.010 38.180 15.720 38.570 ;
      LAYER li1 ;
        RECT 6.340 36.990 9.070 37.990 ;
        RECT 10.180 36.990 12.910 37.990 ;
        RECT 14.970 37.000 15.560 37.960 ;
      LAYER li1 ;
        RECT 15.900 37.130 16.230 38.810 ;
      LAYER li1 ;
        RECT 16.800 37.880 17.130 38.660 ;
        RECT 17.340 38.330 17.670 39.320 ;
        RECT 18.330 38.930 20.000 40.140 ;
      LAYER li1 ;
        RECT 18.370 38.410 19.560 38.750 ;
        RECT 19.740 38.410 20.070 38.750 ;
        RECT 20.260 38.230 20.520 40.390 ;
      LAYER li1 ;
        RECT 20.890 40.360 22.340 40.390 ;
        RECT 20.890 40.190 21.140 40.360 ;
        RECT 21.310 40.190 21.500 40.360 ;
        RECT 21.670 40.190 21.940 40.360 ;
        RECT 22.110 40.190 22.340 40.360 ;
        RECT 20.890 39.320 22.340 40.190 ;
        RECT 22.650 40.310 24.320 40.390 ;
        RECT 22.650 40.140 22.680 40.310 ;
        RECT 22.850 40.140 23.040 40.310 ;
        RECT 23.210 40.140 23.400 40.310 ;
        RECT 23.570 40.140 23.760 40.310 ;
        RECT 23.930 40.140 24.120 40.310 ;
        RECT 24.290 40.140 24.320 40.310 ;
      LAYER li1 ;
        RECT 19.440 38.060 20.520 38.230 ;
      LAYER li1 ;
        RECT 16.800 37.480 18.100 37.880 ;
        RECT 16.490 37.000 18.100 37.480 ;
        RECT 18.330 37.000 19.260 37.960 ;
      LAYER li1 ;
        RECT 19.440 37.130 19.770 38.060 ;
      LAYER li1 ;
        RECT 21.120 37.880 21.450 38.660 ;
        RECT 21.660 38.330 21.990 39.320 ;
        RECT 22.650 38.930 24.320 40.140 ;
      LAYER li1 ;
        RECT 22.690 38.410 23.880 38.750 ;
        RECT 24.060 38.410 24.390 38.750 ;
        RECT 24.580 38.230 24.840 40.390 ;
      LAYER li1 ;
        RECT 25.210 40.360 26.660 40.390 ;
        RECT 25.210 40.190 25.460 40.360 ;
        RECT 25.630 40.190 25.820 40.360 ;
        RECT 25.990 40.190 26.260 40.360 ;
        RECT 26.430 40.190 26.660 40.360 ;
        RECT 25.210 39.320 26.660 40.190 ;
        RECT 26.970 40.310 28.640 40.390 ;
        RECT 26.970 40.140 27.000 40.310 ;
        RECT 27.170 40.140 27.360 40.310 ;
        RECT 27.530 40.140 27.720 40.310 ;
        RECT 27.890 40.140 28.080 40.310 ;
        RECT 28.250 40.140 28.440 40.310 ;
        RECT 28.610 40.140 28.640 40.310 ;
      LAYER li1 ;
        RECT 23.760 38.060 24.840 38.230 ;
      LAYER li1 ;
        RECT 19.960 37.000 20.550 37.880 ;
        RECT 21.120 37.480 22.420 37.880 ;
        RECT 20.810 37.000 22.420 37.480 ;
        RECT 22.650 37.000 23.580 37.960 ;
      LAYER li1 ;
        RECT 23.760 37.130 24.090 38.060 ;
      LAYER li1 ;
        RECT 25.440 37.880 25.770 38.660 ;
        RECT 25.980 38.330 26.310 39.320 ;
        RECT 26.970 38.930 28.640 40.140 ;
      LAYER li1 ;
        RECT 27.010 38.160 27.310 38.750 ;
        RECT 27.490 38.410 28.680 38.750 ;
        RECT 28.860 38.410 29.190 39.890 ;
        RECT 29.370 38.230 29.640 40.390 ;
      LAYER li1 ;
        RECT 30.490 40.360 31.940 40.390 ;
        RECT 30.490 40.190 30.740 40.360 ;
        RECT 30.910 40.190 31.100 40.360 ;
        RECT 31.270 40.190 31.540 40.360 ;
        RECT 31.710 40.190 31.940 40.360 ;
        RECT 30.490 39.320 31.940 40.190 ;
        RECT 32.250 40.310 33.920 40.390 ;
        RECT 32.250 40.140 32.280 40.310 ;
        RECT 32.450 40.140 32.640 40.310 ;
        RECT 32.810 40.140 33.000 40.310 ;
        RECT 33.170 40.140 33.360 40.310 ;
        RECT 33.530 40.140 33.720 40.310 ;
        RECT 33.890 40.140 33.920 40.310 ;
      LAYER li1 ;
        RECT 27.810 38.060 29.640 38.230 ;
      LAYER li1 ;
        RECT 24.280 37.000 24.870 37.880 ;
        RECT 25.440 37.480 26.740 37.880 ;
        RECT 25.130 37.000 26.740 37.480 ;
        RECT 26.970 37.000 27.560 37.960 ;
      LAYER li1 ;
        RECT 27.810 37.130 28.060 38.060 ;
      LAYER li1 ;
        RECT 28.240 37.000 29.190 37.880 ;
      LAYER li1 ;
        RECT 29.370 37.130 29.640 38.060 ;
      LAYER li1 ;
        RECT 30.720 37.880 31.050 38.660 ;
        RECT 31.260 38.330 31.590 39.320 ;
        RECT 32.250 38.930 33.920 40.140 ;
      LAYER li1 ;
        RECT 32.290 38.160 32.590 38.750 ;
        RECT 32.770 38.410 33.960 38.750 ;
        RECT 34.140 38.410 34.470 39.890 ;
        RECT 34.650 38.230 34.920 40.390 ;
      LAYER li1 ;
        RECT 35.770 40.360 37.220 40.390 ;
        RECT 35.770 40.190 36.020 40.360 ;
        RECT 36.190 40.190 36.380 40.360 ;
        RECT 36.550 40.190 36.820 40.360 ;
        RECT 36.990 40.190 37.220 40.360 ;
        RECT 35.770 39.320 37.220 40.190 ;
        RECT 37.530 40.310 38.480 40.390 ;
        RECT 37.530 40.140 37.560 40.310 ;
        RECT 37.730 40.140 37.920 40.310 ;
        RECT 38.090 40.140 38.280 40.310 ;
        RECT 38.450 40.140 38.480 40.310 ;
      LAYER li1 ;
        RECT 33.090 38.060 34.920 38.230 ;
      LAYER li1 ;
        RECT 30.720 37.480 32.020 37.880 ;
        RECT 30.410 37.000 32.020 37.480 ;
        RECT 32.250 37.000 32.840 37.960 ;
      LAYER li1 ;
        RECT 33.090 37.130 33.340 38.060 ;
      LAYER li1 ;
        RECT 33.520 37.000 34.470 37.880 ;
      LAYER li1 ;
        RECT 34.650 37.130 34.920 38.060 ;
      LAYER li1 ;
        RECT 36.000 37.880 36.330 38.660 ;
        RECT 36.540 38.330 36.870 39.320 ;
        RECT 37.530 38.810 38.480 40.140 ;
      LAYER li1 ;
        RECT 38.660 38.710 38.910 40.390 ;
      LAYER li1 ;
        RECT 39.090 40.310 40.040 40.390 ;
        RECT 39.090 40.140 39.120 40.310 ;
        RECT 39.290 40.140 39.480 40.310 ;
        RECT 39.650 40.140 39.840 40.310 ;
        RECT 40.010 40.140 40.040 40.310 ;
        RECT 39.090 38.890 40.040 40.140 ;
      LAYER li1 ;
        RECT 40.220 38.710 40.550 40.390 ;
      LAYER li1 ;
        RECT 40.730 40.310 41.680 40.390 ;
        RECT 40.730 40.140 40.760 40.310 ;
        RECT 40.930 40.140 41.120 40.310 ;
        RECT 41.290 40.140 41.480 40.310 ;
        RECT 41.650 40.140 41.680 40.310 ;
        RECT 40.730 38.930 41.680 40.140 ;
      LAYER li1 ;
        RECT 38.660 38.540 40.550 38.710 ;
        RECT 38.660 38.410 38.830 38.540 ;
        RECT 41.330 38.410 41.660 38.750 ;
        RECT 37.570 38.180 38.830 38.410 ;
      LAYER li1 ;
        RECT 39.010 38.230 41.040 38.360 ;
        RECT 41.860 38.230 42.110 40.390 ;
        RECT 42.490 40.360 43.940 40.390 ;
        RECT 42.490 40.190 42.740 40.360 ;
        RECT 42.910 40.190 43.100 40.360 ;
        RECT 43.270 40.190 43.540 40.360 ;
        RECT 43.710 40.190 43.940 40.360 ;
        RECT 42.490 39.320 43.940 40.190 ;
        RECT 44.250 40.310 45.200 40.390 ;
        RECT 44.250 40.140 44.280 40.310 ;
        RECT 44.450 40.140 44.640 40.310 ;
        RECT 44.810 40.140 45.000 40.310 ;
        RECT 45.170 40.140 45.200 40.310 ;
        RECT 39.010 38.190 42.110 38.230 ;
      LAYER li1 ;
        RECT 38.660 38.010 38.830 38.180 ;
      LAYER li1 ;
        RECT 40.870 38.060 42.110 38.190 ;
        RECT 36.000 37.480 37.300 37.880 ;
        RECT 35.690 37.000 37.300 37.480 ;
        RECT 37.530 37.000 38.480 37.960 ;
      LAYER li1 ;
        RECT 38.660 37.840 40.470 38.010 ;
        RECT 38.660 37.130 38.910 37.840 ;
      LAYER li1 ;
        RECT 39.090 37.000 40.040 37.660 ;
      LAYER li1 ;
        RECT 40.220 37.130 40.470 37.840 ;
      LAYER li1 ;
        RECT 40.650 37.000 41.600 37.880 ;
        RECT 41.780 37.130 42.110 38.060 ;
        RECT 42.720 37.880 43.050 38.660 ;
        RECT 43.260 38.330 43.590 39.320 ;
        RECT 44.250 38.810 45.200 40.140 ;
      LAYER li1 ;
        RECT 45.380 38.710 45.630 40.390 ;
      LAYER li1 ;
        RECT 45.810 40.310 46.760 40.390 ;
        RECT 45.810 40.140 45.840 40.310 ;
        RECT 46.010 40.140 46.200 40.310 ;
        RECT 46.370 40.140 46.560 40.310 ;
        RECT 46.730 40.140 46.760 40.310 ;
        RECT 45.810 38.890 46.760 40.140 ;
      LAYER li1 ;
        RECT 46.940 38.710 47.270 40.390 ;
      LAYER li1 ;
        RECT 47.450 40.310 48.400 40.390 ;
        RECT 47.450 40.140 47.480 40.310 ;
        RECT 47.650 40.140 47.840 40.310 ;
        RECT 48.010 40.140 48.200 40.310 ;
        RECT 48.370 40.140 48.400 40.310 ;
        RECT 47.450 38.930 48.400 40.140 ;
      LAYER li1 ;
        RECT 45.380 38.540 47.270 38.710 ;
        RECT 45.380 38.410 45.550 38.540 ;
        RECT 48.050 38.410 48.380 38.750 ;
        RECT 44.290 38.180 45.550 38.410 ;
      LAYER li1 ;
        RECT 45.730 38.230 47.760 38.360 ;
        RECT 48.580 38.230 48.830 40.390 ;
        RECT 49.210 40.360 50.660 40.390 ;
        RECT 49.210 40.190 49.460 40.360 ;
        RECT 49.630 40.190 49.820 40.360 ;
        RECT 49.990 40.190 50.260 40.360 ;
        RECT 50.430 40.190 50.660 40.360 ;
        RECT 49.210 39.320 50.660 40.190 ;
        RECT 50.970 40.310 51.920 40.390 ;
        RECT 50.970 40.140 51.000 40.310 ;
        RECT 51.170 40.140 51.360 40.310 ;
        RECT 51.530 40.140 51.720 40.310 ;
        RECT 51.890 40.140 51.920 40.310 ;
        RECT 45.730 38.190 48.830 38.230 ;
      LAYER li1 ;
        RECT 45.380 38.010 45.550 38.180 ;
      LAYER li1 ;
        RECT 47.590 38.060 48.830 38.190 ;
        RECT 42.720 37.480 44.020 37.880 ;
        RECT 42.410 37.000 44.020 37.480 ;
        RECT 44.250 37.000 45.200 37.960 ;
      LAYER li1 ;
        RECT 45.380 37.840 47.190 38.010 ;
        RECT 45.380 37.130 45.630 37.840 ;
      LAYER li1 ;
        RECT 45.810 37.000 46.760 37.660 ;
      LAYER li1 ;
        RECT 46.940 37.130 47.190 37.840 ;
      LAYER li1 ;
        RECT 47.370 37.000 48.320 37.880 ;
        RECT 48.500 37.130 48.830 38.060 ;
        RECT 49.440 37.880 49.770 38.660 ;
        RECT 49.980 38.330 50.310 39.320 ;
        RECT 50.970 38.810 51.920 40.140 ;
      LAYER li1 ;
        RECT 52.100 38.710 52.350 40.390 ;
      LAYER li1 ;
        RECT 52.530 40.310 53.480 40.390 ;
        RECT 52.530 40.140 52.560 40.310 ;
        RECT 52.730 40.140 52.920 40.310 ;
        RECT 53.090 40.140 53.280 40.310 ;
        RECT 53.450 40.140 53.480 40.310 ;
        RECT 52.530 38.890 53.480 40.140 ;
      LAYER li1 ;
        RECT 53.660 38.710 53.990 40.390 ;
      LAYER li1 ;
        RECT 54.170 40.310 55.120 40.390 ;
        RECT 54.170 40.140 54.200 40.310 ;
        RECT 54.370 40.140 54.560 40.310 ;
        RECT 54.730 40.140 54.920 40.310 ;
        RECT 55.090 40.140 55.120 40.310 ;
        RECT 54.170 38.930 55.120 40.140 ;
      LAYER li1 ;
        RECT 52.100 38.540 53.990 38.710 ;
        RECT 52.100 38.410 52.270 38.540 ;
        RECT 54.770 38.410 55.100 38.750 ;
        RECT 51.010 38.180 52.270 38.410 ;
      LAYER li1 ;
        RECT 52.450 38.230 54.480 38.360 ;
        RECT 55.300 38.230 55.550 40.390 ;
        RECT 55.930 40.360 57.380 40.390 ;
        RECT 55.930 40.190 56.180 40.360 ;
        RECT 56.350 40.190 56.540 40.360 ;
        RECT 56.710 40.190 56.980 40.360 ;
        RECT 57.150 40.190 57.380 40.360 ;
        RECT 55.930 39.320 57.380 40.190 ;
        RECT 57.690 40.310 58.640 40.390 ;
        RECT 57.690 40.140 57.720 40.310 ;
        RECT 57.890 40.140 58.080 40.310 ;
        RECT 58.250 40.140 58.440 40.310 ;
        RECT 58.610 40.140 58.640 40.310 ;
        RECT 52.450 38.190 55.550 38.230 ;
      LAYER li1 ;
        RECT 52.100 38.010 52.270 38.180 ;
      LAYER li1 ;
        RECT 54.310 38.060 55.550 38.190 ;
        RECT 49.440 37.480 50.740 37.880 ;
        RECT 49.130 37.000 50.740 37.480 ;
        RECT 50.970 37.000 51.920 37.960 ;
      LAYER li1 ;
        RECT 52.100 37.840 53.910 38.010 ;
        RECT 52.100 37.130 52.350 37.840 ;
      LAYER li1 ;
        RECT 52.530 37.000 53.480 37.660 ;
      LAYER li1 ;
        RECT 53.660 37.130 53.910 37.840 ;
      LAYER li1 ;
        RECT 54.090 37.000 55.040 37.880 ;
        RECT 55.220 37.130 55.550 38.060 ;
        RECT 56.160 37.880 56.490 38.660 ;
        RECT 56.700 38.330 57.030 39.320 ;
        RECT 57.690 38.810 58.640 40.140 ;
      LAYER li1 ;
        RECT 58.820 38.710 59.070 40.390 ;
      LAYER li1 ;
        RECT 59.250 40.310 60.200 40.390 ;
        RECT 59.250 40.140 59.280 40.310 ;
        RECT 59.450 40.140 59.640 40.310 ;
        RECT 59.810 40.140 60.000 40.310 ;
        RECT 60.170 40.140 60.200 40.310 ;
        RECT 59.250 38.890 60.200 40.140 ;
      LAYER li1 ;
        RECT 60.380 38.710 60.710 40.390 ;
      LAYER li1 ;
        RECT 60.890 40.310 61.840 40.390 ;
        RECT 60.890 40.140 60.920 40.310 ;
        RECT 61.090 40.140 61.280 40.310 ;
        RECT 61.450 40.140 61.640 40.310 ;
        RECT 61.810 40.140 61.840 40.310 ;
        RECT 60.890 38.930 61.840 40.140 ;
      LAYER li1 ;
        RECT 58.820 38.540 60.710 38.710 ;
        RECT 58.820 38.410 58.990 38.540 ;
        RECT 61.490 38.410 61.820 38.750 ;
        RECT 57.730 38.180 58.990 38.410 ;
      LAYER li1 ;
        RECT 59.170 38.230 61.200 38.360 ;
        RECT 62.020 38.230 62.270 40.390 ;
        RECT 62.650 40.360 64.100 40.390 ;
        RECT 62.650 40.190 62.900 40.360 ;
        RECT 63.070 40.190 63.260 40.360 ;
        RECT 63.430 40.190 63.700 40.360 ;
        RECT 63.870 40.190 64.100 40.360 ;
        RECT 62.650 39.320 64.100 40.190 ;
        RECT 64.410 40.310 65.360 40.390 ;
        RECT 64.410 40.140 64.440 40.310 ;
        RECT 64.610 40.140 64.800 40.310 ;
        RECT 64.970 40.140 65.160 40.310 ;
        RECT 65.330 40.140 65.360 40.310 ;
        RECT 59.170 38.190 62.270 38.230 ;
      LAYER li1 ;
        RECT 58.820 38.010 58.990 38.180 ;
      LAYER li1 ;
        RECT 61.030 38.060 62.270 38.190 ;
        RECT 56.160 37.480 57.460 37.880 ;
        RECT 55.850 37.000 57.460 37.480 ;
        RECT 57.690 37.000 58.640 37.960 ;
      LAYER li1 ;
        RECT 58.820 37.840 60.630 38.010 ;
        RECT 58.820 37.130 59.070 37.840 ;
      LAYER li1 ;
        RECT 59.250 37.000 60.200 37.660 ;
      LAYER li1 ;
        RECT 60.380 37.130 60.630 37.840 ;
      LAYER li1 ;
        RECT 60.810 37.000 61.760 37.880 ;
        RECT 61.940 37.130 62.270 38.060 ;
        RECT 62.880 37.880 63.210 38.660 ;
        RECT 63.420 38.330 63.750 39.320 ;
        RECT 64.410 38.810 65.360 40.140 ;
      LAYER li1 ;
        RECT 65.540 38.710 65.790 40.390 ;
      LAYER li1 ;
        RECT 65.970 40.310 66.920 40.390 ;
        RECT 65.970 40.140 66.000 40.310 ;
        RECT 66.170 40.140 66.360 40.310 ;
        RECT 66.530 40.140 66.720 40.310 ;
        RECT 66.890 40.140 66.920 40.310 ;
        RECT 65.970 38.890 66.920 40.140 ;
      LAYER li1 ;
        RECT 67.100 38.710 67.430 40.390 ;
      LAYER li1 ;
        RECT 67.610 40.310 68.560 40.390 ;
        RECT 67.610 40.140 67.640 40.310 ;
        RECT 67.810 40.140 68.000 40.310 ;
        RECT 68.170 40.140 68.360 40.310 ;
        RECT 68.530 40.140 68.560 40.310 ;
        RECT 67.610 38.930 68.560 40.140 ;
      LAYER li1 ;
        RECT 65.540 38.540 67.430 38.710 ;
        RECT 65.540 38.410 65.710 38.540 ;
        RECT 68.210 38.410 68.540 38.750 ;
        RECT 64.450 38.180 65.710 38.410 ;
      LAYER li1 ;
        RECT 65.890 38.230 67.920 38.360 ;
        RECT 68.740 38.230 68.990 40.390 ;
        RECT 69.370 40.360 70.820 40.390 ;
        RECT 69.370 40.190 69.620 40.360 ;
        RECT 69.790 40.190 69.980 40.360 ;
        RECT 70.150 40.190 70.420 40.360 ;
        RECT 70.590 40.190 70.820 40.360 ;
        RECT 69.370 39.320 70.820 40.190 ;
        RECT 71.130 40.310 72.080 40.390 ;
        RECT 71.130 40.140 71.160 40.310 ;
        RECT 71.330 40.140 71.520 40.310 ;
        RECT 71.690 40.140 71.880 40.310 ;
        RECT 72.050 40.140 72.080 40.310 ;
        RECT 65.890 38.190 68.990 38.230 ;
      LAYER li1 ;
        RECT 65.540 38.010 65.710 38.180 ;
      LAYER li1 ;
        RECT 67.750 38.060 68.990 38.190 ;
        RECT 62.880 37.480 64.180 37.880 ;
        RECT 62.570 37.000 64.180 37.480 ;
        RECT 64.410 37.000 65.360 37.960 ;
      LAYER li1 ;
        RECT 65.540 37.840 67.350 38.010 ;
        RECT 65.540 37.130 65.790 37.840 ;
      LAYER li1 ;
        RECT 65.970 37.000 66.920 37.660 ;
      LAYER li1 ;
        RECT 67.100 37.130 67.350 37.840 ;
      LAYER li1 ;
        RECT 67.530 37.000 68.480 37.880 ;
        RECT 68.660 37.130 68.990 38.060 ;
        RECT 69.600 37.880 69.930 38.660 ;
        RECT 70.140 38.330 70.470 39.320 ;
        RECT 71.130 38.810 72.080 40.140 ;
      LAYER li1 ;
        RECT 72.260 38.710 72.510 40.390 ;
      LAYER li1 ;
        RECT 72.690 40.310 73.640 40.390 ;
        RECT 72.690 40.140 72.720 40.310 ;
        RECT 72.890 40.140 73.080 40.310 ;
        RECT 73.250 40.140 73.440 40.310 ;
        RECT 73.610 40.140 73.640 40.310 ;
        RECT 72.690 38.890 73.640 40.140 ;
      LAYER li1 ;
        RECT 73.820 38.710 74.150 40.390 ;
      LAYER li1 ;
        RECT 74.330 40.310 75.280 40.390 ;
        RECT 74.330 40.140 74.360 40.310 ;
        RECT 74.530 40.140 74.720 40.310 ;
        RECT 74.890 40.140 75.080 40.310 ;
        RECT 75.250 40.140 75.280 40.310 ;
        RECT 74.330 38.930 75.280 40.140 ;
      LAYER li1 ;
        RECT 72.260 38.540 74.150 38.710 ;
        RECT 72.260 38.410 72.430 38.540 ;
        RECT 74.930 38.410 75.260 38.750 ;
        RECT 71.170 38.180 72.430 38.410 ;
      LAYER li1 ;
        RECT 72.610 38.230 74.640 38.360 ;
        RECT 75.460 38.230 75.710 40.390 ;
        RECT 76.090 40.360 77.540 40.390 ;
        RECT 76.090 40.190 76.340 40.360 ;
        RECT 76.510 40.190 76.700 40.360 ;
        RECT 76.870 40.190 77.140 40.360 ;
        RECT 77.310 40.190 77.540 40.360 ;
        RECT 76.090 39.320 77.540 40.190 ;
        RECT 72.610 38.190 75.710 38.230 ;
      LAYER li1 ;
        RECT 72.260 38.010 72.430 38.180 ;
      LAYER li1 ;
        RECT 74.470 38.060 75.710 38.190 ;
        RECT 69.600 37.480 70.900 37.880 ;
        RECT 69.290 37.000 70.900 37.480 ;
        RECT 71.130 37.000 72.080 37.960 ;
      LAYER li1 ;
        RECT 72.260 37.840 74.070 38.010 ;
        RECT 72.260 37.130 72.510 37.840 ;
      LAYER li1 ;
        RECT 72.690 37.000 73.640 37.660 ;
      LAYER li1 ;
        RECT 73.820 37.130 74.070 37.840 ;
      LAYER li1 ;
        RECT 74.250 37.000 75.200 37.880 ;
        RECT 75.380 37.130 75.710 38.060 ;
        RECT 76.320 37.880 76.650 38.660 ;
        RECT 76.860 38.330 77.190 39.320 ;
      LAYER li1 ;
        RECT 78.360 38.810 78.790 40.390 ;
      LAYER li1 ;
        RECT 78.970 40.310 79.530 40.390 ;
        RECT 78.970 40.140 78.980 40.310 ;
        RECT 79.150 40.140 79.340 40.310 ;
        RECT 79.510 40.140 79.530 40.310 ;
        RECT 78.970 38.810 79.530 40.140 ;
        RECT 80.890 40.360 82.340 40.390 ;
        RECT 80.890 40.190 81.140 40.360 ;
        RECT 81.310 40.190 81.500 40.360 ;
        RECT 81.670 40.190 81.940 40.360 ;
        RECT 82.110 40.190 82.340 40.360 ;
        RECT 76.320 37.480 77.620 37.880 ;
        RECT 76.010 37.000 77.620 37.480 ;
      LAYER li1 ;
        RECT 78.360 37.130 78.610 38.810 ;
      LAYER li1 ;
        RECT 78.920 37.920 79.250 38.380 ;
      LAYER li1 ;
        RECT 79.710 38.100 80.040 39.890 ;
      LAYER li1 ;
        RECT 80.220 37.920 80.470 39.640 ;
        RECT 80.890 39.320 82.340 40.190 ;
        RECT 82.650 40.310 83.600 40.390 ;
        RECT 82.650 40.140 82.680 40.310 ;
        RECT 82.850 40.140 83.040 40.310 ;
        RECT 83.210 40.140 83.400 40.310 ;
        RECT 83.570 40.140 83.600 40.310 ;
        RECT 78.920 37.750 80.470 37.920 ;
        RECT 78.790 37.000 80.040 37.570 ;
        RECT 80.220 37.130 80.470 37.750 ;
        RECT 81.120 37.880 81.450 38.660 ;
        RECT 81.660 38.330 81.990 39.320 ;
        RECT 82.650 38.810 83.600 40.140 ;
      LAYER li1 ;
        RECT 83.780 38.710 84.030 40.390 ;
      LAYER li1 ;
        RECT 84.210 40.310 85.160 40.390 ;
        RECT 84.210 40.140 84.240 40.310 ;
        RECT 84.410 40.140 84.600 40.310 ;
        RECT 84.770 40.140 84.960 40.310 ;
        RECT 85.130 40.140 85.160 40.310 ;
        RECT 84.210 38.890 85.160 40.140 ;
      LAYER li1 ;
        RECT 85.340 38.710 85.670 40.390 ;
      LAYER li1 ;
        RECT 85.850 40.310 86.800 40.390 ;
        RECT 85.850 40.140 85.880 40.310 ;
        RECT 86.050 40.140 86.240 40.310 ;
        RECT 86.410 40.140 86.600 40.310 ;
        RECT 86.770 40.140 86.800 40.310 ;
        RECT 85.850 38.930 86.800 40.140 ;
      LAYER li1 ;
        RECT 83.780 38.540 85.670 38.710 ;
        RECT 83.780 38.410 83.950 38.540 ;
        RECT 86.450 38.410 86.780 38.750 ;
        RECT 82.690 38.180 83.950 38.410 ;
      LAYER li1 ;
        RECT 84.130 38.230 86.160 38.360 ;
        RECT 86.980 38.230 87.230 40.390 ;
        RECT 87.610 40.360 89.060 40.390 ;
        RECT 87.610 40.190 87.860 40.360 ;
        RECT 88.030 40.190 88.220 40.360 ;
        RECT 88.390 40.190 88.660 40.360 ;
        RECT 88.830 40.190 89.060 40.360 ;
        RECT 87.610 39.320 89.060 40.190 ;
        RECT 89.370 40.310 90.320 40.390 ;
        RECT 89.370 40.140 89.400 40.310 ;
        RECT 89.570 40.140 89.760 40.310 ;
        RECT 89.930 40.140 90.120 40.310 ;
        RECT 90.290 40.140 90.320 40.310 ;
        RECT 84.130 38.190 87.230 38.230 ;
      LAYER li1 ;
        RECT 83.780 38.010 83.950 38.180 ;
      LAYER li1 ;
        RECT 85.990 38.060 87.230 38.190 ;
        RECT 81.120 37.480 82.420 37.880 ;
        RECT 80.810 37.000 82.420 37.480 ;
        RECT 82.650 37.000 83.600 37.960 ;
      LAYER li1 ;
        RECT 83.780 37.840 85.590 38.010 ;
        RECT 83.780 37.130 84.030 37.840 ;
      LAYER li1 ;
        RECT 84.210 37.000 85.160 37.660 ;
      LAYER li1 ;
        RECT 85.340 37.130 85.590 37.840 ;
      LAYER li1 ;
        RECT 85.770 37.000 86.720 37.880 ;
        RECT 86.900 37.130 87.230 38.060 ;
        RECT 87.840 37.880 88.170 38.660 ;
        RECT 88.380 38.330 88.710 39.320 ;
        RECT 89.370 38.810 90.320 40.140 ;
      LAYER li1 ;
        RECT 90.500 38.710 90.750 40.390 ;
      LAYER li1 ;
        RECT 90.930 40.310 91.880 40.390 ;
        RECT 90.930 40.140 90.960 40.310 ;
        RECT 91.130 40.140 91.320 40.310 ;
        RECT 91.490 40.140 91.680 40.310 ;
        RECT 91.850 40.140 91.880 40.310 ;
        RECT 90.930 38.890 91.880 40.140 ;
      LAYER li1 ;
        RECT 92.060 38.710 92.390 40.390 ;
      LAYER li1 ;
        RECT 92.570 40.310 93.520 40.390 ;
        RECT 92.570 40.140 92.600 40.310 ;
        RECT 92.770 40.140 92.960 40.310 ;
        RECT 93.130 40.140 93.320 40.310 ;
        RECT 93.490 40.140 93.520 40.310 ;
        RECT 92.570 38.930 93.520 40.140 ;
      LAYER li1 ;
        RECT 90.500 38.540 92.390 38.710 ;
        RECT 90.500 38.410 90.670 38.540 ;
        RECT 93.170 38.410 93.500 38.750 ;
        RECT 89.410 38.180 90.670 38.410 ;
      LAYER li1 ;
        RECT 90.850 38.230 92.880 38.360 ;
        RECT 93.700 38.230 93.950 40.390 ;
        RECT 94.330 40.360 95.780 40.390 ;
        RECT 94.330 40.190 94.580 40.360 ;
        RECT 94.750 40.190 94.940 40.360 ;
        RECT 95.110 40.190 95.380 40.360 ;
        RECT 95.550 40.190 95.780 40.360 ;
        RECT 94.330 39.320 95.780 40.190 ;
        RECT 96.090 40.310 97.350 40.390 ;
        RECT 96.090 40.140 96.100 40.310 ;
        RECT 96.270 40.140 96.460 40.310 ;
        RECT 96.630 40.140 96.820 40.310 ;
        RECT 96.990 40.140 97.180 40.310 ;
        RECT 90.850 38.190 93.950 38.230 ;
      LAYER li1 ;
        RECT 90.500 38.010 90.670 38.180 ;
      LAYER li1 ;
        RECT 92.710 38.060 93.950 38.190 ;
        RECT 87.840 37.480 89.140 37.880 ;
        RECT 87.530 37.000 89.140 37.480 ;
        RECT 89.370 37.000 90.320 37.960 ;
      LAYER li1 ;
        RECT 90.500 37.840 92.310 38.010 ;
        RECT 90.500 37.130 90.750 37.840 ;
      LAYER li1 ;
        RECT 90.930 37.000 91.880 37.660 ;
      LAYER li1 ;
        RECT 92.060 37.130 92.310 37.840 ;
      LAYER li1 ;
        RECT 92.490 37.000 93.440 37.880 ;
        RECT 93.620 37.130 93.950 38.060 ;
        RECT 94.560 37.880 94.890 38.660 ;
        RECT 95.100 38.330 95.430 39.320 ;
        RECT 96.090 38.910 97.350 40.140 ;
      LAYER li1 ;
        RECT 97.880 39.890 98.050 40.390 ;
        RECT 97.530 38.810 98.050 39.890 ;
      LAYER li1 ;
        RECT 98.310 40.310 99.620 40.390 ;
        RECT 98.310 40.140 98.340 40.310 ;
        RECT 98.510 40.140 98.700 40.310 ;
        RECT 98.870 40.140 99.060 40.310 ;
        RECT 99.230 40.140 99.420 40.310 ;
        RECT 99.590 40.140 99.620 40.310 ;
        RECT 98.310 38.930 99.620 40.140 ;
        RECT 100.090 40.360 101.540 40.390 ;
        RECT 100.090 40.190 100.340 40.360 ;
        RECT 100.510 40.190 100.700 40.360 ;
        RECT 100.870 40.190 101.140 40.360 ;
        RECT 101.310 40.190 101.540 40.360 ;
        RECT 100.090 39.320 101.540 40.190 ;
        RECT 101.850 40.310 103.520 40.390 ;
        RECT 101.850 40.140 101.880 40.310 ;
        RECT 102.050 40.140 102.240 40.310 ;
        RECT 102.410 40.140 102.600 40.310 ;
        RECT 102.770 40.140 102.960 40.310 ;
        RECT 103.130 40.140 103.320 40.310 ;
        RECT 103.490 40.140 103.520 40.310 ;
      LAYER li1 ;
        RECT 97.530 38.730 97.800 38.810 ;
        RECT 96.740 38.560 97.800 38.730 ;
        RECT 96.130 38.170 96.550 38.500 ;
        RECT 96.740 37.990 96.910 38.560 ;
        RECT 98.250 38.440 98.760 38.750 ;
        RECT 99.010 38.440 99.720 38.750 ;
        RECT 97.090 38.170 97.600 38.380 ;
      LAYER li1 ;
        RECT 97.800 38.090 99.670 38.260 ;
        RECT 94.560 37.480 95.860 37.880 ;
        RECT 94.250 37.000 95.860 37.480 ;
        RECT 96.160 37.070 96.490 37.990 ;
      LAYER li1 ;
        RECT 96.740 37.250 97.270 37.990 ;
      LAYER li1 ;
        RECT 97.800 37.070 97.970 38.090 ;
        RECT 96.160 36.900 97.970 37.070 ;
        RECT 98.150 37.000 99.250 37.910 ;
        RECT 99.420 37.160 99.670 38.090 ;
        RECT 100.320 37.880 100.650 38.660 ;
        RECT 100.860 38.330 101.190 39.320 ;
        RECT 101.850 38.930 103.520 40.140 ;
      LAYER li1 ;
        RECT 101.890 38.160 102.190 38.750 ;
        RECT 102.370 38.410 103.560 38.750 ;
        RECT 103.740 38.410 104.070 39.890 ;
        RECT 104.250 38.230 104.520 40.390 ;
      LAYER li1 ;
        RECT 105.370 40.360 106.820 40.390 ;
        RECT 105.370 40.190 105.620 40.360 ;
        RECT 105.790 40.190 105.980 40.360 ;
        RECT 106.150 40.190 106.420 40.360 ;
        RECT 106.590 40.190 106.820 40.360 ;
      LAYER li1 ;
        RECT 102.690 38.060 104.520 38.230 ;
        RECT 104.790 38.210 104.960 39.490 ;
      LAYER li1 ;
        RECT 105.370 39.320 106.820 40.190 ;
        RECT 107.130 40.310 107.720 40.390 ;
        RECT 107.130 40.140 107.160 40.310 ;
        RECT 107.330 40.140 107.520 40.310 ;
        RECT 107.690 40.140 107.720 40.310 ;
        RECT 100.320 37.480 101.620 37.880 ;
        RECT 100.010 37.000 101.620 37.480 ;
        RECT 101.850 37.000 102.440 37.960 ;
      LAYER li1 ;
        RECT 102.690 37.130 102.940 38.060 ;
      LAYER li1 ;
        RECT 103.120 37.000 104.070 37.880 ;
      LAYER li1 ;
        RECT 104.250 37.130 104.520 38.060 ;
      LAYER li1 ;
        RECT 105.600 37.880 105.930 38.660 ;
        RECT 106.140 38.330 106.470 39.320 ;
        RECT 107.130 38.810 107.720 40.140 ;
      LAYER li1 ;
        RECT 108.000 38.810 108.390 40.390 ;
      LAYER li1 ;
        RECT 108.730 40.360 110.180 40.390 ;
        RECT 108.730 40.190 108.980 40.360 ;
        RECT 109.150 40.190 109.340 40.360 ;
        RECT 109.510 40.190 109.780 40.360 ;
        RECT 109.950 40.190 110.180 40.360 ;
        RECT 108.730 39.320 110.180 40.190 ;
        RECT 110.970 40.310 111.920 40.390 ;
        RECT 110.970 40.140 111.000 40.310 ;
        RECT 111.170 40.140 111.360 40.310 ;
        RECT 111.530 40.140 111.720 40.310 ;
        RECT 111.890 40.140 111.920 40.310 ;
      LAYER li1 ;
        RECT 107.170 38.180 107.880 38.570 ;
      LAYER li1 ;
        RECT 105.600 37.480 106.900 37.880 ;
        RECT 105.290 37.000 106.900 37.480 ;
        RECT 107.130 37.000 107.720 37.960 ;
      LAYER li1 ;
        RECT 108.060 37.130 108.390 38.810 ;
      LAYER li1 ;
        RECT 108.960 37.880 109.290 38.660 ;
        RECT 109.500 38.330 109.830 39.320 ;
        RECT 110.970 38.810 111.920 40.140 ;
      LAYER li1 ;
        RECT 112.100 38.710 112.350 40.390 ;
      LAYER li1 ;
        RECT 112.530 40.310 113.480 40.390 ;
        RECT 112.530 40.140 112.560 40.310 ;
        RECT 112.730 40.140 112.920 40.310 ;
        RECT 113.090 40.140 113.280 40.310 ;
        RECT 113.450 40.140 113.480 40.310 ;
        RECT 112.530 38.890 113.480 40.140 ;
      LAYER li1 ;
        RECT 113.660 38.710 113.990 40.390 ;
      LAYER li1 ;
        RECT 114.170 40.310 115.120 40.390 ;
        RECT 114.170 40.140 114.200 40.310 ;
        RECT 114.370 40.140 114.560 40.310 ;
        RECT 114.730 40.140 114.920 40.310 ;
        RECT 115.090 40.140 115.120 40.310 ;
        RECT 114.170 38.930 115.120 40.140 ;
      LAYER li1 ;
        RECT 112.100 38.540 113.990 38.710 ;
        RECT 112.100 38.410 112.270 38.540 ;
        RECT 114.770 38.410 115.100 38.750 ;
        RECT 111.010 38.180 112.270 38.410 ;
      LAYER li1 ;
        RECT 112.450 38.230 114.480 38.360 ;
        RECT 115.300 38.230 115.550 40.390 ;
        RECT 116.180 40.360 118.920 40.380 ;
        RECT 116.180 40.190 116.390 40.360 ;
        RECT 116.560 40.190 116.830 40.360 ;
        RECT 117.000 40.190 117.240 40.360 ;
        RECT 117.410 40.190 117.670 40.360 ;
        RECT 117.840 40.190 118.110 40.360 ;
        RECT 118.280 40.190 118.520 40.360 ;
        RECT 118.690 40.190 118.920 40.360 ;
        RECT 116.180 39.310 118.920 40.190 ;
        RECT 120.570 40.310 121.520 40.390 ;
        RECT 120.570 40.140 120.600 40.310 ;
        RECT 120.770 40.140 120.960 40.310 ;
        RECT 121.130 40.140 121.320 40.310 ;
        RECT 121.490 40.140 121.520 40.310 ;
        RECT 112.450 38.190 115.550 38.230 ;
      LAYER li1 ;
        RECT 112.100 38.010 112.270 38.180 ;
      LAYER li1 ;
        RECT 114.310 38.060 115.550 38.190 ;
        RECT 108.960 37.480 110.260 37.880 ;
        RECT 108.650 37.000 110.260 37.480 ;
        RECT 110.970 37.000 111.920 37.960 ;
      LAYER li1 ;
        RECT 112.100 37.840 113.910 38.010 ;
        RECT 112.100 37.130 112.350 37.840 ;
      LAYER li1 ;
        RECT 112.530 37.000 113.480 37.660 ;
      LAYER li1 ;
        RECT 113.660 37.130 113.910 37.840 ;
      LAYER li1 ;
        RECT 114.090 37.000 115.040 37.880 ;
        RECT 115.220 37.130 115.550 38.060 ;
        RECT 116.420 37.990 116.750 38.660 ;
        RECT 117.150 38.330 117.480 39.310 ;
        RECT 117.700 37.990 118.030 38.660 ;
        RECT 118.430 38.330 118.760 39.310 ;
        RECT 120.570 38.810 121.520 40.140 ;
      LAYER li1 ;
        RECT 121.700 38.710 121.950 40.390 ;
      LAYER li1 ;
        RECT 122.130 40.310 123.080 40.390 ;
        RECT 122.130 40.140 122.160 40.310 ;
        RECT 122.330 40.140 122.520 40.310 ;
        RECT 122.690 40.140 122.880 40.310 ;
        RECT 123.050 40.140 123.080 40.310 ;
        RECT 122.130 38.890 123.080 40.140 ;
      LAYER li1 ;
        RECT 123.260 38.710 123.590 40.390 ;
      LAYER li1 ;
        RECT 123.770 40.310 124.720 40.390 ;
        RECT 123.770 40.140 123.800 40.310 ;
        RECT 123.970 40.140 124.160 40.310 ;
        RECT 124.330 40.140 124.520 40.310 ;
        RECT 124.690 40.140 124.720 40.310 ;
        RECT 123.770 38.930 124.720 40.140 ;
      LAYER li1 ;
        RECT 121.700 38.540 123.590 38.710 ;
        RECT 121.700 38.410 121.870 38.540 ;
        RECT 124.370 38.410 124.700 38.750 ;
        RECT 120.610 38.180 121.870 38.410 ;
      LAYER li1 ;
        RECT 122.050 38.230 124.080 38.360 ;
        RECT 124.900 38.230 125.150 40.390 ;
        RECT 125.530 40.360 126.980 40.390 ;
        RECT 125.530 40.190 125.780 40.360 ;
        RECT 125.950 40.190 126.140 40.360 ;
        RECT 126.310 40.190 126.580 40.360 ;
        RECT 126.750 40.190 126.980 40.360 ;
        RECT 125.530 39.320 126.980 40.190 ;
        RECT 122.050 38.190 125.150 38.230 ;
      LAYER li1 ;
        RECT 121.700 38.010 121.870 38.180 ;
      LAYER li1 ;
        RECT 123.910 38.060 125.150 38.190 ;
        RECT 116.260 36.990 118.990 37.990 ;
        RECT 120.570 37.000 121.520 37.960 ;
      LAYER li1 ;
        RECT 121.700 37.840 123.510 38.010 ;
        RECT 121.700 37.130 121.950 37.840 ;
      LAYER li1 ;
        RECT 122.130 37.000 123.080 37.660 ;
      LAYER li1 ;
        RECT 123.260 37.130 123.510 37.840 ;
      LAYER li1 ;
        RECT 123.690 37.000 124.640 37.880 ;
        RECT 124.820 37.130 125.150 38.060 ;
        RECT 125.760 37.880 126.090 38.660 ;
        RECT 126.300 38.330 126.630 39.320 ;
      LAYER li1 ;
        RECT 127.330 38.610 127.800 40.390 ;
      LAYER li1 ;
        RECT 127.980 40.310 129.230 40.390 ;
        RECT 128.150 40.140 128.340 40.310 ;
        RECT 128.510 40.140 128.700 40.310 ;
        RECT 128.870 40.140 129.060 40.310 ;
        RECT 127.980 38.930 129.230 40.140 ;
        RECT 125.760 37.480 127.060 37.880 ;
        RECT 125.450 37.000 127.060 37.480 ;
      LAYER li1 ;
        RECT 127.330 37.160 127.580 38.610 ;
        RECT 128.290 38.440 129.200 38.750 ;
      LAYER li1 ;
        RECT 127.750 38.260 128.040 38.430 ;
        RECT 129.410 38.260 129.580 40.390 ;
        RECT 130.170 40.310 131.430 40.390 ;
        RECT 130.340 40.140 130.530 40.310 ;
        RECT 130.700 40.140 130.890 40.310 ;
        RECT 131.060 40.140 131.250 40.310 ;
        RECT 131.420 40.140 131.430 40.310 ;
      LAYER li1 ;
        RECT 129.760 39.860 129.990 39.890 ;
        RECT 129.750 39.690 129.990 39.860 ;
      LAYER li1 ;
        RECT 127.750 38.090 129.580 38.260 ;
      LAYER li1 ;
        RECT 129.760 38.180 129.990 39.690 ;
      LAYER li1 ;
        RECT 130.170 38.810 131.430 40.140 ;
        RECT 131.770 40.360 133.220 40.390 ;
        RECT 131.770 40.190 132.020 40.360 ;
        RECT 132.190 40.190 132.380 40.360 ;
        RECT 132.550 40.190 132.820 40.360 ;
        RECT 132.990 40.190 133.220 40.360 ;
        RECT 131.770 39.320 133.220 40.190 ;
      LAYER li1 ;
        RECT 130.210 38.140 131.400 38.470 ;
      LAYER li1 ;
        RECT 127.750 37.000 128.520 37.910 ;
        RECT 128.700 37.130 129.030 38.090 ;
        RECT 131.060 37.910 131.390 37.960 ;
        RECT 129.480 37.740 131.390 37.910 ;
        RECT 129.480 37.130 129.810 37.740 ;
        RECT 129.990 37.000 130.880 37.560 ;
        RECT 131.060 37.130 131.390 37.740 ;
        RECT 132.000 37.880 132.330 38.660 ;
        RECT 132.540 38.330 132.870 39.320 ;
      LAYER li1 ;
        RECT 133.560 38.810 133.990 40.390 ;
      LAYER li1 ;
        RECT 134.170 40.310 134.730 40.390 ;
        RECT 134.170 40.140 134.180 40.310 ;
        RECT 134.350 40.140 134.540 40.310 ;
        RECT 134.710 40.140 134.730 40.310 ;
        RECT 134.170 38.810 134.730 40.140 ;
        RECT 136.090 40.360 137.540 40.390 ;
        RECT 136.090 40.190 136.340 40.360 ;
        RECT 136.510 40.190 136.700 40.360 ;
        RECT 136.870 40.190 137.140 40.360 ;
        RECT 137.310 40.190 137.540 40.360 ;
        RECT 132.000 37.480 133.300 37.880 ;
        RECT 131.690 37.000 133.300 37.480 ;
      LAYER li1 ;
        RECT 133.560 37.130 133.810 38.810 ;
      LAYER li1 ;
        RECT 134.120 37.920 134.450 38.380 ;
      LAYER li1 ;
        RECT 134.910 38.100 135.240 39.890 ;
      LAYER li1 ;
        RECT 135.420 37.920 135.670 39.640 ;
        RECT 136.090 39.320 137.540 40.190 ;
        RECT 137.980 40.310 138.630 40.420 ;
        RECT 137.980 40.140 138.040 40.310 ;
        RECT 138.210 40.140 138.400 40.310 ;
        RECT 138.570 40.140 138.630 40.310 ;
        RECT 137.980 40.080 138.630 40.140 ;
        RECT 137.980 39.810 138.380 40.080 ;
      LAYER li1 ;
        RECT 139.290 39.810 139.870 40.450 ;
      LAYER li1 ;
        RECT 140.410 40.360 141.860 40.390 ;
        RECT 140.410 40.190 140.660 40.360 ;
        RECT 140.830 40.190 141.020 40.360 ;
        RECT 141.190 40.190 141.460 40.360 ;
        RECT 141.630 40.190 141.860 40.360 ;
        RECT 134.120 37.750 135.670 37.920 ;
        RECT 133.990 37.000 135.240 37.570 ;
        RECT 135.420 37.130 135.670 37.750 ;
        RECT 136.320 37.880 136.650 38.660 ;
        RECT 136.860 38.330 137.190 39.320 ;
      LAYER li1 ;
        RECT 139.290 38.400 139.560 39.810 ;
      LAYER li1 ;
        RECT 140.410 39.320 141.860 40.190 ;
      LAYER li1 ;
        RECT 138.800 38.130 139.560 38.400 ;
      LAYER li1 ;
        RECT 136.320 37.480 137.620 37.880 ;
        RECT 136.010 37.000 137.620 37.480 ;
      LAYER li1 ;
        RECT 138.800 37.130 139.130 38.130 ;
      LAYER li1 ;
        RECT 140.640 37.880 140.970 38.660 ;
        RECT 141.180 38.330 141.510 39.320 ;
        RECT 139.540 37.260 139.950 37.700 ;
        RECT 140.640 37.480 141.940 37.880 ;
        RECT 139.300 36.920 139.950 37.260 ;
        RECT 140.330 37.000 141.940 37.480 ;
        RECT 5.760 36.540 5.920 36.720 ;
        RECT 6.090 36.540 6.400 36.720 ;
        RECT 6.570 36.540 6.880 36.720 ;
        RECT 7.050 36.540 7.360 36.720 ;
        RECT 7.530 36.540 7.840 36.720 ;
        RECT 8.010 36.540 8.320 36.720 ;
        RECT 8.490 36.540 8.800 36.720 ;
        RECT 8.970 36.540 9.280 36.720 ;
        RECT 9.450 36.540 9.760 36.720 ;
        RECT 9.930 36.540 10.240 36.720 ;
        RECT 10.410 36.540 10.720 36.720 ;
        RECT 10.890 36.540 11.200 36.720 ;
        RECT 11.370 36.540 11.680 36.720 ;
        RECT 11.850 36.540 12.160 36.720 ;
        RECT 12.330 36.540 12.640 36.720 ;
        RECT 12.810 36.540 13.120 36.720 ;
        RECT 13.290 36.540 13.600 36.720 ;
        RECT 13.770 36.540 14.080 36.720 ;
        RECT 14.250 36.540 14.400 36.720 ;
        RECT 14.880 36.540 15.040 36.720 ;
        RECT 15.210 36.540 15.520 36.720 ;
        RECT 15.690 36.540 16.000 36.720 ;
        RECT 16.170 36.540 16.480 36.720 ;
        RECT 16.650 36.540 16.960 36.720 ;
        RECT 17.130 36.540 17.440 36.720 ;
        RECT 17.610 36.540 17.920 36.720 ;
        RECT 18.090 36.540 18.400 36.720 ;
        RECT 18.570 36.540 18.880 36.720 ;
        RECT 19.050 36.540 19.360 36.720 ;
        RECT 19.530 36.540 19.840 36.720 ;
        RECT 20.010 36.540 20.320 36.720 ;
        RECT 20.490 36.540 20.800 36.720 ;
        RECT 20.970 36.540 21.280 36.720 ;
        RECT 21.450 36.540 21.760 36.720 ;
        RECT 21.930 36.540 22.240 36.720 ;
        RECT 22.410 36.540 22.720 36.720 ;
        RECT 22.890 36.540 23.200 36.720 ;
        RECT 23.370 36.540 23.680 36.720 ;
        RECT 23.850 36.540 24.160 36.720 ;
        RECT 24.330 36.540 24.640 36.720 ;
        RECT 24.810 36.540 25.120 36.720 ;
        RECT 25.290 36.540 25.600 36.720 ;
        RECT 25.770 36.540 26.080 36.720 ;
        RECT 26.250 36.540 26.560 36.720 ;
        RECT 26.730 36.540 27.040 36.720 ;
        RECT 27.210 36.540 27.520 36.720 ;
        RECT 27.690 36.540 28.000 36.720 ;
        RECT 28.170 36.540 28.480 36.720 ;
        RECT 28.650 36.540 28.960 36.720 ;
        RECT 29.130 36.540 29.440 36.720 ;
        RECT 29.610 36.540 29.920 36.720 ;
        RECT 30.090 36.540 30.400 36.720 ;
        RECT 30.570 36.540 30.880 36.720 ;
        RECT 31.050 36.540 31.360 36.720 ;
        RECT 31.530 36.540 31.840 36.720 ;
        RECT 32.010 36.540 32.320 36.720 ;
        RECT 32.490 36.540 32.800 36.720 ;
        RECT 32.970 36.540 33.280 36.720 ;
        RECT 33.450 36.540 33.760 36.720 ;
        RECT 33.930 36.540 34.240 36.720 ;
        RECT 34.410 36.540 34.720 36.720 ;
        RECT 34.890 36.540 35.200 36.720 ;
        RECT 35.370 36.540 35.680 36.720 ;
        RECT 35.850 36.540 36.160 36.720 ;
        RECT 36.330 36.540 36.640 36.720 ;
        RECT 36.810 36.540 37.120 36.720 ;
        RECT 37.290 36.540 37.600 36.720 ;
        RECT 37.770 36.540 38.080 36.720 ;
        RECT 38.250 36.540 38.560 36.720 ;
        RECT 38.730 36.540 39.040 36.720 ;
        RECT 39.210 36.540 39.520 36.720 ;
        RECT 39.690 36.540 40.000 36.720 ;
        RECT 40.170 36.540 40.480 36.720 ;
        RECT 40.650 36.540 40.960 36.720 ;
        RECT 41.130 36.540 41.440 36.720 ;
        RECT 41.610 36.540 41.920 36.720 ;
        RECT 42.090 36.540 42.400 36.720 ;
        RECT 42.570 36.540 42.880 36.720 ;
        RECT 43.050 36.540 43.360 36.720 ;
        RECT 43.530 36.540 43.840 36.720 ;
        RECT 44.010 36.540 44.320 36.720 ;
        RECT 44.490 36.540 44.800 36.720 ;
        RECT 44.970 36.540 45.280 36.720 ;
        RECT 45.450 36.540 45.760 36.720 ;
        RECT 45.930 36.540 46.240 36.720 ;
        RECT 46.410 36.540 46.720 36.720 ;
        RECT 46.890 36.540 47.200 36.720 ;
        RECT 47.370 36.540 47.680 36.720 ;
        RECT 47.850 36.540 48.160 36.720 ;
        RECT 48.330 36.540 48.640 36.720 ;
        RECT 48.810 36.540 49.120 36.720 ;
        RECT 49.290 36.540 49.600 36.720 ;
        RECT 49.770 36.540 50.080 36.720 ;
        RECT 50.250 36.540 50.560 36.720 ;
        RECT 50.730 36.540 51.040 36.720 ;
        RECT 51.210 36.540 51.520 36.720 ;
        RECT 51.690 36.540 52.000 36.720 ;
        RECT 52.170 36.540 52.480 36.720 ;
        RECT 52.650 36.540 52.960 36.720 ;
        RECT 53.130 36.540 53.440 36.720 ;
        RECT 53.610 36.540 53.920 36.720 ;
        RECT 54.090 36.540 54.400 36.720 ;
        RECT 54.570 36.540 54.880 36.720 ;
        RECT 55.050 36.540 55.360 36.720 ;
        RECT 55.530 36.540 55.840 36.720 ;
        RECT 56.010 36.540 56.320 36.720 ;
        RECT 56.490 36.540 56.800 36.720 ;
        RECT 56.970 36.540 57.280 36.720 ;
        RECT 57.450 36.540 57.760 36.720 ;
        RECT 57.930 36.540 58.240 36.720 ;
        RECT 58.410 36.540 58.720 36.720 ;
        RECT 58.890 36.540 59.200 36.720 ;
        RECT 59.370 36.540 59.680 36.720 ;
        RECT 59.850 36.540 60.160 36.720 ;
        RECT 60.330 36.540 60.640 36.720 ;
        RECT 60.810 36.540 61.120 36.720 ;
        RECT 61.290 36.540 61.600 36.720 ;
        RECT 61.770 36.540 62.080 36.720 ;
        RECT 62.250 36.540 62.560 36.720 ;
        RECT 62.730 36.540 63.040 36.720 ;
        RECT 63.210 36.540 63.520 36.720 ;
        RECT 63.690 36.540 64.000 36.720 ;
        RECT 64.170 36.540 64.480 36.720 ;
        RECT 64.650 36.540 64.960 36.720 ;
        RECT 65.130 36.540 65.440 36.720 ;
        RECT 65.610 36.540 65.920 36.720 ;
        RECT 66.090 36.540 66.400 36.720 ;
        RECT 66.570 36.540 66.880 36.720 ;
        RECT 67.050 36.540 67.360 36.720 ;
        RECT 67.530 36.540 67.840 36.720 ;
        RECT 68.010 36.540 68.320 36.720 ;
        RECT 68.490 36.540 68.800 36.720 ;
        RECT 68.970 36.540 69.280 36.720 ;
        RECT 69.450 36.540 69.760 36.720 ;
        RECT 69.930 36.540 70.240 36.720 ;
        RECT 70.410 36.540 70.720 36.720 ;
        RECT 70.890 36.540 71.200 36.720 ;
        RECT 71.370 36.540 71.680 36.720 ;
        RECT 71.850 36.540 72.160 36.720 ;
        RECT 72.330 36.540 72.640 36.720 ;
        RECT 72.810 36.540 73.120 36.720 ;
        RECT 73.290 36.540 73.600 36.720 ;
        RECT 73.770 36.540 74.080 36.720 ;
        RECT 74.250 36.540 74.560 36.720 ;
        RECT 74.730 36.540 75.040 36.720 ;
        RECT 75.210 36.540 75.520 36.720 ;
        RECT 75.690 36.540 76.000 36.720 ;
        RECT 76.170 36.540 76.480 36.720 ;
        RECT 76.650 36.540 76.960 36.720 ;
        RECT 77.130 36.540 77.440 36.720 ;
        RECT 77.610 36.540 77.760 36.720 ;
        RECT 78.240 36.540 78.400 36.720 ;
        RECT 78.570 36.540 78.880 36.720 ;
        RECT 79.050 36.540 79.360 36.720 ;
        RECT 79.530 36.540 79.840 36.720 ;
        RECT 80.010 36.540 80.320 36.720 ;
        RECT 80.490 36.540 80.800 36.720 ;
        RECT 80.970 36.540 81.280 36.720 ;
        RECT 81.450 36.540 81.760 36.720 ;
        RECT 81.930 36.540 82.240 36.720 ;
        RECT 82.410 36.540 82.720 36.720 ;
        RECT 82.890 36.540 83.200 36.720 ;
        RECT 83.370 36.540 83.680 36.720 ;
        RECT 83.850 36.540 84.160 36.720 ;
        RECT 84.330 36.540 84.640 36.720 ;
        RECT 84.810 36.540 85.120 36.720 ;
        RECT 85.290 36.540 85.600 36.720 ;
        RECT 85.770 36.540 86.080 36.720 ;
        RECT 86.250 36.540 86.560 36.720 ;
        RECT 86.730 36.540 87.040 36.720 ;
        RECT 87.210 36.540 87.520 36.720 ;
        RECT 87.690 36.540 88.000 36.720 ;
        RECT 88.170 36.540 88.480 36.720 ;
        RECT 88.650 36.540 88.960 36.720 ;
        RECT 89.130 36.540 89.440 36.720 ;
        RECT 89.610 36.540 89.920 36.720 ;
        RECT 90.090 36.540 90.400 36.720 ;
        RECT 90.570 36.540 90.880 36.720 ;
        RECT 91.050 36.540 91.360 36.720 ;
        RECT 91.530 36.540 91.840 36.720 ;
        RECT 92.010 36.540 92.320 36.720 ;
        RECT 92.490 36.540 92.800 36.720 ;
        RECT 92.970 36.540 93.280 36.720 ;
        RECT 93.450 36.540 93.760 36.720 ;
        RECT 93.930 36.540 94.240 36.720 ;
        RECT 94.410 36.540 94.720 36.720 ;
        RECT 94.890 36.540 95.200 36.720 ;
        RECT 95.370 36.540 95.680 36.720 ;
        RECT 95.850 36.540 96.160 36.720 ;
        RECT 96.330 36.540 96.640 36.720 ;
        RECT 96.810 36.540 97.120 36.720 ;
        RECT 97.290 36.540 97.600 36.720 ;
        RECT 97.770 36.540 98.080 36.720 ;
        RECT 98.250 36.540 98.560 36.720 ;
        RECT 98.730 36.540 99.040 36.720 ;
        RECT 99.210 36.540 99.520 36.720 ;
        RECT 99.690 36.540 100.000 36.720 ;
        RECT 100.170 36.540 100.480 36.720 ;
        RECT 100.650 36.540 100.960 36.720 ;
        RECT 101.130 36.540 101.440 36.720 ;
        RECT 101.610 36.540 101.920 36.720 ;
        RECT 102.090 36.540 102.400 36.720 ;
        RECT 102.570 36.540 102.880 36.720 ;
        RECT 103.050 36.540 103.360 36.720 ;
        RECT 103.530 36.540 103.840 36.720 ;
        RECT 104.010 36.540 104.320 36.720 ;
        RECT 104.490 36.540 104.800 36.720 ;
        RECT 104.970 36.540 105.280 36.720 ;
        RECT 105.450 36.540 105.760 36.720 ;
        RECT 105.930 36.540 106.240 36.720 ;
        RECT 106.410 36.540 106.720 36.720 ;
        RECT 106.890 36.540 107.200 36.720 ;
        RECT 107.370 36.540 107.680 36.720 ;
        RECT 107.850 36.540 108.160 36.720 ;
        RECT 108.330 36.540 108.640 36.720 ;
        RECT 108.810 36.540 109.120 36.720 ;
        RECT 109.290 36.540 109.600 36.720 ;
        RECT 109.770 36.540 110.080 36.720 ;
        RECT 110.250 36.540 110.400 36.720 ;
        RECT 110.880 36.540 111.040 36.720 ;
        RECT 111.210 36.540 111.520 36.720 ;
        RECT 111.690 36.540 112.000 36.720 ;
        RECT 112.170 36.540 112.480 36.720 ;
        RECT 112.650 36.540 112.960 36.720 ;
        RECT 113.130 36.540 113.440 36.720 ;
        RECT 113.610 36.540 113.920 36.720 ;
        RECT 114.090 36.540 114.400 36.720 ;
        RECT 114.570 36.540 114.880 36.720 ;
        RECT 115.050 36.540 115.360 36.720 ;
        RECT 115.530 36.540 115.840 36.720 ;
        RECT 116.010 36.540 116.320 36.720 ;
        RECT 116.490 36.540 116.800 36.720 ;
        RECT 116.970 36.540 117.280 36.720 ;
        RECT 117.450 36.540 117.760 36.720 ;
        RECT 117.930 36.540 118.240 36.720 ;
        RECT 118.410 36.540 118.720 36.720 ;
        RECT 118.890 36.540 119.200 36.720 ;
        RECT 119.370 36.540 119.680 36.720 ;
        RECT 119.850 36.540 120.160 36.720 ;
        RECT 120.330 36.540 120.640 36.720 ;
        RECT 120.810 36.540 121.120 36.720 ;
        RECT 121.290 36.540 121.600 36.720 ;
        RECT 121.770 36.540 122.080 36.720 ;
        RECT 122.250 36.540 122.560 36.720 ;
        RECT 122.730 36.540 123.040 36.720 ;
        RECT 123.210 36.540 123.520 36.720 ;
        RECT 123.690 36.540 124.000 36.720 ;
        RECT 124.170 36.540 124.480 36.720 ;
        RECT 124.650 36.540 124.960 36.720 ;
        RECT 125.130 36.540 125.440 36.720 ;
        RECT 125.610 36.540 125.920 36.720 ;
        RECT 126.090 36.540 126.400 36.720 ;
        RECT 126.570 36.540 126.880 36.720 ;
        RECT 127.050 36.540 127.360 36.720 ;
        RECT 127.530 36.540 127.840 36.720 ;
        RECT 128.010 36.540 128.320 36.720 ;
        RECT 128.490 36.540 128.800 36.720 ;
        RECT 128.970 36.540 129.280 36.720 ;
        RECT 129.450 36.540 129.760 36.720 ;
        RECT 129.930 36.540 130.240 36.720 ;
        RECT 130.410 36.540 130.720 36.720 ;
        RECT 130.890 36.540 131.200 36.720 ;
        RECT 131.370 36.540 131.680 36.720 ;
        RECT 131.850 36.540 132.160 36.720 ;
        RECT 132.330 36.540 132.640 36.720 ;
        RECT 132.810 36.540 133.120 36.720 ;
        RECT 133.290 36.540 133.600 36.720 ;
        RECT 133.770 36.540 134.080 36.720 ;
        RECT 134.250 36.540 134.560 36.720 ;
        RECT 134.730 36.540 135.040 36.720 ;
        RECT 135.210 36.540 135.520 36.720 ;
        RECT 135.690 36.540 136.000 36.720 ;
        RECT 136.170 36.540 136.480 36.720 ;
        RECT 136.650 36.540 136.960 36.720 ;
        RECT 137.130 36.540 137.440 36.720 ;
        RECT 137.610 36.540 137.920 36.720 ;
        RECT 138.090 36.540 138.400 36.720 ;
        RECT 138.570 36.540 138.880 36.720 ;
        RECT 139.050 36.540 139.360 36.720 ;
        RECT 139.530 36.540 139.840 36.720 ;
        RECT 140.010 36.540 140.320 36.720 ;
        RECT 140.490 36.540 140.800 36.720 ;
        RECT 140.970 36.540 141.280 36.720 ;
        RECT 141.450 36.540 141.760 36.720 ;
        RECT 141.930 36.540 142.080 36.720 ;
        RECT 6.340 36.240 9.070 36.270 ;
        RECT 6.340 36.070 6.510 36.240 ;
        RECT 6.680 36.070 6.950 36.240 ;
        RECT 7.120 36.070 7.360 36.240 ;
        RECT 7.530 36.070 7.790 36.240 ;
        RECT 7.960 36.070 8.230 36.240 ;
        RECT 8.400 36.070 8.640 36.240 ;
        RECT 8.810 36.070 9.070 36.240 ;
        RECT 6.340 35.270 9.070 36.070 ;
        RECT 10.650 36.230 11.240 36.260 ;
        RECT 10.650 36.060 10.680 36.230 ;
        RECT 10.850 36.060 11.040 36.230 ;
        RECT 11.210 36.060 11.240 36.230 ;
        RECT 12.170 36.230 13.780 36.260 ;
        RECT 14.470 36.230 15.720 36.260 ;
        RECT 16.900 36.240 19.630 36.270 ;
        RECT 10.650 35.300 11.240 36.060 ;
        RECT 6.500 34.600 6.830 35.270 ;
        RECT 7.230 33.950 7.560 34.930 ;
        RECT 7.780 34.600 8.110 35.270 ;
        RECT 8.510 33.950 8.840 34.930 ;
      LAYER li1 ;
        RECT 10.690 34.690 11.400 35.080 ;
        RECT 11.580 34.450 11.910 36.130 ;
      LAYER li1 ;
        RECT 12.170 36.060 12.220 36.230 ;
        RECT 12.390 36.060 12.660 36.230 ;
        RECT 12.830 36.060 13.100 36.230 ;
        RECT 13.270 36.060 13.510 36.230 ;
        RECT 13.680 36.060 13.780 36.230 ;
        RECT 12.170 35.780 13.780 36.060 ;
        RECT 12.480 35.380 13.780 35.780 ;
        RECT 12.480 34.600 12.810 35.380 ;
        RECT 6.260 33.070 9.000 33.950 ;
        RECT 6.260 32.900 6.470 33.070 ;
        RECT 6.640 32.900 6.910 33.070 ;
        RECT 7.080 32.900 7.320 33.070 ;
        RECT 7.490 32.900 7.750 33.070 ;
        RECT 7.920 32.900 8.190 33.070 ;
        RECT 8.360 32.900 8.600 33.070 ;
        RECT 8.770 32.900 9.000 33.070 ;
        RECT 6.260 32.880 9.000 32.900 ;
        RECT 10.650 33.120 11.240 34.450 ;
        RECT 10.650 32.950 10.680 33.120 ;
        RECT 10.850 32.950 11.040 33.120 ;
        RECT 11.210 32.950 11.240 33.120 ;
        RECT 10.650 32.870 11.240 32.950 ;
      LAYER li1 ;
        RECT 11.520 32.870 11.910 34.450 ;
      LAYER li1 ;
        RECT 13.020 33.940 13.350 34.930 ;
      LAYER li1 ;
        RECT 14.040 34.450 14.290 36.130 ;
      LAYER li1 ;
        RECT 14.640 36.060 14.830 36.230 ;
        RECT 15.000 36.060 15.190 36.230 ;
        RECT 15.360 36.060 15.550 36.230 ;
        RECT 14.470 35.690 15.720 36.060 ;
        RECT 15.900 35.510 16.150 36.130 ;
        RECT 14.600 35.340 16.150 35.510 ;
        RECT 14.600 34.880 14.930 35.340 ;
        RECT 12.250 33.070 13.700 33.940 ;
        RECT 12.250 32.900 12.500 33.070 ;
        RECT 12.670 32.900 12.860 33.070 ;
        RECT 13.030 32.900 13.300 33.070 ;
        RECT 13.470 32.900 13.700 33.070 ;
        RECT 12.250 32.870 13.700 32.900 ;
      LAYER li1 ;
        RECT 14.040 32.870 14.470 34.450 ;
      LAYER li1 ;
        RECT 14.650 33.120 15.210 34.450 ;
      LAYER li1 ;
        RECT 15.390 33.370 15.720 35.160 ;
      LAYER li1 ;
        RECT 15.900 33.620 16.150 35.340 ;
        RECT 16.900 36.070 17.070 36.240 ;
        RECT 17.240 36.070 17.510 36.240 ;
        RECT 17.680 36.070 17.920 36.240 ;
        RECT 18.090 36.070 18.350 36.240 ;
        RECT 18.520 36.070 18.790 36.240 ;
        RECT 18.960 36.070 19.200 36.240 ;
        RECT 19.370 36.070 19.630 36.240 ;
        RECT 16.900 35.270 19.630 36.070 ;
        RECT 21.210 36.230 22.520 36.260 ;
        RECT 21.210 36.060 21.240 36.230 ;
        RECT 21.410 36.060 21.600 36.230 ;
        RECT 21.770 36.060 21.960 36.230 ;
        RECT 22.130 36.060 22.320 36.230 ;
        RECT 22.490 36.060 22.520 36.230 ;
        RECT 23.690 36.230 25.300 36.260 ;
        RECT 21.210 35.280 22.520 36.060 ;
      LAYER li1 ;
        RECT 22.970 35.450 23.300 36.110 ;
      LAYER li1 ;
        RECT 23.690 36.060 23.740 36.230 ;
        RECT 23.910 36.060 24.180 36.230 ;
        RECT 24.350 36.060 24.620 36.230 ;
        RECT 24.790 36.060 25.030 36.230 ;
        RECT 25.200 36.060 25.300 36.230 ;
        RECT 23.690 35.780 25.300 36.060 ;
      LAYER li1 ;
        RECT 22.700 35.280 23.300 35.450 ;
      LAYER li1 ;
        RECT 24.000 35.380 25.300 35.780 ;
        RECT 25.600 36.190 27.410 36.360 ;
        RECT 17.060 34.600 17.390 35.270 ;
        RECT 17.790 33.950 18.120 34.930 ;
        RECT 18.340 34.600 18.670 35.270 ;
      LAYER li1 ;
        RECT 22.700 35.100 22.920 35.280 ;
      LAYER li1 ;
        RECT 19.070 33.950 19.400 34.930 ;
      LAYER li1 ;
        RECT 21.250 34.690 22.140 35.080 ;
        RECT 22.340 34.930 22.920 35.100 ;
      LAYER li1 ;
        RECT 14.650 32.950 14.660 33.120 ;
        RECT 14.830 32.950 15.020 33.120 ;
        RECT 15.190 32.950 15.210 33.120 ;
        RECT 14.650 32.870 15.210 32.950 ;
        RECT 16.820 33.070 19.560 33.950 ;
        RECT 16.820 32.900 17.030 33.070 ;
        RECT 17.200 32.900 17.470 33.070 ;
        RECT 17.640 32.900 17.880 33.070 ;
        RECT 18.050 32.900 18.310 33.070 ;
        RECT 18.480 32.900 18.750 33.070 ;
        RECT 18.920 32.900 19.160 33.070 ;
        RECT 19.330 32.900 19.560 33.070 ;
        RECT 16.820 32.880 19.560 32.900 ;
        RECT 21.210 33.120 22.160 34.450 ;
        RECT 21.210 32.950 21.240 33.120 ;
        RECT 21.410 32.950 21.600 33.120 ;
        RECT 21.770 32.950 21.960 33.120 ;
        RECT 22.130 32.950 22.160 33.120 ;
        RECT 21.210 32.870 22.160 32.950 ;
      LAYER li1 ;
        RECT 22.340 32.870 22.590 34.930 ;
        RECT 23.100 34.770 23.400 35.100 ;
      LAYER li1 ;
        RECT 24.000 34.600 24.330 35.380 ;
        RECT 25.600 35.270 25.930 36.190 ;
      LAYER li1 ;
        RECT 26.180 35.270 26.710 36.010 ;
      LAYER li1 ;
        RECT 22.780 33.120 23.370 34.450 ;
        RECT 24.540 33.940 24.870 34.930 ;
      LAYER li1 ;
        RECT 25.570 34.760 25.990 35.090 ;
        RECT 26.180 34.700 26.350 35.270 ;
      LAYER li1 ;
        RECT 27.240 35.170 27.410 36.190 ;
        RECT 27.590 36.230 28.690 36.260 ;
        RECT 27.590 36.060 27.640 36.230 ;
        RECT 27.810 36.060 28.000 36.230 ;
        RECT 28.170 36.060 28.360 36.230 ;
        RECT 28.530 36.060 28.690 36.230 ;
        RECT 29.450 36.230 31.060 36.260 ;
        RECT 31.760 36.230 32.650 36.260 ;
        RECT 27.590 35.350 28.690 36.060 ;
        RECT 28.860 35.170 29.110 36.100 ;
        RECT 29.450 36.060 29.500 36.230 ;
        RECT 29.670 36.060 29.940 36.230 ;
        RECT 30.110 36.060 30.380 36.230 ;
        RECT 30.550 36.060 30.790 36.230 ;
        RECT 30.960 36.060 31.060 36.230 ;
        RECT 29.450 35.780 31.060 36.060 ;
      LAYER li1 ;
        RECT 26.530 34.880 27.040 35.090 ;
      LAYER li1 ;
        RECT 27.240 35.000 29.110 35.170 ;
        RECT 29.760 35.380 31.060 35.780 ;
      LAYER li1 ;
        RECT 26.180 34.530 27.240 34.700 ;
        RECT 26.970 34.450 27.240 34.530 ;
        RECT 27.690 34.510 28.200 34.820 ;
        RECT 28.450 34.510 29.160 34.820 ;
      LAYER li1 ;
        RECT 29.760 34.600 30.090 35.380 ;
        RECT 22.780 32.950 22.810 33.120 ;
        RECT 22.980 32.950 23.170 33.120 ;
        RECT 23.340 32.950 23.370 33.120 ;
        RECT 22.780 32.870 23.370 32.950 ;
        RECT 23.770 33.070 25.220 33.940 ;
        RECT 23.770 32.900 24.020 33.070 ;
        RECT 24.190 32.900 24.380 33.070 ;
        RECT 24.550 32.900 24.820 33.070 ;
        RECT 24.990 32.900 25.220 33.070 ;
        RECT 23.770 32.870 25.220 32.900 ;
        RECT 25.530 33.120 26.790 34.350 ;
      LAYER li1 ;
        RECT 26.970 33.370 27.490 34.450 ;
      LAYER li1 ;
        RECT 25.530 32.950 25.540 33.120 ;
        RECT 25.710 32.950 25.900 33.120 ;
        RECT 26.070 32.950 26.260 33.120 ;
        RECT 26.430 32.950 26.620 33.120 ;
        RECT 25.530 32.870 26.790 32.950 ;
      LAYER li1 ;
        RECT 27.320 32.870 27.490 33.370 ;
      LAYER li1 ;
        RECT 27.750 33.120 29.060 34.330 ;
        RECT 30.300 33.940 30.630 34.930 ;
        RECT 27.750 32.950 27.780 33.120 ;
        RECT 27.950 32.950 28.140 33.120 ;
        RECT 28.310 32.950 28.500 33.120 ;
        RECT 28.670 32.950 28.860 33.120 ;
        RECT 29.030 32.950 29.060 33.120 ;
        RECT 27.750 32.870 29.060 32.950 ;
        RECT 29.530 33.070 30.980 33.940 ;
        RECT 29.530 32.900 29.780 33.070 ;
        RECT 29.950 32.900 30.140 33.070 ;
        RECT 30.310 32.900 30.580 33.070 ;
        RECT 30.750 32.900 30.980 33.070 ;
        RECT 29.530 32.870 30.980 32.900 ;
      LAYER li1 ;
        RECT 31.330 32.870 31.580 36.130 ;
      LAYER li1 ;
        RECT 31.930 36.060 32.120 36.230 ;
        RECT 32.290 36.060 32.480 36.230 ;
        RECT 32.950 36.190 34.880 36.360 ;
        RECT 31.760 35.380 32.650 36.060 ;
        RECT 32.950 35.760 33.280 36.190 ;
        RECT 33.730 35.750 34.060 36.010 ;
        RECT 33.460 35.580 34.060 35.750 ;
        RECT 34.550 35.600 34.880 36.190 ;
        RECT 35.090 36.230 36.390 36.260 ;
        RECT 35.090 36.060 35.120 36.230 ;
        RECT 35.290 36.060 35.480 36.230 ;
        RECT 35.650 36.060 35.840 36.230 ;
        RECT 36.010 36.060 36.200 36.230 ;
        RECT 36.370 36.060 36.390 36.230 ;
        RECT 35.090 35.580 36.390 36.060 ;
        RECT 37.060 36.240 39.790 36.270 ;
        RECT 37.060 36.070 37.230 36.240 ;
        RECT 37.400 36.070 37.670 36.240 ;
        RECT 37.840 36.070 38.080 36.240 ;
        RECT 38.250 36.070 38.510 36.240 ;
        RECT 38.680 36.070 38.950 36.240 ;
        RECT 39.120 36.070 39.360 36.240 ;
        RECT 39.530 36.070 39.790 36.240 ;
        RECT 32.830 35.410 33.630 35.580 ;
        RECT 32.830 35.200 33.000 35.410 ;
      LAYER li1 ;
        RECT 34.240 35.400 34.910 35.420 ;
        RECT 33.810 35.230 36.080 35.400 ;
      LAYER li1 ;
        RECT 37.060 35.270 39.790 36.070 ;
        RECT 40.890 36.230 41.840 36.260 ;
        RECT 40.890 36.060 40.920 36.230 ;
        RECT 41.090 36.060 41.280 36.230 ;
        RECT 41.450 36.060 41.640 36.230 ;
        RECT 41.810 36.060 41.840 36.230 ;
        RECT 42.450 36.230 43.400 36.260 ;
        RECT 40.890 35.300 41.840 36.060 ;
      LAYER li1 ;
        RECT 42.020 35.420 42.270 36.130 ;
      LAYER li1 ;
        RECT 42.450 36.060 42.480 36.230 ;
        RECT 42.650 36.060 42.840 36.230 ;
        RECT 43.010 36.060 43.200 36.230 ;
        RECT 43.370 36.060 43.400 36.230 ;
        RECT 44.010 36.230 44.960 36.260 ;
        RECT 42.450 35.600 43.400 36.060 ;
      LAYER li1 ;
        RECT 43.580 35.420 43.830 36.130 ;
      LAYER li1 ;
        RECT 31.790 35.030 33.000 35.200 ;
      LAYER li1 ;
        RECT 33.180 35.060 33.980 35.230 ;
      LAYER li1 ;
        RECT 31.790 34.330 32.120 35.030 ;
      LAYER li1 ;
        RECT 33.180 34.850 33.350 35.060 ;
        RECT 32.620 34.570 33.350 34.850 ;
        RECT 32.790 34.510 32.960 34.570 ;
        RECT 33.530 34.510 33.960 34.880 ;
        RECT 34.160 34.510 34.450 35.050 ;
        RECT 34.690 34.720 35.400 35.050 ;
        RECT 35.750 34.610 36.080 35.230 ;
      LAYER li1 ;
        RECT 37.220 34.600 37.550 35.270 ;
        RECT 34.630 34.330 34.880 34.450 ;
        RECT 31.790 34.160 34.880 34.330 ;
        RECT 31.760 33.120 34.450 33.980 ;
        RECT 31.930 32.950 32.120 33.120 ;
        RECT 32.290 32.950 32.480 33.120 ;
        RECT 32.650 32.950 32.840 33.120 ;
        RECT 33.010 32.950 33.200 33.120 ;
        RECT 33.370 32.950 33.560 33.120 ;
        RECT 33.730 32.950 33.920 33.120 ;
        RECT 34.090 32.950 34.280 33.120 ;
        RECT 31.760 32.870 34.450 32.950 ;
        RECT 34.630 32.870 34.880 34.160 ;
        RECT 35.060 33.120 36.370 34.430 ;
        RECT 37.950 33.950 38.280 34.930 ;
        RECT 38.500 34.600 38.830 35.270 ;
      LAYER li1 ;
        RECT 42.020 35.250 43.830 35.420 ;
      LAYER li1 ;
        RECT 44.010 36.060 44.040 36.230 ;
        RECT 44.210 36.060 44.400 36.230 ;
        RECT 44.570 36.060 44.760 36.230 ;
        RECT 44.930 36.060 44.960 36.230 ;
        RECT 45.770 36.230 47.380 36.260 ;
        RECT 44.010 35.380 44.960 36.060 ;
      LAYER li1 ;
        RECT 42.020 35.080 42.190 35.250 ;
      LAYER li1 ;
        RECT 45.140 35.200 45.470 36.130 ;
        RECT 45.770 36.060 45.820 36.230 ;
        RECT 45.990 36.060 46.260 36.230 ;
        RECT 46.430 36.060 46.700 36.230 ;
        RECT 46.870 36.060 47.110 36.230 ;
        RECT 47.280 36.060 47.380 36.230 ;
        RECT 45.770 35.780 47.380 36.060 ;
        RECT 39.230 33.950 39.560 34.930 ;
      LAYER li1 ;
        RECT 40.930 34.850 42.190 35.080 ;
      LAYER li1 ;
        RECT 44.230 35.070 45.470 35.200 ;
        RECT 42.370 35.030 45.470 35.070 ;
        RECT 42.370 34.900 44.400 35.030 ;
      LAYER li1 ;
        RECT 42.020 34.720 42.190 34.850 ;
        RECT 42.020 34.550 43.910 34.720 ;
      LAYER li1 ;
        RECT 35.060 32.950 35.090 33.120 ;
        RECT 35.260 32.950 35.450 33.120 ;
        RECT 35.620 32.950 35.810 33.120 ;
        RECT 35.980 32.950 36.170 33.120 ;
        RECT 36.340 32.950 36.370 33.120 ;
        RECT 35.060 32.890 36.370 32.950 ;
        RECT 36.980 33.070 39.720 33.950 ;
        RECT 36.980 32.900 37.190 33.070 ;
        RECT 37.360 32.900 37.630 33.070 ;
        RECT 37.800 32.900 38.040 33.070 ;
        RECT 38.210 32.900 38.470 33.070 ;
        RECT 38.640 32.900 38.910 33.070 ;
        RECT 39.080 32.900 39.320 33.070 ;
        RECT 39.490 32.900 39.720 33.070 ;
        RECT 36.980 32.880 39.720 32.900 ;
        RECT 40.890 33.120 41.840 34.450 ;
        RECT 40.890 32.950 40.920 33.120 ;
        RECT 41.090 32.950 41.280 33.120 ;
        RECT 41.450 32.950 41.640 33.120 ;
        RECT 41.810 32.950 41.840 33.120 ;
        RECT 40.890 32.870 41.840 32.950 ;
      LAYER li1 ;
        RECT 42.020 32.870 42.270 34.550 ;
      LAYER li1 ;
        RECT 42.450 33.120 43.400 34.370 ;
        RECT 42.450 32.950 42.480 33.120 ;
        RECT 42.650 32.950 42.840 33.120 ;
        RECT 43.010 32.950 43.200 33.120 ;
        RECT 43.370 32.950 43.400 33.120 ;
        RECT 42.450 32.870 43.400 32.950 ;
      LAYER li1 ;
        RECT 43.580 32.870 43.910 34.550 ;
        RECT 44.690 34.510 45.020 34.850 ;
      LAYER li1 ;
        RECT 44.090 33.120 45.040 34.330 ;
        RECT 44.090 32.950 44.120 33.120 ;
        RECT 44.290 32.950 44.480 33.120 ;
        RECT 44.650 32.950 44.840 33.120 ;
        RECT 45.010 32.950 45.040 33.120 ;
        RECT 44.090 32.870 45.040 32.950 ;
        RECT 45.220 32.870 45.470 35.030 ;
        RECT 46.080 35.380 47.380 35.780 ;
        RECT 47.610 36.230 48.560 36.260 ;
        RECT 47.610 36.060 47.640 36.230 ;
        RECT 47.810 36.060 48.000 36.230 ;
        RECT 48.170 36.060 48.360 36.230 ;
        RECT 48.530 36.060 48.560 36.230 ;
        RECT 49.170 36.230 50.120 36.260 ;
        RECT 46.080 34.600 46.410 35.380 ;
        RECT 47.610 35.300 48.560 36.060 ;
      LAYER li1 ;
        RECT 48.740 35.420 48.990 36.130 ;
      LAYER li1 ;
        RECT 49.170 36.060 49.200 36.230 ;
        RECT 49.370 36.060 49.560 36.230 ;
        RECT 49.730 36.060 49.920 36.230 ;
        RECT 50.090 36.060 50.120 36.230 ;
        RECT 50.730 36.230 51.680 36.260 ;
        RECT 49.170 35.600 50.120 36.060 ;
      LAYER li1 ;
        RECT 50.300 35.420 50.550 36.130 ;
        RECT 48.740 35.250 50.550 35.420 ;
      LAYER li1 ;
        RECT 50.730 36.060 50.760 36.230 ;
        RECT 50.930 36.060 51.120 36.230 ;
        RECT 51.290 36.060 51.480 36.230 ;
        RECT 51.650 36.060 51.680 36.230 ;
        RECT 52.490 36.230 54.100 36.260 ;
        RECT 50.730 35.380 51.680 36.060 ;
      LAYER li1 ;
        RECT 48.740 35.080 48.910 35.250 ;
      LAYER li1 ;
        RECT 51.860 35.200 52.190 36.130 ;
        RECT 52.490 36.060 52.540 36.230 ;
        RECT 52.710 36.060 52.980 36.230 ;
        RECT 53.150 36.060 53.420 36.230 ;
        RECT 53.590 36.060 53.830 36.230 ;
        RECT 54.000 36.060 54.100 36.230 ;
        RECT 52.490 35.780 54.100 36.060 ;
        RECT 46.620 33.940 46.950 34.930 ;
      LAYER li1 ;
        RECT 47.650 34.850 48.910 35.080 ;
      LAYER li1 ;
        RECT 50.950 35.070 52.190 35.200 ;
        RECT 49.090 35.030 52.190 35.070 ;
        RECT 49.090 34.900 51.120 35.030 ;
      LAYER li1 ;
        RECT 48.740 34.720 48.910 34.850 ;
        RECT 48.740 34.550 50.630 34.720 ;
      LAYER li1 ;
        RECT 45.850 33.070 47.300 33.940 ;
        RECT 45.850 32.900 46.100 33.070 ;
        RECT 46.270 32.900 46.460 33.070 ;
        RECT 46.630 32.900 46.900 33.070 ;
        RECT 47.070 32.900 47.300 33.070 ;
        RECT 45.850 32.870 47.300 32.900 ;
        RECT 47.610 33.120 48.560 34.450 ;
        RECT 47.610 32.950 47.640 33.120 ;
        RECT 47.810 32.950 48.000 33.120 ;
        RECT 48.170 32.950 48.360 33.120 ;
        RECT 48.530 32.950 48.560 33.120 ;
        RECT 47.610 32.870 48.560 32.950 ;
      LAYER li1 ;
        RECT 48.740 32.870 48.990 34.550 ;
      LAYER li1 ;
        RECT 49.170 33.120 50.120 34.370 ;
        RECT 49.170 32.950 49.200 33.120 ;
        RECT 49.370 32.950 49.560 33.120 ;
        RECT 49.730 32.950 49.920 33.120 ;
        RECT 50.090 32.950 50.120 33.120 ;
        RECT 49.170 32.870 50.120 32.950 ;
      LAYER li1 ;
        RECT 50.300 32.870 50.630 34.550 ;
        RECT 51.410 34.510 51.740 34.850 ;
      LAYER li1 ;
        RECT 50.810 33.120 51.760 34.330 ;
        RECT 50.810 32.950 50.840 33.120 ;
        RECT 51.010 32.950 51.200 33.120 ;
        RECT 51.370 32.950 51.560 33.120 ;
        RECT 51.730 32.950 51.760 33.120 ;
        RECT 50.810 32.870 51.760 32.950 ;
        RECT 51.940 32.870 52.190 35.030 ;
        RECT 52.800 35.380 54.100 35.780 ;
        RECT 54.330 36.230 55.280 36.260 ;
        RECT 54.330 36.060 54.360 36.230 ;
        RECT 54.530 36.060 54.720 36.230 ;
        RECT 54.890 36.060 55.080 36.230 ;
        RECT 55.250 36.060 55.280 36.230 ;
        RECT 55.890 36.230 56.840 36.260 ;
        RECT 52.800 34.600 53.130 35.380 ;
        RECT 54.330 35.300 55.280 36.060 ;
      LAYER li1 ;
        RECT 55.460 35.420 55.710 36.130 ;
      LAYER li1 ;
        RECT 55.890 36.060 55.920 36.230 ;
        RECT 56.090 36.060 56.280 36.230 ;
        RECT 56.450 36.060 56.640 36.230 ;
        RECT 56.810 36.060 56.840 36.230 ;
        RECT 57.450 36.230 58.400 36.260 ;
        RECT 55.890 35.600 56.840 36.060 ;
      LAYER li1 ;
        RECT 57.020 35.420 57.270 36.130 ;
        RECT 55.460 35.250 57.270 35.420 ;
      LAYER li1 ;
        RECT 57.450 36.060 57.480 36.230 ;
        RECT 57.650 36.060 57.840 36.230 ;
        RECT 58.010 36.060 58.200 36.230 ;
        RECT 58.370 36.060 58.400 36.230 ;
        RECT 59.210 36.230 60.820 36.260 ;
        RECT 57.450 35.380 58.400 36.060 ;
      LAYER li1 ;
        RECT 55.460 35.080 55.630 35.250 ;
      LAYER li1 ;
        RECT 58.580 35.200 58.910 36.130 ;
        RECT 59.210 36.060 59.260 36.230 ;
        RECT 59.430 36.060 59.700 36.230 ;
        RECT 59.870 36.060 60.140 36.230 ;
        RECT 60.310 36.060 60.550 36.230 ;
        RECT 60.720 36.060 60.820 36.230 ;
        RECT 61.520 36.230 62.470 36.260 ;
        RECT 59.210 35.780 60.820 36.060 ;
        RECT 53.340 33.940 53.670 34.930 ;
      LAYER li1 ;
        RECT 54.370 34.850 55.630 35.080 ;
      LAYER li1 ;
        RECT 57.670 35.070 58.910 35.200 ;
        RECT 55.810 35.030 58.910 35.070 ;
        RECT 55.810 34.900 57.840 35.030 ;
      LAYER li1 ;
        RECT 55.460 34.720 55.630 34.850 ;
        RECT 55.460 34.550 57.350 34.720 ;
      LAYER li1 ;
        RECT 52.570 33.070 54.020 33.940 ;
        RECT 52.570 32.900 52.820 33.070 ;
        RECT 52.990 32.900 53.180 33.070 ;
        RECT 53.350 32.900 53.620 33.070 ;
        RECT 53.790 32.900 54.020 33.070 ;
        RECT 52.570 32.870 54.020 32.900 ;
        RECT 54.330 33.120 55.280 34.450 ;
        RECT 54.330 32.950 54.360 33.120 ;
        RECT 54.530 32.950 54.720 33.120 ;
        RECT 54.890 32.950 55.080 33.120 ;
        RECT 55.250 32.950 55.280 33.120 ;
        RECT 54.330 32.870 55.280 32.950 ;
      LAYER li1 ;
        RECT 55.460 32.870 55.710 34.550 ;
      LAYER li1 ;
        RECT 55.890 33.120 56.840 34.370 ;
        RECT 55.890 32.950 55.920 33.120 ;
        RECT 56.090 32.950 56.280 33.120 ;
        RECT 56.450 32.950 56.640 33.120 ;
        RECT 56.810 32.950 56.840 33.120 ;
        RECT 55.890 32.870 56.840 32.950 ;
      LAYER li1 ;
        RECT 57.020 32.870 57.350 34.550 ;
        RECT 58.130 34.510 58.460 34.850 ;
      LAYER li1 ;
        RECT 57.530 33.120 58.480 34.330 ;
        RECT 57.530 32.950 57.560 33.120 ;
        RECT 57.730 32.950 57.920 33.120 ;
        RECT 58.090 32.950 58.280 33.120 ;
        RECT 58.450 32.950 58.480 33.120 ;
        RECT 57.530 32.870 58.480 32.950 ;
        RECT 58.660 32.870 58.910 35.030 ;
        RECT 59.520 35.380 60.820 35.780 ;
        RECT 59.520 34.600 59.850 35.380 ;
        RECT 60.060 33.940 60.390 34.930 ;
        RECT 61.070 34.270 61.340 36.130 ;
        RECT 61.520 36.060 61.550 36.230 ;
        RECT 61.720 36.060 61.910 36.230 ;
        RECT 62.080 36.060 62.270 36.230 ;
        RECT 62.440 36.060 62.470 36.230 ;
        RECT 63.160 36.230 63.750 36.260 ;
        RECT 61.520 35.630 62.470 36.060 ;
        RECT 62.650 35.630 62.980 36.130 ;
        RECT 62.200 34.270 62.530 34.770 ;
        RECT 61.070 34.100 62.530 34.270 ;
        RECT 59.290 33.070 60.740 33.940 ;
        RECT 61.070 33.170 61.400 34.100 ;
        RECT 59.290 32.900 59.540 33.070 ;
        RECT 59.710 32.900 59.900 33.070 ;
        RECT 60.070 32.900 60.340 33.070 ;
        RECT 60.510 32.900 60.740 33.070 ;
        RECT 61.590 33.120 62.180 33.900 ;
        RECT 61.590 32.950 61.620 33.120 ;
        RECT 61.790 32.950 61.980 33.120 ;
        RECT 62.150 32.950 62.180 33.120 ;
        RECT 61.590 32.920 62.180 32.950 ;
        RECT 62.360 32.990 62.530 34.100 ;
        RECT 62.710 34.710 62.980 35.630 ;
        RECT 63.160 36.060 63.190 36.230 ;
        RECT 63.360 36.060 63.550 36.230 ;
        RECT 63.720 36.060 63.750 36.230 ;
        RECT 68.120 36.230 69.070 36.260 ;
        RECT 63.160 35.380 63.750 36.060 ;
      LAYER li1 ;
        RECT 64.030 36.000 66.970 36.170 ;
        RECT 64.030 35.010 64.200 36.000 ;
      LAYER li1 ;
        RECT 62.710 34.480 63.240 34.710 ;
        RECT 62.710 33.170 62.960 34.480 ;
      LAYER li1 ;
        RECT 63.660 34.140 64.200 35.010 ;
        RECT 64.380 34.520 64.710 35.820 ;
      LAYER li1 ;
        RECT 64.890 35.300 65.160 35.800 ;
        RECT 65.610 35.550 65.940 35.800 ;
        RECT 65.610 35.380 66.620 35.550 ;
        RECT 64.890 34.310 65.060 35.300 ;
        RECT 65.940 34.710 66.270 35.200 ;
        RECT 64.840 34.140 65.060 34.310 ;
        RECT 65.240 34.480 66.270 34.710 ;
        RECT 66.450 35.150 66.620 35.380 ;
      LAYER li1 ;
        RECT 66.800 35.500 66.970 36.000 ;
      LAYER li1 ;
        RECT 68.120 36.060 68.150 36.230 ;
        RECT 68.320 36.060 68.510 36.230 ;
        RECT 68.680 36.060 68.870 36.230 ;
        RECT 69.040 36.060 69.070 36.230 ;
        RECT 68.120 35.680 69.070 36.060 ;
      LAYER li1 ;
        RECT 69.250 36.190 71.910 36.360 ;
        RECT 69.250 35.500 69.420 36.190 ;
        RECT 66.800 35.330 69.420 35.500 ;
      LAYER li1 ;
        RECT 66.450 34.980 69.070 35.150 ;
        RECT 64.840 33.960 65.010 34.140 ;
        RECT 65.240 33.960 65.410 34.480 ;
        RECT 66.450 34.300 66.620 34.980 ;
      LAYER li1 ;
        RECT 69.250 34.800 69.420 35.330 ;
      LAYER li1 ;
        RECT 63.200 33.790 65.010 33.960 ;
        RECT 63.200 33.170 63.450 33.790 ;
        RECT 63.630 33.440 64.660 33.610 ;
        RECT 63.630 32.990 63.800 33.440 ;
        RECT 59.290 32.870 60.740 32.900 ;
        RECT 62.360 32.820 63.800 32.990 ;
        RECT 63.980 33.120 64.310 33.260 ;
        RECT 63.980 32.950 64.010 33.120 ;
        RECT 64.180 32.950 64.310 33.120 ;
        RECT 63.980 32.920 64.310 32.950 ;
        RECT 64.490 32.990 64.660 33.440 ;
        RECT 64.840 33.170 65.010 33.790 ;
        RECT 65.190 33.630 65.410 33.960 ;
        RECT 65.590 34.130 66.620 34.300 ;
        RECT 66.800 34.450 67.130 34.800 ;
      LAYER li1 ;
        RECT 67.570 34.630 69.420 34.800 ;
      LAYER li1 ;
        RECT 69.600 35.300 69.930 36.010 ;
        RECT 70.390 35.840 71.560 36.010 ;
        RECT 70.390 35.300 70.720 35.840 ;
        RECT 69.600 34.450 69.860 35.300 ;
        RECT 70.930 35.040 71.210 35.540 ;
        RECT 66.800 34.280 69.860 34.450 ;
        RECT 65.590 33.430 65.760 34.130 ;
        RECT 66.450 34.100 66.620 34.130 ;
        RECT 65.940 33.750 66.270 33.950 ;
        RECT 66.450 33.930 68.220 34.100 ;
        RECT 65.940 33.630 67.710 33.750 ;
        RECT 66.060 33.580 67.710 33.630 ;
        RECT 65.540 33.170 65.870 33.430 ;
        RECT 66.060 32.990 66.230 33.580 ;
        RECT 64.490 32.820 66.230 32.990 ;
        RECT 66.410 33.120 67.360 33.400 ;
        RECT 66.410 32.950 66.440 33.120 ;
        RECT 66.610 32.950 66.800 33.120 ;
        RECT 66.970 32.950 67.160 33.120 ;
        RECT 67.330 32.950 67.360 33.120 ;
        RECT 66.410 32.920 67.360 32.950 ;
        RECT 67.540 32.990 67.710 33.580 ;
        RECT 67.890 33.170 68.220 33.930 ;
        RECT 69.530 33.700 69.860 34.280 ;
        RECT 70.040 34.870 71.210 35.040 ;
        RECT 70.040 33.520 70.210 34.870 ;
        RECT 70.590 34.190 70.920 34.690 ;
        RECT 71.390 34.440 71.560 35.840 ;
      LAYER li1 ;
        RECT 71.740 35.530 71.910 36.190 ;
      LAYER li1 ;
        RECT 72.090 36.230 73.040 36.260 ;
        RECT 72.090 36.060 72.120 36.230 ;
        RECT 72.290 36.060 72.480 36.230 ;
        RECT 72.650 36.060 72.840 36.230 ;
        RECT 73.010 36.060 73.040 36.230 ;
        RECT 74.700 36.230 75.650 36.260 ;
        RECT 72.090 35.710 73.040 36.060 ;
        RECT 73.580 35.630 73.910 36.130 ;
        RECT 74.700 36.060 74.730 36.230 ;
        RECT 74.900 36.060 75.090 36.230 ;
        RECT 75.260 36.060 75.450 36.230 ;
        RECT 75.620 36.060 75.650 36.230 ;
      LAYER li1 ;
        RECT 71.740 35.360 72.750 35.530 ;
      LAYER li1 ;
        RECT 71.770 34.790 72.100 35.180 ;
      LAYER li1 ;
        RECT 72.420 34.970 72.750 35.360 ;
      LAYER li1 ;
        RECT 73.580 34.790 73.810 35.630 ;
        RECT 74.190 35.130 74.520 35.630 ;
        RECT 74.700 35.130 75.650 36.060 ;
        RECT 76.490 36.230 78.100 36.260 ;
        RECT 76.490 36.060 76.540 36.230 ;
        RECT 76.710 36.060 76.980 36.230 ;
        RECT 77.150 36.060 77.420 36.230 ;
        RECT 77.590 36.060 77.830 36.230 ;
        RECT 78.000 36.060 78.100 36.230 ;
        RECT 71.770 34.620 73.810 34.790 ;
        RECT 71.100 34.270 73.460 34.440 ;
        RECT 71.100 33.950 71.270 34.270 ;
        RECT 73.640 34.090 73.810 34.620 ;
        RECT 68.400 33.350 70.210 33.520 ;
        RECT 70.390 33.780 71.270 33.950 ;
        RECT 68.400 32.990 68.570 33.350 ;
        RECT 67.540 32.820 68.570 32.990 ;
        RECT 68.750 33.120 69.700 33.170 ;
        RECT 68.750 32.950 68.780 33.120 ;
        RECT 68.950 32.950 69.140 33.120 ;
        RECT 69.310 32.950 69.500 33.120 ;
        RECT 69.670 32.950 69.700 33.120 ;
        RECT 68.750 32.870 69.700 32.950 ;
        RECT 70.390 32.870 70.640 33.780 ;
        RECT 71.450 33.120 72.400 33.950 ;
        RECT 72.800 33.920 73.810 34.090 ;
        RECT 74.310 34.950 74.520 35.130 ;
        RECT 74.310 34.620 75.680 34.950 ;
        RECT 72.800 33.450 73.050 33.920 ;
        RECT 73.230 33.120 74.130 33.740 ;
        RECT 74.310 33.620 74.560 34.620 ;
        RECT 71.450 32.950 71.480 33.120 ;
        RECT 71.650 32.950 71.840 33.120 ;
        RECT 72.010 32.950 72.200 33.120 ;
        RECT 72.370 32.950 72.400 33.120 ;
        RECT 73.400 32.950 73.590 33.120 ;
        RECT 73.760 32.950 73.950 33.120 ;
        RECT 74.120 32.950 74.130 33.120 ;
        RECT 71.450 32.920 72.400 32.950 ;
        RECT 73.230 32.920 74.130 32.950 ;
        RECT 74.740 33.120 75.680 34.430 ;
        RECT 74.740 32.950 74.760 33.120 ;
        RECT 74.930 32.950 75.120 33.120 ;
        RECT 75.290 32.950 75.480 33.120 ;
        RECT 75.650 32.950 75.680 33.120 ;
        RECT 74.740 32.890 75.680 32.950 ;
      LAYER li1 ;
        RECT 75.860 32.890 76.200 35.960 ;
      LAYER li1 ;
        RECT 76.490 35.780 78.100 36.060 ;
        RECT 76.800 35.380 78.100 35.780 ;
        RECT 78.330 36.230 78.920 36.260 ;
        RECT 78.330 36.060 78.360 36.230 ;
        RECT 78.530 36.060 78.720 36.230 ;
        RECT 78.890 36.060 78.920 36.230 ;
        RECT 79.850 36.230 81.460 36.260 ;
        RECT 76.800 34.600 77.130 35.380 ;
        RECT 78.330 35.300 78.920 36.060 ;
        RECT 77.340 33.940 77.670 34.930 ;
      LAYER li1 ;
        RECT 78.370 34.690 79.080 35.080 ;
        RECT 79.260 34.450 79.590 36.130 ;
      LAYER li1 ;
        RECT 79.850 36.060 79.900 36.230 ;
        RECT 80.070 36.060 80.340 36.230 ;
        RECT 80.510 36.060 80.780 36.230 ;
        RECT 80.950 36.060 81.190 36.230 ;
        RECT 81.360 36.060 81.460 36.230 ;
        RECT 79.850 35.780 81.460 36.060 ;
        RECT 80.160 35.380 81.460 35.780 ;
        RECT 81.690 36.230 82.640 36.260 ;
        RECT 81.690 36.060 81.720 36.230 ;
        RECT 81.890 36.060 82.080 36.230 ;
        RECT 82.250 36.060 82.440 36.230 ;
        RECT 82.610 36.060 82.640 36.230 ;
        RECT 83.250 36.230 84.200 36.260 ;
        RECT 80.160 34.600 80.490 35.380 ;
        RECT 81.690 35.300 82.640 36.060 ;
      LAYER li1 ;
        RECT 82.820 35.420 83.070 36.130 ;
      LAYER li1 ;
        RECT 83.250 36.060 83.280 36.230 ;
        RECT 83.450 36.060 83.640 36.230 ;
        RECT 83.810 36.060 84.000 36.230 ;
        RECT 84.170 36.060 84.200 36.230 ;
        RECT 84.810 36.230 85.760 36.260 ;
        RECT 83.250 35.600 84.200 36.060 ;
      LAYER li1 ;
        RECT 84.380 35.420 84.630 36.130 ;
        RECT 82.820 35.250 84.630 35.420 ;
      LAYER li1 ;
        RECT 84.810 36.060 84.840 36.230 ;
        RECT 85.010 36.060 85.200 36.230 ;
        RECT 85.370 36.060 85.560 36.230 ;
        RECT 85.730 36.060 85.760 36.230 ;
        RECT 86.570 36.230 88.180 36.260 ;
        RECT 84.810 35.380 85.760 36.060 ;
      LAYER li1 ;
        RECT 82.820 35.080 82.990 35.250 ;
      LAYER li1 ;
        RECT 85.940 35.200 86.270 36.130 ;
        RECT 86.570 36.060 86.620 36.230 ;
        RECT 86.790 36.060 87.060 36.230 ;
        RECT 87.230 36.060 87.500 36.230 ;
        RECT 87.670 36.060 87.910 36.230 ;
        RECT 88.080 36.060 88.180 36.230 ;
        RECT 86.570 35.780 88.180 36.060 ;
        RECT 76.570 33.070 78.020 33.940 ;
        RECT 76.570 32.900 76.820 33.070 ;
        RECT 76.990 32.900 77.180 33.070 ;
        RECT 77.350 32.900 77.620 33.070 ;
        RECT 77.790 32.900 78.020 33.070 ;
        RECT 76.570 32.870 78.020 32.900 ;
        RECT 78.330 33.120 78.920 34.450 ;
        RECT 78.330 32.950 78.360 33.120 ;
        RECT 78.530 32.950 78.720 33.120 ;
        RECT 78.890 32.950 78.920 33.120 ;
        RECT 78.330 32.870 78.920 32.950 ;
      LAYER li1 ;
        RECT 79.200 32.870 79.590 34.450 ;
      LAYER li1 ;
        RECT 80.700 33.940 81.030 34.930 ;
      LAYER li1 ;
        RECT 81.730 34.850 82.990 35.080 ;
      LAYER li1 ;
        RECT 85.030 35.070 86.270 35.200 ;
        RECT 83.170 35.030 86.270 35.070 ;
        RECT 83.170 34.900 85.200 35.030 ;
      LAYER li1 ;
        RECT 82.820 34.720 82.990 34.850 ;
        RECT 82.820 34.550 84.710 34.720 ;
      LAYER li1 ;
        RECT 79.930 33.070 81.380 33.940 ;
        RECT 79.930 32.900 80.180 33.070 ;
        RECT 80.350 32.900 80.540 33.070 ;
        RECT 80.710 32.900 80.980 33.070 ;
        RECT 81.150 32.900 81.380 33.070 ;
        RECT 79.930 32.870 81.380 32.900 ;
        RECT 81.690 33.120 82.640 34.450 ;
        RECT 81.690 32.950 81.720 33.120 ;
        RECT 81.890 32.950 82.080 33.120 ;
        RECT 82.250 32.950 82.440 33.120 ;
        RECT 82.610 32.950 82.640 33.120 ;
        RECT 81.690 32.870 82.640 32.950 ;
      LAYER li1 ;
        RECT 82.820 32.870 83.070 34.550 ;
      LAYER li1 ;
        RECT 83.250 33.120 84.200 34.370 ;
        RECT 83.250 32.950 83.280 33.120 ;
        RECT 83.450 32.950 83.640 33.120 ;
        RECT 83.810 32.950 84.000 33.120 ;
        RECT 84.170 32.950 84.200 33.120 ;
        RECT 83.250 32.870 84.200 32.950 ;
      LAYER li1 ;
        RECT 84.380 32.870 84.710 34.550 ;
        RECT 85.490 34.510 85.820 34.850 ;
      LAYER li1 ;
        RECT 84.890 33.120 85.840 34.330 ;
        RECT 84.890 32.950 84.920 33.120 ;
        RECT 85.090 32.950 85.280 33.120 ;
        RECT 85.450 32.950 85.640 33.120 ;
        RECT 85.810 32.950 85.840 33.120 ;
        RECT 84.890 32.870 85.840 32.950 ;
        RECT 86.020 32.870 86.270 35.030 ;
        RECT 86.880 35.380 88.180 35.780 ;
        RECT 89.370 36.230 90.320 36.260 ;
        RECT 89.370 36.060 89.400 36.230 ;
        RECT 89.570 36.060 89.760 36.230 ;
        RECT 89.930 36.060 90.120 36.230 ;
        RECT 90.290 36.060 90.320 36.230 ;
        RECT 90.930 36.230 91.880 36.260 ;
        RECT 86.880 34.600 87.210 35.380 ;
        RECT 89.370 35.300 90.320 36.060 ;
      LAYER li1 ;
        RECT 90.500 35.420 90.750 36.130 ;
      LAYER li1 ;
        RECT 90.930 36.060 90.960 36.230 ;
        RECT 91.130 36.060 91.320 36.230 ;
        RECT 91.490 36.060 91.680 36.230 ;
        RECT 91.850 36.060 91.880 36.230 ;
        RECT 92.490 36.230 93.440 36.260 ;
        RECT 90.930 35.600 91.880 36.060 ;
      LAYER li1 ;
        RECT 92.060 35.420 92.310 36.130 ;
        RECT 90.500 35.250 92.310 35.420 ;
      LAYER li1 ;
        RECT 92.490 36.060 92.520 36.230 ;
        RECT 92.690 36.060 92.880 36.230 ;
        RECT 93.050 36.060 93.240 36.230 ;
        RECT 93.410 36.060 93.440 36.230 ;
        RECT 94.250 36.230 95.860 36.260 ;
        RECT 92.490 35.380 93.440 36.060 ;
      LAYER li1 ;
        RECT 90.500 35.080 90.670 35.250 ;
      LAYER li1 ;
        RECT 93.620 35.200 93.950 36.130 ;
        RECT 94.250 36.060 94.300 36.230 ;
        RECT 94.470 36.060 94.740 36.230 ;
        RECT 94.910 36.060 95.180 36.230 ;
        RECT 95.350 36.060 95.590 36.230 ;
        RECT 95.760 36.060 95.860 36.230 ;
        RECT 94.250 35.780 95.860 36.060 ;
        RECT 87.420 33.940 87.750 34.930 ;
      LAYER li1 ;
        RECT 89.410 34.850 90.670 35.080 ;
      LAYER li1 ;
        RECT 92.710 35.070 93.950 35.200 ;
        RECT 90.850 35.030 93.950 35.070 ;
        RECT 90.850 34.900 92.880 35.030 ;
      LAYER li1 ;
        RECT 90.500 34.720 90.670 34.850 ;
        RECT 90.500 34.550 92.390 34.720 ;
      LAYER li1 ;
        RECT 86.650 33.070 88.100 33.940 ;
        RECT 86.650 32.900 86.900 33.070 ;
        RECT 87.070 32.900 87.260 33.070 ;
        RECT 87.430 32.900 87.700 33.070 ;
        RECT 87.870 32.900 88.100 33.070 ;
        RECT 86.650 32.870 88.100 32.900 ;
        RECT 89.370 33.120 90.320 34.450 ;
        RECT 89.370 32.950 89.400 33.120 ;
        RECT 89.570 32.950 89.760 33.120 ;
        RECT 89.930 32.950 90.120 33.120 ;
        RECT 90.290 32.950 90.320 33.120 ;
        RECT 89.370 32.870 90.320 32.950 ;
      LAYER li1 ;
        RECT 90.500 32.870 90.750 34.550 ;
      LAYER li1 ;
        RECT 90.930 33.120 91.880 34.370 ;
        RECT 90.930 32.950 90.960 33.120 ;
        RECT 91.130 32.950 91.320 33.120 ;
        RECT 91.490 32.950 91.680 33.120 ;
        RECT 91.850 32.950 91.880 33.120 ;
        RECT 90.930 32.870 91.880 32.950 ;
      LAYER li1 ;
        RECT 92.060 32.870 92.390 34.550 ;
        RECT 93.170 34.510 93.500 34.850 ;
      LAYER li1 ;
        RECT 92.570 33.120 93.520 34.330 ;
        RECT 92.570 32.950 92.600 33.120 ;
        RECT 92.770 32.950 92.960 33.120 ;
        RECT 93.130 32.950 93.320 33.120 ;
        RECT 93.490 32.950 93.520 33.120 ;
        RECT 92.570 32.870 93.520 32.950 ;
        RECT 93.700 32.870 93.950 35.030 ;
        RECT 94.560 35.380 95.860 35.780 ;
        RECT 96.160 36.190 97.970 36.360 ;
        RECT 94.560 34.600 94.890 35.380 ;
        RECT 96.160 35.270 96.490 36.190 ;
      LAYER li1 ;
        RECT 96.740 35.790 97.270 36.010 ;
        RECT 96.740 35.620 97.280 35.790 ;
        RECT 96.740 35.270 97.270 35.620 ;
      LAYER li1 ;
        RECT 95.100 33.940 95.430 34.930 ;
      LAYER li1 ;
        RECT 96.130 34.760 96.550 35.090 ;
        RECT 96.740 34.700 96.910 35.270 ;
      LAYER li1 ;
        RECT 97.800 35.170 97.970 36.190 ;
        RECT 98.150 36.230 99.250 36.260 ;
        RECT 98.150 36.060 98.200 36.230 ;
        RECT 98.370 36.060 98.560 36.230 ;
        RECT 98.730 36.060 98.920 36.230 ;
        RECT 99.090 36.060 99.250 36.230 ;
        RECT 100.420 36.240 103.150 36.270 ;
        RECT 98.150 35.350 99.250 36.060 ;
        RECT 99.420 35.170 99.670 36.100 ;
        RECT 100.420 36.070 100.590 36.240 ;
        RECT 100.760 36.070 101.030 36.240 ;
        RECT 101.200 36.070 101.440 36.240 ;
        RECT 101.610 36.070 101.870 36.240 ;
        RECT 102.040 36.070 102.310 36.240 ;
        RECT 102.480 36.070 102.720 36.240 ;
        RECT 102.890 36.070 103.150 36.240 ;
        RECT 100.420 35.270 103.150 36.070 ;
        RECT 104.730 36.230 105.640 36.260 ;
        RECT 104.730 36.060 104.740 36.230 ;
        RECT 104.910 36.060 105.100 36.230 ;
        RECT 105.270 36.060 105.460 36.230 ;
        RECT 105.630 36.060 105.640 36.230 ;
        RECT 106.680 36.230 107.270 36.260 ;
        RECT 104.730 35.630 105.640 36.060 ;
        RECT 105.820 35.630 106.150 36.130 ;
        RECT 106.680 36.060 106.710 36.230 ;
        RECT 106.880 36.060 107.070 36.230 ;
        RECT 107.240 36.060 107.270 36.230 ;
        RECT 108.170 36.230 109.780 36.260 ;
      LAYER li1 ;
        RECT 97.090 34.880 97.600 35.090 ;
      LAYER li1 ;
        RECT 97.800 35.000 99.670 35.170 ;
      LAYER li1 ;
        RECT 96.740 34.530 97.800 34.700 ;
        RECT 97.530 34.450 97.800 34.530 ;
        RECT 98.250 34.510 98.760 34.820 ;
        RECT 99.010 34.510 99.720 34.820 ;
      LAYER li1 ;
        RECT 100.580 34.600 100.910 35.270 ;
        RECT 94.330 33.070 95.780 33.940 ;
        RECT 94.330 32.900 94.580 33.070 ;
        RECT 94.750 32.900 94.940 33.070 ;
        RECT 95.110 32.900 95.380 33.070 ;
        RECT 95.550 32.900 95.780 33.070 ;
        RECT 94.330 32.870 95.780 32.900 ;
        RECT 96.090 33.120 97.350 34.350 ;
      LAYER li1 ;
        RECT 97.530 33.370 98.050 34.450 ;
      LAYER li1 ;
        RECT 96.090 32.950 96.100 33.120 ;
        RECT 96.270 32.950 96.460 33.120 ;
        RECT 96.630 32.950 96.820 33.120 ;
        RECT 96.990 32.950 97.180 33.120 ;
        RECT 96.090 32.870 97.350 32.950 ;
      LAYER li1 ;
        RECT 97.880 32.870 98.050 33.370 ;
      LAYER li1 ;
        RECT 98.310 33.120 99.620 34.330 ;
        RECT 101.310 33.950 101.640 34.930 ;
        RECT 101.860 34.600 102.190 35.270 ;
        RECT 102.590 33.950 102.920 34.930 ;
      LAYER li1 ;
        RECT 105.250 34.900 105.580 35.450 ;
      LAYER li1 ;
        RECT 105.820 34.720 105.990 35.630 ;
      LAYER li1 ;
        RECT 106.170 34.900 106.500 35.450 ;
      LAYER li1 ;
        RECT 106.680 35.300 107.270 36.060 ;
        RECT 107.090 34.720 107.420 34.900 ;
        RECT 105.040 34.550 107.420 34.720 ;
        RECT 105.040 33.950 105.290 34.550 ;
        RECT 98.310 32.950 98.340 33.120 ;
        RECT 98.510 32.950 98.700 33.120 ;
        RECT 98.870 32.950 99.060 33.120 ;
        RECT 99.230 32.950 99.420 33.120 ;
        RECT 99.590 32.950 99.620 33.120 ;
        RECT 98.310 32.870 99.620 32.950 ;
        RECT 100.340 33.070 103.080 33.950 ;
        RECT 105.470 33.120 107.440 34.370 ;
        RECT 100.340 32.900 100.550 33.070 ;
        RECT 100.720 32.900 100.990 33.070 ;
        RECT 101.160 32.900 101.400 33.070 ;
        RECT 101.570 32.900 101.830 33.070 ;
        RECT 102.000 32.900 102.270 33.070 ;
        RECT 102.440 32.900 102.680 33.070 ;
        RECT 102.850 32.900 103.080 33.070 ;
        RECT 105.640 32.950 105.830 33.120 ;
        RECT 106.000 32.950 106.190 33.120 ;
        RECT 106.360 32.950 106.550 33.120 ;
        RECT 106.720 32.950 106.910 33.120 ;
        RECT 107.080 32.950 107.270 33.120 ;
        RECT 100.340 32.880 103.080 32.900 ;
        RECT 105.470 32.870 107.440 32.950 ;
      LAYER li1 ;
        RECT 107.620 32.870 107.880 36.130 ;
      LAYER li1 ;
        RECT 108.170 36.060 108.220 36.230 ;
        RECT 108.390 36.060 108.660 36.230 ;
        RECT 108.830 36.060 109.100 36.230 ;
        RECT 109.270 36.060 109.510 36.230 ;
        RECT 109.680 36.060 109.780 36.230 ;
        RECT 108.170 35.780 109.780 36.060 ;
        RECT 108.480 35.380 109.780 35.780 ;
        RECT 110.010 36.230 110.600 36.260 ;
        RECT 110.010 36.060 110.040 36.230 ;
        RECT 110.210 36.060 110.400 36.230 ;
        RECT 110.570 36.060 110.600 36.230 ;
        RECT 111.280 36.230 112.230 36.260 ;
        RECT 108.480 34.600 108.810 35.380 ;
        RECT 110.010 35.300 110.600 36.060 ;
      LAYER li1 ;
        RECT 110.850 35.200 111.100 36.130 ;
      LAYER li1 ;
        RECT 111.280 36.060 111.310 36.230 ;
        RECT 111.480 36.060 111.670 36.230 ;
        RECT 111.840 36.060 112.030 36.230 ;
        RECT 112.200 36.060 112.230 36.230 ;
        RECT 113.450 36.230 115.060 36.260 ;
        RECT 111.280 35.380 112.230 36.060 ;
      LAYER li1 ;
        RECT 112.410 35.200 112.680 36.130 ;
      LAYER li1 ;
        RECT 113.450 36.060 113.500 36.230 ;
        RECT 113.670 36.060 113.940 36.230 ;
        RECT 114.110 36.060 114.380 36.230 ;
        RECT 114.550 36.060 114.790 36.230 ;
        RECT 114.960 36.060 115.060 36.230 ;
        RECT 113.450 35.780 115.060 36.060 ;
        RECT 116.250 36.230 117.200 36.260 ;
        RECT 116.250 36.060 116.280 36.230 ;
        RECT 116.450 36.060 116.640 36.230 ;
        RECT 116.810 36.060 117.000 36.230 ;
        RECT 117.170 36.060 117.200 36.230 ;
        RECT 117.810 36.230 118.760 36.260 ;
        RECT 109.020 33.940 109.350 34.930 ;
      LAYER li1 ;
        RECT 110.050 34.510 110.350 35.100 ;
        RECT 110.850 35.030 112.680 35.200 ;
        RECT 110.530 34.510 111.720 34.850 ;
      LAYER li1 ;
        RECT 108.250 33.070 109.700 33.940 ;
        RECT 108.250 32.900 108.500 33.070 ;
        RECT 108.670 32.900 108.860 33.070 ;
        RECT 109.030 32.900 109.300 33.070 ;
        RECT 109.470 32.900 109.700 33.070 ;
        RECT 108.250 32.870 109.700 32.900 ;
        RECT 110.010 33.120 111.680 34.330 ;
      LAYER li1 ;
        RECT 111.900 33.370 112.230 34.850 ;
      LAYER li1 ;
        RECT 110.010 32.950 110.040 33.120 ;
        RECT 110.210 32.950 110.400 33.120 ;
        RECT 110.570 32.950 110.760 33.120 ;
        RECT 110.930 32.950 111.120 33.120 ;
        RECT 111.290 32.950 111.480 33.120 ;
        RECT 111.650 32.950 111.680 33.120 ;
        RECT 110.010 32.870 111.680 32.950 ;
      LAYER li1 ;
        RECT 112.410 32.870 112.680 35.030 ;
      LAYER li1 ;
        RECT 113.760 35.380 115.060 35.780 ;
        RECT 113.760 34.600 114.090 35.380 ;
        RECT 114.300 33.940 114.630 34.930 ;
        RECT 113.530 33.070 114.980 33.940 ;
      LAYER li1 ;
        RECT 115.830 33.770 116.000 35.790 ;
      LAYER li1 ;
        RECT 116.250 35.300 117.200 36.060 ;
      LAYER li1 ;
        RECT 117.380 35.420 117.630 36.130 ;
      LAYER li1 ;
        RECT 117.810 36.060 117.840 36.230 ;
        RECT 118.010 36.060 118.200 36.230 ;
        RECT 118.370 36.060 118.560 36.230 ;
        RECT 118.730 36.060 118.760 36.230 ;
        RECT 119.370 36.230 120.320 36.260 ;
        RECT 117.810 35.600 118.760 36.060 ;
      LAYER li1 ;
        RECT 118.940 35.420 119.190 36.130 ;
        RECT 117.380 35.250 119.190 35.420 ;
      LAYER li1 ;
        RECT 119.370 36.060 119.400 36.230 ;
        RECT 119.570 36.060 119.760 36.230 ;
        RECT 119.930 36.060 120.120 36.230 ;
        RECT 120.290 36.060 120.320 36.230 ;
        RECT 121.130 36.230 122.740 36.260 ;
        RECT 119.370 35.380 120.320 36.060 ;
      LAYER li1 ;
        RECT 117.380 35.080 117.550 35.250 ;
      LAYER li1 ;
        RECT 120.500 35.200 120.830 36.130 ;
        RECT 121.130 36.060 121.180 36.230 ;
        RECT 121.350 36.060 121.620 36.230 ;
        RECT 121.790 36.060 122.060 36.230 ;
        RECT 122.230 36.060 122.470 36.230 ;
        RECT 122.640 36.060 122.740 36.230 ;
        RECT 123.410 36.230 124.270 36.260 ;
        RECT 121.130 35.780 122.740 36.060 ;
      LAYER li1 ;
        RECT 116.290 34.850 117.550 35.080 ;
      LAYER li1 ;
        RECT 119.590 35.070 120.830 35.200 ;
        RECT 117.730 35.030 120.830 35.070 ;
        RECT 117.730 34.900 119.760 35.030 ;
      LAYER li1 ;
        RECT 117.380 34.720 117.550 34.850 ;
        RECT 117.380 34.550 119.270 34.720 ;
      LAYER li1 ;
        RECT 113.530 32.900 113.780 33.070 ;
        RECT 113.950 32.900 114.140 33.070 ;
        RECT 114.310 32.900 114.580 33.070 ;
        RECT 114.750 32.900 114.980 33.070 ;
        RECT 113.530 32.870 114.980 32.900 ;
        RECT 116.250 33.120 117.200 34.450 ;
        RECT 116.250 32.950 116.280 33.120 ;
        RECT 116.450 32.950 116.640 33.120 ;
        RECT 116.810 32.950 117.000 33.120 ;
        RECT 117.170 32.950 117.200 33.120 ;
        RECT 116.250 32.870 117.200 32.950 ;
      LAYER li1 ;
        RECT 117.380 32.870 117.630 34.550 ;
      LAYER li1 ;
        RECT 117.810 33.120 118.760 34.370 ;
        RECT 117.810 32.950 117.840 33.120 ;
        RECT 118.010 32.950 118.200 33.120 ;
        RECT 118.370 32.950 118.560 33.120 ;
        RECT 118.730 32.950 118.760 33.120 ;
        RECT 117.810 32.870 118.760 32.950 ;
      LAYER li1 ;
        RECT 118.940 32.870 119.270 34.550 ;
        RECT 120.050 34.510 120.380 34.850 ;
      LAYER li1 ;
        RECT 119.450 33.120 120.400 34.330 ;
        RECT 119.450 32.950 119.480 33.120 ;
        RECT 119.650 32.950 119.840 33.120 ;
        RECT 120.010 32.950 120.200 33.120 ;
        RECT 120.370 32.950 120.400 33.120 ;
        RECT 119.450 32.870 120.400 32.950 ;
        RECT 120.580 32.870 120.830 35.030 ;
        RECT 121.440 35.380 122.740 35.780 ;
        RECT 121.440 34.600 121.770 35.380 ;
        RECT 123.030 35.070 123.240 36.130 ;
        RECT 123.410 36.060 123.460 36.230 ;
        RECT 123.630 36.060 124.050 36.230 ;
        RECT 124.220 36.060 124.270 36.230 ;
        RECT 125.500 36.230 126.170 36.260 ;
        RECT 123.410 35.720 124.270 36.060 ;
        RECT 124.450 35.720 124.850 36.130 ;
        RECT 125.500 36.060 125.570 36.230 ;
        RECT 125.740 36.060 125.930 36.230 ;
        RECT 126.100 36.060 126.170 36.230 ;
        RECT 126.890 36.230 128.500 36.260 ;
      LAYER li1 ;
        RECT 123.410 35.240 124.200 35.550 ;
      LAYER li1 ;
        RECT 124.450 35.070 124.620 35.720 ;
      LAYER li1 ;
        RECT 124.800 35.240 125.330 35.550 ;
      LAYER li1 ;
        RECT 125.500 35.300 126.170 36.060 ;
        RECT 121.980 33.940 122.310 34.930 ;
        RECT 123.030 34.900 126.140 35.070 ;
        RECT 121.210 33.070 122.660 33.940 ;
        RECT 123.030 33.850 123.280 34.900 ;
      LAYER li1 ;
        RECT 123.490 33.370 124.420 34.720 ;
      LAYER li1 ;
        RECT 125.810 34.690 126.140 34.900 ;
        RECT 124.590 33.200 126.160 34.450 ;
        RECT 121.210 32.900 121.460 33.070 ;
        RECT 121.630 32.900 121.820 33.070 ;
        RECT 121.990 32.900 122.260 33.070 ;
        RECT 122.430 32.900 122.660 33.070 ;
        RECT 121.210 32.870 122.660 32.900 ;
        RECT 124.500 33.120 126.160 33.200 ;
        RECT 124.500 32.950 124.550 33.120 ;
        RECT 124.720 32.950 124.910 33.120 ;
        RECT 125.080 32.950 125.270 33.120 ;
        RECT 125.440 32.950 125.630 33.120 ;
        RECT 125.800 32.950 125.990 33.120 ;
        RECT 124.500 32.870 126.160 32.950 ;
      LAYER li1 ;
        RECT 126.340 32.870 126.600 36.130 ;
      LAYER li1 ;
        RECT 126.890 36.060 126.940 36.230 ;
        RECT 127.110 36.060 127.380 36.230 ;
        RECT 127.550 36.060 127.820 36.230 ;
        RECT 127.990 36.060 128.230 36.230 ;
        RECT 128.400 36.060 128.500 36.230 ;
        RECT 126.890 35.780 128.500 36.060 ;
        RECT 127.200 35.380 128.500 35.780 ;
        RECT 128.730 36.230 129.660 36.260 ;
        RECT 128.730 36.060 128.750 36.230 ;
        RECT 128.920 36.060 129.110 36.230 ;
        RECT 129.280 36.060 129.470 36.230 ;
        RECT 129.640 36.060 129.660 36.230 ;
        RECT 130.360 36.230 130.950 36.260 ;
        RECT 127.200 34.600 127.530 35.380 ;
        RECT 128.730 35.300 129.660 36.060 ;
      LAYER li1 ;
        RECT 129.840 35.200 130.170 36.130 ;
      LAYER li1 ;
        RECT 130.360 36.060 130.390 36.230 ;
        RECT 130.560 36.060 130.750 36.230 ;
        RECT 130.920 36.060 130.950 36.230 ;
        RECT 130.360 35.380 130.950 36.060 ;
        RECT 131.620 36.240 134.350 36.270 ;
        RECT 131.620 36.070 131.790 36.240 ;
        RECT 131.960 36.070 132.230 36.240 ;
        RECT 132.400 36.070 132.640 36.240 ;
        RECT 132.810 36.070 133.070 36.240 ;
        RECT 133.240 36.070 133.510 36.240 ;
        RECT 133.680 36.070 133.920 36.240 ;
        RECT 134.090 36.070 134.350 36.240 ;
        RECT 131.620 35.270 134.350 36.070 ;
        RECT 134.970 36.230 135.560 36.260 ;
        RECT 134.970 36.060 135.000 36.230 ;
        RECT 135.170 36.060 135.360 36.230 ;
        RECT 135.530 36.060 135.560 36.230 ;
        RECT 136.490 36.230 138.100 36.260 ;
        RECT 134.970 35.300 135.560 36.060 ;
      LAYER li1 ;
        RECT 129.840 35.030 130.920 35.200 ;
      LAYER li1 ;
        RECT 127.740 33.940 128.070 34.930 ;
      LAYER li1 ;
        RECT 128.770 34.510 129.960 34.850 ;
        RECT 130.140 34.510 130.470 34.850 ;
      LAYER li1 ;
        RECT 126.970 33.070 128.420 33.940 ;
        RECT 126.970 32.900 127.220 33.070 ;
        RECT 127.390 32.900 127.580 33.070 ;
        RECT 127.750 32.900 128.020 33.070 ;
        RECT 128.190 32.900 128.420 33.070 ;
        RECT 126.970 32.870 128.420 32.900 ;
        RECT 128.730 33.120 130.400 34.330 ;
        RECT 128.730 32.950 128.760 33.120 ;
        RECT 128.930 32.950 129.120 33.120 ;
        RECT 129.290 32.950 129.480 33.120 ;
        RECT 129.650 32.950 129.840 33.120 ;
        RECT 130.010 32.950 130.200 33.120 ;
        RECT 130.370 32.950 130.400 33.120 ;
        RECT 128.730 32.870 130.400 32.950 ;
      LAYER li1 ;
        RECT 130.660 32.870 130.920 35.030 ;
      LAYER li1 ;
        RECT 131.780 34.600 132.110 35.270 ;
        RECT 132.510 33.950 132.840 34.930 ;
        RECT 133.060 34.600 133.390 35.270 ;
        RECT 133.790 33.950 134.120 34.930 ;
      LAYER li1 ;
        RECT 135.010 34.690 135.720 35.080 ;
        RECT 135.900 34.450 136.230 36.130 ;
      LAYER li1 ;
        RECT 136.490 36.060 136.540 36.230 ;
        RECT 136.710 36.060 136.980 36.230 ;
        RECT 137.150 36.060 137.420 36.230 ;
        RECT 137.590 36.060 137.830 36.230 ;
        RECT 138.000 36.060 138.100 36.230 ;
        RECT 136.490 35.780 138.100 36.060 ;
        RECT 136.800 35.380 138.100 35.780 ;
        RECT 138.330 36.230 138.920 36.260 ;
        RECT 138.330 36.060 138.360 36.230 ;
        RECT 138.530 36.060 138.720 36.230 ;
        RECT 138.890 36.060 138.920 36.230 ;
        RECT 139.850 36.230 141.460 36.260 ;
        RECT 136.800 34.600 137.130 35.380 ;
        RECT 138.330 35.300 138.920 36.060 ;
        RECT 131.540 33.070 134.280 33.950 ;
        RECT 131.540 32.900 131.750 33.070 ;
        RECT 131.920 32.900 132.190 33.070 ;
        RECT 132.360 32.900 132.600 33.070 ;
        RECT 132.770 32.900 133.030 33.070 ;
        RECT 133.200 32.900 133.470 33.070 ;
        RECT 133.640 32.900 133.880 33.070 ;
        RECT 134.050 32.900 134.280 33.070 ;
        RECT 131.540 32.880 134.280 32.900 ;
        RECT 134.970 33.120 135.560 34.450 ;
        RECT 134.970 32.950 135.000 33.120 ;
        RECT 135.170 32.950 135.360 33.120 ;
        RECT 135.530 32.950 135.560 33.120 ;
        RECT 134.970 32.870 135.560 32.950 ;
      LAYER li1 ;
        RECT 135.840 32.870 136.230 34.450 ;
      LAYER li1 ;
        RECT 137.340 33.940 137.670 34.930 ;
      LAYER li1 ;
        RECT 138.370 34.690 139.080 35.080 ;
        RECT 139.260 34.450 139.590 36.130 ;
      LAYER li1 ;
        RECT 139.850 36.060 139.900 36.230 ;
        RECT 140.070 36.060 140.340 36.230 ;
        RECT 140.510 36.060 140.780 36.230 ;
        RECT 140.950 36.060 141.190 36.230 ;
        RECT 141.360 36.060 141.460 36.230 ;
        RECT 139.850 35.780 141.460 36.060 ;
        RECT 140.160 35.380 141.460 35.780 ;
        RECT 140.160 34.600 140.490 35.380 ;
        RECT 136.570 33.070 138.020 33.940 ;
        RECT 136.570 32.900 136.820 33.070 ;
        RECT 136.990 32.900 137.180 33.070 ;
        RECT 137.350 32.900 137.620 33.070 ;
        RECT 137.790 32.900 138.020 33.070 ;
        RECT 136.570 32.870 138.020 32.900 ;
        RECT 138.330 33.120 138.920 34.450 ;
        RECT 138.330 32.950 138.360 33.120 ;
        RECT 138.530 32.950 138.720 33.120 ;
        RECT 138.890 32.950 138.920 33.120 ;
        RECT 138.330 32.870 138.920 32.950 ;
      LAYER li1 ;
        RECT 139.200 32.870 139.590 34.450 ;
      LAYER li1 ;
        RECT 140.700 33.940 141.030 34.930 ;
        RECT 139.930 33.070 141.380 33.940 ;
        RECT 139.930 32.900 140.180 33.070 ;
        RECT 140.350 32.900 140.540 33.070 ;
        RECT 140.710 32.900 140.980 33.070 ;
        RECT 141.150 32.900 141.380 33.070 ;
        RECT 139.930 32.870 141.380 32.900 ;
        RECT 5.760 32.470 5.920 32.650 ;
        RECT 6.090 32.470 6.400 32.650 ;
        RECT 6.570 32.470 6.880 32.650 ;
        RECT 7.050 32.470 7.360 32.650 ;
        RECT 7.530 32.470 7.840 32.650 ;
        RECT 8.010 32.470 8.320 32.650 ;
        RECT 8.490 32.470 8.800 32.650 ;
        RECT 8.970 32.470 9.280 32.650 ;
        RECT 9.450 32.470 9.760 32.650 ;
        RECT 9.930 32.470 10.240 32.650 ;
        RECT 10.410 32.470 10.720 32.650 ;
        RECT 10.890 32.470 11.200 32.650 ;
        RECT 11.370 32.470 11.680 32.650 ;
        RECT 11.850 32.470 12.160 32.650 ;
        RECT 12.330 32.470 12.640 32.650 ;
        RECT 12.810 32.470 13.120 32.650 ;
        RECT 13.290 32.470 13.600 32.650 ;
        RECT 13.770 32.470 14.080 32.650 ;
        RECT 14.250 32.470 14.560 32.650 ;
        RECT 14.730 32.470 15.040 32.650 ;
        RECT 15.210 32.470 15.520 32.650 ;
        RECT 15.690 32.470 16.000 32.650 ;
        RECT 16.170 32.470 16.480 32.650 ;
        RECT 16.650 32.470 16.960 32.650 ;
        RECT 17.130 32.470 17.440 32.650 ;
        RECT 17.610 32.470 17.920 32.650 ;
        RECT 18.090 32.470 18.400 32.650 ;
        RECT 18.570 32.470 18.880 32.650 ;
        RECT 19.050 32.470 19.360 32.650 ;
        RECT 19.530 32.470 19.840 32.650 ;
        RECT 20.010 32.470 20.320 32.650 ;
        RECT 20.490 32.470 20.800 32.650 ;
        RECT 20.970 32.470 21.280 32.650 ;
        RECT 21.450 32.470 21.760 32.650 ;
        RECT 21.930 32.470 22.240 32.650 ;
        RECT 22.410 32.470 22.720 32.650 ;
        RECT 22.890 32.470 23.200 32.650 ;
        RECT 23.370 32.470 23.680 32.650 ;
        RECT 23.850 32.470 24.160 32.650 ;
        RECT 24.330 32.470 24.640 32.650 ;
        RECT 24.810 32.470 25.120 32.650 ;
        RECT 25.290 32.470 25.600 32.650 ;
        RECT 25.770 32.470 26.080 32.650 ;
        RECT 26.250 32.470 26.560 32.650 ;
        RECT 26.730 32.470 27.040 32.650 ;
        RECT 27.210 32.470 27.520 32.650 ;
        RECT 27.690 32.470 28.000 32.650 ;
        RECT 28.170 32.470 28.480 32.650 ;
        RECT 28.650 32.470 28.960 32.650 ;
        RECT 29.130 32.470 29.440 32.650 ;
        RECT 29.610 32.470 29.920 32.650 ;
        RECT 30.090 32.470 30.400 32.650 ;
        RECT 30.570 32.470 30.880 32.650 ;
        RECT 31.050 32.470 31.360 32.650 ;
        RECT 31.530 32.470 31.840 32.650 ;
        RECT 32.010 32.470 32.320 32.650 ;
        RECT 32.490 32.470 32.800 32.650 ;
        RECT 32.970 32.470 33.280 32.650 ;
        RECT 33.450 32.470 33.760 32.650 ;
        RECT 33.930 32.470 34.240 32.650 ;
        RECT 34.410 32.470 34.720 32.650 ;
        RECT 34.890 32.470 35.200 32.650 ;
        RECT 35.370 32.470 35.680 32.650 ;
        RECT 35.850 32.470 36.160 32.650 ;
        RECT 36.330 32.470 36.640 32.650 ;
        RECT 36.810 32.470 37.120 32.650 ;
        RECT 37.290 32.470 37.600 32.650 ;
        RECT 37.770 32.470 38.080 32.650 ;
        RECT 38.250 32.470 38.560 32.650 ;
        RECT 38.730 32.470 39.040 32.650 ;
        RECT 39.210 32.470 39.520 32.650 ;
        RECT 39.690 32.470 40.000 32.650 ;
        RECT 40.170 32.640 40.480 32.650 ;
        RECT 40.650 32.640 40.960 32.650 ;
        RECT 40.170 32.470 40.320 32.640 ;
        RECT 40.800 32.470 40.960 32.640 ;
        RECT 41.130 32.470 41.440 32.650 ;
        RECT 41.610 32.470 41.920 32.650 ;
        RECT 42.090 32.470 42.400 32.650 ;
        RECT 42.570 32.470 42.880 32.650 ;
        RECT 43.050 32.470 43.360 32.650 ;
        RECT 43.530 32.470 43.840 32.650 ;
        RECT 44.010 32.470 44.320 32.650 ;
        RECT 44.490 32.470 44.800 32.650 ;
        RECT 44.970 32.470 45.280 32.650 ;
        RECT 45.450 32.470 45.760 32.650 ;
        RECT 45.930 32.470 46.240 32.650 ;
        RECT 46.410 32.470 46.720 32.650 ;
        RECT 46.890 32.470 47.200 32.650 ;
        RECT 47.370 32.470 47.680 32.650 ;
        RECT 47.850 32.470 48.160 32.650 ;
        RECT 48.330 32.470 48.640 32.650 ;
        RECT 48.810 32.470 49.120 32.650 ;
        RECT 49.290 32.470 49.600 32.650 ;
        RECT 49.770 32.470 50.080 32.650 ;
        RECT 50.250 32.470 50.560 32.650 ;
        RECT 50.730 32.470 51.040 32.650 ;
        RECT 51.210 32.470 51.520 32.650 ;
        RECT 51.690 32.470 52.000 32.650 ;
        RECT 52.170 32.470 52.480 32.650 ;
        RECT 52.650 32.470 52.960 32.650 ;
        RECT 53.130 32.470 53.440 32.650 ;
        RECT 53.610 32.470 53.920 32.650 ;
        RECT 54.090 32.470 54.400 32.650 ;
        RECT 54.570 32.470 54.880 32.650 ;
        RECT 55.050 32.470 55.360 32.650 ;
        RECT 55.530 32.470 55.840 32.650 ;
        RECT 56.010 32.470 56.320 32.650 ;
        RECT 56.490 32.470 56.800 32.650 ;
        RECT 56.970 32.470 57.280 32.650 ;
        RECT 57.450 32.470 57.760 32.650 ;
        RECT 57.930 32.470 58.240 32.650 ;
        RECT 58.410 32.470 58.720 32.650 ;
        RECT 58.890 32.470 59.200 32.650 ;
        RECT 59.370 32.470 59.680 32.650 ;
        RECT 59.850 32.470 60.160 32.650 ;
        RECT 60.330 32.470 60.640 32.650 ;
        RECT 60.810 32.470 61.120 32.650 ;
        RECT 61.290 32.470 61.600 32.650 ;
        RECT 61.770 32.470 62.080 32.650 ;
        RECT 62.250 32.470 62.560 32.650 ;
        RECT 62.730 32.470 63.040 32.650 ;
        RECT 63.210 32.470 63.520 32.650 ;
        RECT 63.690 32.470 64.000 32.650 ;
        RECT 64.170 32.470 64.480 32.650 ;
        RECT 64.650 32.470 64.960 32.650 ;
        RECT 65.130 32.470 65.440 32.650 ;
        RECT 65.610 32.470 65.920 32.650 ;
        RECT 66.090 32.470 66.400 32.650 ;
        RECT 66.570 32.470 66.880 32.650 ;
        RECT 67.050 32.470 67.360 32.650 ;
        RECT 67.530 32.470 67.840 32.650 ;
        RECT 68.010 32.470 68.320 32.650 ;
        RECT 68.490 32.470 68.800 32.650 ;
        RECT 68.970 32.470 69.280 32.650 ;
        RECT 69.450 32.470 69.760 32.650 ;
        RECT 69.930 32.470 70.240 32.650 ;
        RECT 70.410 32.470 70.720 32.650 ;
        RECT 70.890 32.470 71.200 32.650 ;
        RECT 71.370 32.470 71.680 32.650 ;
        RECT 71.850 32.470 72.160 32.650 ;
        RECT 72.330 32.470 72.640 32.650 ;
        RECT 72.810 32.470 73.120 32.650 ;
        RECT 73.290 32.470 73.600 32.650 ;
        RECT 73.770 32.470 74.080 32.650 ;
        RECT 74.250 32.470 74.560 32.650 ;
        RECT 74.730 32.470 75.040 32.650 ;
        RECT 75.210 32.470 75.520 32.650 ;
        RECT 75.690 32.470 76.000 32.650 ;
        RECT 76.170 32.470 76.480 32.650 ;
        RECT 76.650 32.470 76.960 32.650 ;
        RECT 77.130 32.470 77.440 32.650 ;
        RECT 77.610 32.470 77.920 32.650 ;
        RECT 78.090 32.470 78.400 32.650 ;
        RECT 78.570 32.470 78.880 32.650 ;
        RECT 79.050 32.470 79.360 32.650 ;
        RECT 79.530 32.470 79.840 32.650 ;
        RECT 80.010 32.470 80.320 32.650 ;
        RECT 80.490 32.470 80.800 32.650 ;
        RECT 80.970 32.470 81.280 32.650 ;
        RECT 81.450 32.470 81.760 32.650 ;
        RECT 81.930 32.470 82.240 32.650 ;
        RECT 82.410 32.470 82.720 32.650 ;
        RECT 82.890 32.470 83.200 32.650 ;
        RECT 83.370 32.470 83.680 32.650 ;
        RECT 83.850 32.470 84.160 32.650 ;
        RECT 84.330 32.470 84.640 32.650 ;
        RECT 84.810 32.470 85.120 32.650 ;
        RECT 85.290 32.470 85.600 32.650 ;
        RECT 85.770 32.470 86.080 32.650 ;
        RECT 86.250 32.470 86.560 32.650 ;
        RECT 86.730 32.470 87.040 32.650 ;
        RECT 87.210 32.470 87.520 32.650 ;
        RECT 87.690 32.470 88.000 32.650 ;
        RECT 88.170 32.470 88.480 32.650 ;
        RECT 88.650 32.470 88.960 32.650 ;
        RECT 89.130 32.470 89.440 32.650 ;
        RECT 89.610 32.470 89.920 32.650 ;
        RECT 90.090 32.470 90.400 32.650 ;
        RECT 90.570 32.470 90.880 32.650 ;
        RECT 91.050 32.470 91.360 32.650 ;
        RECT 91.530 32.470 91.840 32.650 ;
        RECT 92.010 32.470 92.320 32.650 ;
        RECT 92.490 32.470 92.800 32.650 ;
        RECT 92.970 32.470 93.280 32.650 ;
        RECT 93.450 32.470 93.760 32.650 ;
        RECT 93.930 32.470 94.240 32.650 ;
        RECT 94.410 32.470 94.720 32.650 ;
        RECT 94.890 32.470 95.200 32.650 ;
        RECT 95.370 32.470 95.680 32.650 ;
        RECT 95.850 32.470 96.160 32.650 ;
        RECT 96.330 32.470 96.640 32.650 ;
        RECT 96.810 32.470 97.120 32.650 ;
        RECT 97.290 32.470 97.600 32.650 ;
        RECT 97.770 32.470 98.080 32.650 ;
        RECT 98.250 32.470 98.560 32.650 ;
        RECT 98.730 32.470 99.040 32.650 ;
        RECT 99.210 32.470 99.520 32.650 ;
        RECT 99.690 32.470 100.000 32.650 ;
        RECT 100.170 32.470 100.480 32.650 ;
        RECT 100.650 32.470 100.960 32.650 ;
        RECT 101.130 32.470 101.440 32.650 ;
        RECT 101.610 32.470 101.920 32.650 ;
        RECT 102.090 32.470 102.400 32.650 ;
        RECT 102.570 32.470 102.880 32.650 ;
        RECT 103.050 32.470 103.360 32.650 ;
        RECT 103.530 32.470 103.840 32.650 ;
        RECT 104.010 32.640 104.160 32.650 ;
        RECT 104.640 32.640 104.800 32.650 ;
        RECT 104.010 32.470 104.320 32.640 ;
        RECT 104.490 32.470 104.800 32.640 ;
        RECT 104.970 32.470 105.280 32.650 ;
        RECT 105.450 32.470 105.760 32.650 ;
        RECT 105.930 32.470 106.240 32.650 ;
        RECT 106.410 32.470 106.720 32.650 ;
        RECT 106.890 32.470 107.200 32.650 ;
        RECT 107.370 32.470 107.680 32.650 ;
        RECT 107.850 32.470 108.160 32.650 ;
        RECT 108.330 32.470 108.640 32.650 ;
        RECT 108.810 32.470 109.120 32.650 ;
        RECT 109.290 32.470 109.600 32.650 ;
        RECT 109.770 32.470 110.080 32.650 ;
        RECT 110.250 32.470 110.560 32.650 ;
        RECT 110.730 32.470 111.040 32.650 ;
        RECT 111.210 32.470 111.520 32.650 ;
        RECT 111.690 32.470 112.000 32.650 ;
        RECT 112.170 32.470 112.480 32.650 ;
        RECT 112.650 32.470 112.960 32.650 ;
        RECT 113.130 32.470 113.440 32.650 ;
        RECT 113.610 32.470 113.920 32.650 ;
        RECT 114.090 32.470 114.400 32.650 ;
        RECT 114.570 32.470 114.880 32.650 ;
        RECT 115.050 32.470 115.360 32.650 ;
        RECT 115.530 32.470 115.840 32.650 ;
        RECT 116.010 32.470 116.320 32.650 ;
        RECT 116.490 32.470 116.800 32.650 ;
        RECT 116.970 32.470 117.280 32.650 ;
        RECT 117.450 32.470 117.760 32.650 ;
        RECT 117.930 32.470 118.240 32.650 ;
        RECT 118.410 32.470 118.720 32.650 ;
        RECT 118.890 32.470 119.200 32.650 ;
        RECT 119.370 32.640 119.520 32.650 ;
        RECT 120.000 32.640 120.160 32.650 ;
        RECT 119.370 32.470 119.680 32.640 ;
        RECT 119.850 32.470 120.160 32.640 ;
        RECT 120.330 32.470 120.640 32.650 ;
        RECT 120.810 32.470 121.120 32.650 ;
        RECT 121.290 32.470 121.600 32.650 ;
        RECT 121.770 32.470 122.080 32.650 ;
        RECT 122.250 32.470 122.560 32.650 ;
        RECT 122.730 32.470 123.040 32.650 ;
        RECT 123.210 32.470 123.520 32.650 ;
        RECT 123.690 32.470 124.000 32.650 ;
        RECT 124.170 32.470 124.480 32.650 ;
        RECT 124.650 32.470 124.960 32.650 ;
        RECT 125.130 32.470 125.440 32.650 ;
        RECT 125.610 32.470 125.920 32.650 ;
        RECT 126.090 32.470 126.400 32.650 ;
        RECT 126.570 32.470 126.880 32.650 ;
        RECT 127.050 32.470 127.360 32.650 ;
        RECT 127.530 32.470 127.840 32.650 ;
        RECT 128.010 32.470 128.320 32.650 ;
        RECT 128.490 32.470 128.800 32.650 ;
        RECT 128.970 32.470 129.280 32.650 ;
        RECT 129.450 32.470 129.760 32.650 ;
        RECT 129.930 32.470 130.240 32.650 ;
        RECT 130.410 32.470 130.720 32.650 ;
        RECT 130.890 32.470 131.200 32.650 ;
        RECT 131.370 32.470 131.680 32.650 ;
        RECT 131.850 32.640 132.000 32.650 ;
        RECT 132.480 32.640 132.640 32.650 ;
        RECT 131.850 32.470 132.160 32.640 ;
        RECT 132.330 32.470 132.640 32.640 ;
        RECT 132.810 32.470 133.120 32.650 ;
        RECT 133.290 32.470 133.600 32.650 ;
        RECT 133.770 32.470 134.080 32.650 ;
        RECT 134.250 32.470 134.560 32.650 ;
        RECT 134.730 32.470 135.040 32.650 ;
        RECT 135.210 32.470 135.520 32.650 ;
        RECT 135.690 32.470 136.000 32.650 ;
        RECT 136.170 32.470 136.480 32.650 ;
        RECT 136.650 32.470 136.960 32.650 ;
        RECT 137.130 32.470 137.440 32.650 ;
        RECT 137.610 32.470 137.920 32.650 ;
        RECT 138.090 32.470 138.400 32.650 ;
        RECT 138.570 32.470 138.880 32.650 ;
        RECT 139.050 32.470 139.360 32.650 ;
        RECT 139.530 32.470 139.840 32.650 ;
        RECT 140.010 32.470 140.320 32.650 ;
        RECT 140.490 32.470 140.800 32.650 ;
        RECT 140.970 32.470 141.280 32.650 ;
        RECT 141.450 32.470 141.600 32.650 ;
        RECT 7.350 32.170 7.940 32.200 ;
        RECT 7.350 32.000 7.380 32.170 ;
        RECT 7.550 32.000 7.740 32.170 ;
        RECT 7.910 32.000 7.940 32.170 ;
        RECT 6.830 31.020 7.160 31.950 ;
        RECT 7.350 31.220 7.940 32.000 ;
        RECT 8.120 32.130 9.560 32.300 ;
        RECT 8.120 31.020 8.290 32.130 ;
        RECT 6.830 30.850 8.290 31.020 ;
        RECT 6.830 28.990 7.100 30.850 ;
        RECT 7.960 30.350 8.290 30.850 ;
        RECT 8.470 30.640 8.720 31.950 ;
        RECT 8.960 31.330 9.210 31.950 ;
        RECT 9.390 31.680 9.560 32.130 ;
        RECT 9.740 32.170 10.070 32.200 ;
        RECT 9.740 32.000 9.770 32.170 ;
        RECT 9.940 32.000 10.070 32.170 ;
        RECT 9.740 31.860 10.070 32.000 ;
        RECT 10.250 32.130 11.990 32.300 ;
        RECT 10.250 31.680 10.420 32.130 ;
        RECT 9.390 31.510 10.420 31.680 ;
        RECT 10.600 31.330 10.770 31.950 ;
        RECT 11.300 31.690 11.630 31.950 ;
        RECT 8.960 31.160 10.770 31.330 ;
        RECT 10.950 31.160 11.170 31.490 ;
        RECT 10.600 30.980 10.770 31.160 ;
        RECT 8.470 30.410 9.000 30.640 ;
        RECT 8.470 29.490 8.740 30.410 ;
      LAYER li1 ;
        RECT 9.420 30.110 9.960 30.980 ;
      LAYER li1 ;
        RECT 10.600 30.810 10.820 30.980 ;
        RECT 7.280 28.860 8.230 29.490 ;
        RECT 8.410 28.990 8.740 29.490 ;
        RECT 8.920 28.860 9.510 29.740 ;
      LAYER li1 ;
        RECT 9.790 29.120 9.960 30.110 ;
        RECT 10.140 29.300 10.470 30.600 ;
      LAYER li1 ;
        RECT 10.650 29.820 10.820 30.810 ;
        RECT 11.000 30.640 11.170 31.160 ;
        RECT 11.350 30.990 11.520 31.690 ;
        RECT 11.820 31.540 11.990 32.130 ;
        RECT 12.170 32.170 13.120 32.200 ;
        RECT 12.170 32.000 12.200 32.170 ;
        RECT 12.370 32.000 12.560 32.170 ;
        RECT 12.730 32.000 12.920 32.170 ;
        RECT 13.090 32.000 13.120 32.170 ;
        RECT 12.170 31.720 13.120 32.000 ;
        RECT 13.300 32.130 14.330 32.300 ;
        RECT 13.300 31.540 13.470 32.130 ;
        RECT 11.820 31.490 13.470 31.540 ;
        RECT 11.700 31.370 13.470 31.490 ;
        RECT 11.700 31.170 12.030 31.370 ;
        RECT 13.650 31.190 13.980 31.950 ;
        RECT 14.160 31.770 14.330 32.130 ;
        RECT 14.510 32.170 15.460 32.250 ;
        RECT 14.510 32.000 14.540 32.170 ;
        RECT 14.710 32.000 14.900 32.170 ;
        RECT 15.070 32.000 15.260 32.170 ;
        RECT 15.430 32.000 15.460 32.170 ;
        RECT 14.510 31.950 15.460 32.000 ;
        RECT 14.160 31.600 15.970 31.770 ;
        RECT 12.210 31.020 13.980 31.190 ;
        RECT 12.210 30.990 12.380 31.020 ;
        RECT 11.350 30.820 12.380 30.990 ;
        RECT 15.290 30.840 15.620 31.420 ;
        RECT 11.000 30.410 12.030 30.640 ;
        RECT 11.700 29.920 12.030 30.410 ;
        RECT 12.210 30.140 12.380 30.820 ;
        RECT 12.560 30.670 15.620 30.840 ;
        RECT 12.560 30.320 12.890 30.670 ;
      LAYER li1 ;
        RECT 13.330 30.320 15.180 30.490 ;
      LAYER li1 ;
        RECT 12.210 29.970 14.830 30.140 ;
        RECT 10.650 29.320 10.920 29.820 ;
        RECT 12.210 29.740 12.380 29.970 ;
      LAYER li1 ;
        RECT 15.010 29.790 15.180 30.320 ;
      LAYER li1 ;
        RECT 11.370 29.570 12.380 29.740 ;
      LAYER li1 ;
        RECT 12.560 29.620 15.180 29.790 ;
      LAYER li1 ;
        RECT 11.370 29.320 11.700 29.570 ;
      LAYER li1 ;
        RECT 12.560 29.120 12.730 29.620 ;
        RECT 9.790 28.950 12.730 29.120 ;
      LAYER li1 ;
        RECT 13.880 28.860 14.830 29.440 ;
      LAYER li1 ;
        RECT 15.010 28.930 15.180 29.620 ;
      LAYER li1 ;
        RECT 15.360 29.820 15.620 30.670 ;
        RECT 15.800 30.250 15.970 31.600 ;
        RECT 16.150 31.340 16.400 32.250 ;
        RECT 17.210 32.170 18.160 32.200 ;
        RECT 18.990 32.170 19.890 32.200 ;
        RECT 17.210 32.000 17.240 32.170 ;
        RECT 17.410 32.000 17.600 32.170 ;
        RECT 17.770 32.000 17.960 32.170 ;
        RECT 18.130 32.000 18.160 32.170 ;
        RECT 19.160 32.000 19.350 32.170 ;
        RECT 19.520 32.000 19.710 32.170 ;
        RECT 19.880 32.000 19.890 32.170 ;
        RECT 16.150 31.170 17.030 31.340 ;
        RECT 17.210 31.170 18.160 32.000 ;
        RECT 18.560 31.200 18.810 31.670 ;
        RECT 18.990 31.380 19.890 32.000 ;
        RECT 20.500 32.170 21.440 32.230 ;
        RECT 20.500 32.000 20.520 32.170 ;
        RECT 20.690 32.000 20.880 32.170 ;
        RECT 21.050 32.000 21.240 32.170 ;
        RECT 21.410 32.000 21.440 32.170 ;
        RECT 16.350 30.430 16.680 30.930 ;
        RECT 16.860 30.850 17.030 31.170 ;
        RECT 18.560 31.030 19.570 31.200 ;
        RECT 16.860 30.680 19.220 30.850 ;
        RECT 15.800 30.080 16.970 30.250 ;
        RECT 15.360 29.110 15.690 29.820 ;
        RECT 16.150 29.280 16.480 29.820 ;
        RECT 16.690 29.580 16.970 30.080 ;
        RECT 17.150 29.280 17.320 30.680 ;
        RECT 19.400 30.500 19.570 31.030 ;
        RECT 17.530 30.330 19.570 30.500 ;
        RECT 17.530 29.940 17.860 30.330 ;
      LAYER li1 ;
        RECT 18.180 29.760 18.510 30.150 ;
      LAYER li1 ;
        RECT 16.150 29.110 17.320 29.280 ;
      LAYER li1 ;
        RECT 17.500 29.590 18.510 29.760 ;
        RECT 17.500 28.930 17.670 29.590 ;
      LAYER li1 ;
        RECT 19.340 29.490 19.570 30.330 ;
        RECT 20.070 30.500 20.320 31.500 ;
        RECT 20.500 30.690 21.440 32.000 ;
        RECT 20.070 30.170 21.440 30.500 ;
        RECT 20.070 29.990 20.280 30.170 ;
        RECT 19.950 29.490 20.280 29.990 ;
      LAYER li1 ;
        RECT 15.010 28.760 17.670 28.930 ;
      LAYER li1 ;
        RECT 17.850 28.860 18.800 29.410 ;
        RECT 19.340 28.990 19.670 29.490 ;
        RECT 20.460 28.860 21.410 29.990 ;
      LAYER li1 ;
        RECT 21.620 29.160 21.960 32.230 ;
      LAYER li1 ;
        RECT 22.330 32.220 23.780 32.250 ;
        RECT 22.330 32.050 22.580 32.220 ;
        RECT 22.750 32.050 22.940 32.220 ;
        RECT 23.110 32.050 23.380 32.220 ;
        RECT 23.550 32.050 23.780 32.220 ;
        RECT 22.330 31.180 23.780 32.050 ;
        RECT 24.090 32.170 24.680 32.250 ;
        RECT 24.090 32.000 24.120 32.170 ;
        RECT 24.290 32.000 24.480 32.170 ;
        RECT 24.650 32.000 24.680 32.170 ;
        RECT 22.560 29.740 22.890 30.520 ;
        RECT 23.100 30.190 23.430 31.180 ;
        RECT 24.090 30.670 24.680 32.000 ;
      LAYER li1 ;
        RECT 24.960 30.670 25.350 32.250 ;
      LAYER li1 ;
        RECT 25.690 32.220 27.140 32.250 ;
        RECT 25.690 32.050 25.940 32.220 ;
        RECT 26.110 32.050 26.300 32.220 ;
        RECT 26.470 32.050 26.740 32.220 ;
        RECT 26.910 32.050 27.140 32.220 ;
        RECT 25.690 31.180 27.140 32.050 ;
      LAYER li1 ;
        RECT 24.130 30.040 24.840 30.430 ;
      LAYER li1 ;
        RECT 22.560 29.340 23.860 29.740 ;
        RECT 22.250 28.860 23.860 29.340 ;
        RECT 24.090 28.860 24.680 29.820 ;
      LAYER li1 ;
        RECT 25.020 28.990 25.350 30.670 ;
      LAYER li1 ;
        RECT 25.920 29.740 26.250 30.520 ;
        RECT 26.460 30.190 26.790 31.180 ;
        RECT 27.620 30.590 27.870 32.250 ;
        RECT 28.050 32.170 29.300 32.250 ;
        RECT 28.220 32.000 28.410 32.170 ;
        RECT 28.580 32.000 28.770 32.170 ;
        RECT 28.940 32.000 29.130 32.170 ;
        RECT 28.050 30.770 29.300 32.000 ;
        RECT 29.480 30.590 29.650 32.250 ;
        RECT 27.620 30.420 29.650 30.590 ;
      LAYER li1 ;
        RECT 29.830 30.300 30.160 31.750 ;
        RECT 27.490 30.000 28.680 30.240 ;
        RECT 28.930 30.000 29.280 30.240 ;
        RECT 30.340 30.120 30.600 32.250 ;
      LAYER li1 ;
        RECT 30.970 32.220 32.420 32.250 ;
        RECT 30.970 32.050 31.220 32.220 ;
        RECT 31.390 32.050 31.580 32.220 ;
        RECT 31.750 32.050 32.020 32.220 ;
        RECT 32.190 32.050 32.420 32.220 ;
        RECT 30.970 31.180 32.420 32.050 ;
      LAYER li1 ;
        RECT 29.580 29.950 30.600 30.120 ;
      LAYER li1 ;
        RECT 25.920 29.340 27.220 29.740 ;
        RECT 25.610 28.860 27.220 29.340 ;
        RECT 27.690 28.860 29.400 29.820 ;
      LAYER li1 ;
        RECT 29.580 28.990 29.830 29.950 ;
      LAYER li1 ;
        RECT 30.040 28.860 30.630 29.770 ;
        RECT 31.200 29.740 31.530 30.520 ;
        RECT 31.740 30.190 32.070 31.180 ;
        RECT 32.900 30.590 33.150 32.250 ;
        RECT 33.330 32.170 34.580 32.250 ;
        RECT 33.500 32.000 33.690 32.170 ;
        RECT 33.860 32.000 34.050 32.170 ;
        RECT 34.220 32.000 34.410 32.170 ;
        RECT 33.330 30.770 34.580 32.000 ;
        RECT 34.760 30.590 34.930 32.250 ;
        RECT 32.900 30.420 34.930 30.590 ;
      LAYER li1 ;
        RECT 35.110 30.300 35.440 31.750 ;
        RECT 32.770 30.000 33.960 30.240 ;
        RECT 34.210 30.000 34.560 30.240 ;
        RECT 35.620 30.120 35.880 32.250 ;
      LAYER li1 ;
        RECT 36.250 32.220 37.700 32.250 ;
        RECT 36.250 32.050 36.500 32.220 ;
        RECT 36.670 32.050 36.860 32.220 ;
        RECT 37.030 32.050 37.300 32.220 ;
        RECT 37.470 32.050 37.700 32.220 ;
        RECT 36.250 31.180 37.700 32.050 ;
        RECT 38.970 32.170 40.230 32.250 ;
        RECT 38.970 32.000 38.980 32.170 ;
        RECT 39.150 32.000 39.340 32.170 ;
        RECT 39.510 32.000 39.700 32.170 ;
        RECT 39.870 32.000 40.060 32.170 ;
      LAYER li1 ;
        RECT 34.860 29.950 35.880 30.120 ;
      LAYER li1 ;
        RECT 31.200 29.340 32.500 29.740 ;
        RECT 30.890 28.860 32.500 29.340 ;
        RECT 32.970 28.860 34.680 29.820 ;
      LAYER li1 ;
        RECT 34.860 28.990 35.110 29.950 ;
      LAYER li1 ;
        RECT 35.320 28.860 35.910 29.770 ;
        RECT 36.480 29.740 36.810 30.520 ;
        RECT 37.020 30.190 37.350 31.180 ;
        RECT 38.970 30.770 40.230 32.000 ;
      LAYER li1 ;
        RECT 40.760 31.750 40.930 32.250 ;
        RECT 40.410 30.670 40.930 31.750 ;
      LAYER li1 ;
        RECT 41.190 32.170 42.500 32.250 ;
        RECT 41.190 32.000 41.220 32.170 ;
        RECT 41.390 32.000 41.580 32.170 ;
        RECT 41.750 32.000 41.940 32.170 ;
        RECT 42.110 32.000 42.300 32.170 ;
        RECT 42.470 32.000 42.500 32.170 ;
        RECT 41.190 30.790 42.500 32.000 ;
        RECT 42.970 32.220 44.420 32.250 ;
        RECT 42.970 32.050 43.220 32.220 ;
        RECT 43.390 32.050 43.580 32.220 ;
        RECT 43.750 32.050 44.020 32.220 ;
        RECT 44.190 32.050 44.420 32.220 ;
        RECT 42.970 31.180 44.420 32.050 ;
        RECT 44.730 32.170 45.680 32.250 ;
        RECT 44.730 32.000 44.760 32.170 ;
        RECT 44.930 32.000 45.120 32.170 ;
        RECT 45.290 32.000 45.480 32.170 ;
        RECT 45.650 32.000 45.680 32.170 ;
      LAYER li1 ;
        RECT 40.410 30.590 40.680 30.670 ;
        RECT 39.620 30.420 40.680 30.590 ;
        RECT 39.010 30.030 39.430 30.360 ;
        RECT 39.620 29.850 39.790 30.420 ;
        RECT 41.130 30.300 41.640 30.610 ;
        RECT 41.890 30.300 42.600 30.610 ;
        RECT 39.970 30.030 40.480 30.240 ;
      LAYER li1 ;
        RECT 40.680 29.950 42.550 30.120 ;
        RECT 36.480 29.340 37.780 29.740 ;
        RECT 36.170 28.860 37.780 29.340 ;
        RECT 39.040 28.930 39.370 29.850 ;
      LAYER li1 ;
        RECT 39.620 29.500 40.150 29.850 ;
        RECT 39.620 29.330 40.160 29.500 ;
        RECT 39.620 29.110 40.150 29.330 ;
      LAYER li1 ;
        RECT 40.680 28.930 40.850 29.950 ;
        RECT 39.040 28.760 40.850 28.930 ;
        RECT 41.030 28.860 42.130 29.770 ;
        RECT 42.300 29.020 42.550 29.950 ;
        RECT 43.200 29.740 43.530 30.520 ;
        RECT 43.740 30.190 44.070 31.180 ;
        RECT 44.730 30.670 45.680 32.000 ;
      LAYER li1 ;
        RECT 45.860 30.570 46.110 32.250 ;
      LAYER li1 ;
        RECT 46.290 32.170 47.240 32.250 ;
        RECT 46.290 32.000 46.320 32.170 ;
        RECT 46.490 32.000 46.680 32.170 ;
        RECT 46.850 32.000 47.040 32.170 ;
        RECT 47.210 32.000 47.240 32.170 ;
        RECT 46.290 30.750 47.240 32.000 ;
      LAYER li1 ;
        RECT 47.420 30.570 47.750 32.250 ;
      LAYER li1 ;
        RECT 47.930 32.170 48.880 32.250 ;
        RECT 47.930 32.000 47.960 32.170 ;
        RECT 48.130 32.000 48.320 32.170 ;
        RECT 48.490 32.000 48.680 32.170 ;
        RECT 48.850 32.000 48.880 32.170 ;
        RECT 47.930 30.790 48.880 32.000 ;
      LAYER li1 ;
        RECT 45.860 30.400 47.750 30.570 ;
        RECT 45.860 30.270 46.030 30.400 ;
        RECT 48.530 30.270 48.860 30.610 ;
        RECT 44.770 30.040 46.030 30.270 ;
      LAYER li1 ;
        RECT 46.210 30.090 48.240 30.220 ;
        RECT 49.060 30.090 49.310 32.250 ;
        RECT 49.690 32.220 51.140 32.250 ;
        RECT 49.690 32.050 49.940 32.220 ;
        RECT 50.110 32.050 50.300 32.220 ;
        RECT 50.470 32.050 50.740 32.220 ;
        RECT 50.910 32.050 51.140 32.220 ;
        RECT 49.690 31.180 51.140 32.050 ;
        RECT 51.450 32.170 52.400 32.250 ;
        RECT 51.450 32.000 51.480 32.170 ;
        RECT 51.650 32.000 51.840 32.170 ;
        RECT 52.010 32.000 52.200 32.170 ;
        RECT 52.370 32.000 52.400 32.170 ;
        RECT 46.210 30.050 49.310 30.090 ;
      LAYER li1 ;
        RECT 45.860 29.870 46.030 30.040 ;
      LAYER li1 ;
        RECT 48.070 29.920 49.310 30.050 ;
        RECT 43.200 29.340 44.500 29.740 ;
        RECT 42.890 28.860 44.500 29.340 ;
        RECT 44.730 28.860 45.680 29.820 ;
      LAYER li1 ;
        RECT 45.860 29.700 47.670 29.870 ;
        RECT 45.860 28.990 46.110 29.700 ;
      LAYER li1 ;
        RECT 46.290 28.860 47.240 29.520 ;
      LAYER li1 ;
        RECT 47.420 28.990 47.670 29.700 ;
      LAYER li1 ;
        RECT 47.850 28.860 48.800 29.740 ;
        RECT 48.980 28.990 49.310 29.920 ;
        RECT 49.920 29.740 50.250 30.520 ;
        RECT 50.460 30.190 50.790 31.180 ;
        RECT 51.450 30.670 52.400 32.000 ;
      LAYER li1 ;
        RECT 52.580 30.570 52.830 32.250 ;
      LAYER li1 ;
        RECT 53.010 32.170 53.960 32.250 ;
        RECT 53.010 32.000 53.040 32.170 ;
        RECT 53.210 32.000 53.400 32.170 ;
        RECT 53.570 32.000 53.760 32.170 ;
        RECT 53.930 32.000 53.960 32.170 ;
        RECT 53.010 30.750 53.960 32.000 ;
      LAYER li1 ;
        RECT 54.140 30.570 54.470 32.250 ;
      LAYER li1 ;
        RECT 54.650 32.170 55.600 32.250 ;
        RECT 54.650 32.000 54.680 32.170 ;
        RECT 54.850 32.000 55.040 32.170 ;
        RECT 55.210 32.000 55.400 32.170 ;
        RECT 55.570 32.000 55.600 32.170 ;
        RECT 54.650 30.790 55.600 32.000 ;
      LAYER li1 ;
        RECT 52.580 30.400 54.470 30.570 ;
        RECT 52.580 30.270 52.750 30.400 ;
        RECT 55.250 30.270 55.580 30.610 ;
        RECT 51.490 30.040 52.750 30.270 ;
      LAYER li1 ;
        RECT 52.930 30.090 54.960 30.220 ;
        RECT 55.780 30.090 56.030 32.250 ;
        RECT 56.660 32.220 59.400 32.240 ;
        RECT 56.660 32.050 56.870 32.220 ;
        RECT 57.040 32.050 57.310 32.220 ;
        RECT 57.480 32.050 57.720 32.220 ;
        RECT 57.890 32.050 58.150 32.220 ;
        RECT 58.320 32.050 58.590 32.220 ;
        RECT 58.760 32.050 59.000 32.220 ;
        RECT 59.170 32.050 59.400 32.220 ;
        RECT 56.660 31.170 59.400 32.050 ;
        RECT 60.090 32.170 61.040 32.250 ;
        RECT 60.090 32.000 60.120 32.170 ;
        RECT 60.290 32.000 60.480 32.170 ;
        RECT 60.650 32.000 60.840 32.170 ;
        RECT 61.010 32.000 61.040 32.170 ;
        RECT 52.930 30.050 56.030 30.090 ;
      LAYER li1 ;
        RECT 52.580 29.870 52.750 30.040 ;
      LAYER li1 ;
        RECT 54.790 29.920 56.030 30.050 ;
        RECT 49.920 29.340 51.220 29.740 ;
        RECT 49.610 28.860 51.220 29.340 ;
        RECT 51.450 28.860 52.400 29.820 ;
      LAYER li1 ;
        RECT 52.580 29.700 54.390 29.870 ;
        RECT 52.580 28.990 52.830 29.700 ;
      LAYER li1 ;
        RECT 53.010 28.860 53.960 29.520 ;
      LAYER li1 ;
        RECT 54.140 28.990 54.390 29.700 ;
      LAYER li1 ;
        RECT 54.570 28.860 55.520 29.740 ;
        RECT 55.700 28.990 56.030 29.920 ;
        RECT 56.900 29.850 57.230 30.520 ;
        RECT 57.630 30.190 57.960 31.170 ;
        RECT 58.180 29.850 58.510 30.520 ;
        RECT 58.910 30.190 59.240 31.170 ;
        RECT 60.090 30.670 61.040 32.000 ;
      LAYER li1 ;
        RECT 61.220 30.570 61.470 32.250 ;
      LAYER li1 ;
        RECT 61.650 32.170 62.600 32.250 ;
        RECT 61.650 32.000 61.680 32.170 ;
        RECT 61.850 32.000 62.040 32.170 ;
        RECT 62.210 32.000 62.400 32.170 ;
        RECT 62.570 32.000 62.600 32.170 ;
        RECT 61.650 30.750 62.600 32.000 ;
      LAYER li1 ;
        RECT 62.780 30.570 63.110 32.250 ;
      LAYER li1 ;
        RECT 63.290 32.170 64.240 32.250 ;
        RECT 63.290 32.000 63.320 32.170 ;
        RECT 63.490 32.000 63.680 32.170 ;
        RECT 63.850 32.000 64.040 32.170 ;
        RECT 64.210 32.000 64.240 32.170 ;
        RECT 63.290 30.790 64.240 32.000 ;
      LAYER li1 ;
        RECT 61.220 30.400 63.110 30.570 ;
        RECT 61.220 30.270 61.390 30.400 ;
        RECT 63.890 30.270 64.220 30.610 ;
        RECT 60.130 30.040 61.390 30.270 ;
      LAYER li1 ;
        RECT 61.570 30.090 63.600 30.220 ;
        RECT 64.420 30.090 64.670 32.250 ;
        RECT 65.050 32.220 66.500 32.250 ;
        RECT 65.050 32.050 65.300 32.220 ;
        RECT 65.470 32.050 65.660 32.220 ;
        RECT 65.830 32.050 66.100 32.220 ;
        RECT 66.270 32.050 66.500 32.220 ;
        RECT 65.050 31.180 66.500 32.050 ;
        RECT 66.810 32.170 67.760 32.250 ;
        RECT 66.810 32.000 66.840 32.170 ;
        RECT 67.010 32.000 67.200 32.170 ;
        RECT 67.370 32.000 67.560 32.170 ;
        RECT 67.730 32.000 67.760 32.170 ;
        RECT 61.570 30.050 64.670 30.090 ;
      LAYER li1 ;
        RECT 61.220 29.870 61.390 30.040 ;
      LAYER li1 ;
        RECT 63.430 29.920 64.670 30.050 ;
        RECT 56.740 28.850 59.470 29.850 ;
        RECT 60.090 28.860 61.040 29.820 ;
      LAYER li1 ;
        RECT 61.220 29.700 63.030 29.870 ;
        RECT 61.220 28.990 61.470 29.700 ;
      LAYER li1 ;
        RECT 61.650 28.860 62.600 29.520 ;
      LAYER li1 ;
        RECT 62.780 28.990 63.030 29.700 ;
      LAYER li1 ;
        RECT 63.210 28.860 64.160 29.740 ;
        RECT 64.340 28.990 64.670 29.920 ;
        RECT 65.280 29.740 65.610 30.520 ;
        RECT 65.820 30.190 66.150 31.180 ;
        RECT 66.810 30.670 67.760 32.000 ;
      LAYER li1 ;
        RECT 67.940 30.570 68.190 32.250 ;
      LAYER li1 ;
        RECT 68.370 32.170 69.320 32.250 ;
        RECT 68.370 32.000 68.400 32.170 ;
        RECT 68.570 32.000 68.760 32.170 ;
        RECT 68.930 32.000 69.120 32.170 ;
        RECT 69.290 32.000 69.320 32.170 ;
        RECT 68.370 30.750 69.320 32.000 ;
      LAYER li1 ;
        RECT 69.500 30.570 69.830 32.250 ;
      LAYER li1 ;
        RECT 70.010 32.170 70.960 32.250 ;
        RECT 70.010 32.000 70.040 32.170 ;
        RECT 70.210 32.000 70.400 32.170 ;
        RECT 70.570 32.000 70.760 32.170 ;
        RECT 70.930 32.000 70.960 32.170 ;
        RECT 70.010 30.790 70.960 32.000 ;
      LAYER li1 ;
        RECT 67.940 30.400 69.830 30.570 ;
        RECT 67.940 30.270 68.110 30.400 ;
        RECT 70.610 30.270 70.940 30.610 ;
        RECT 66.850 30.040 68.110 30.270 ;
      LAYER li1 ;
        RECT 68.290 30.090 70.320 30.220 ;
        RECT 71.140 30.090 71.390 32.250 ;
        RECT 71.770 32.220 73.220 32.250 ;
        RECT 71.770 32.050 72.020 32.220 ;
        RECT 72.190 32.050 72.380 32.220 ;
        RECT 72.550 32.050 72.820 32.220 ;
        RECT 72.990 32.050 73.220 32.220 ;
        RECT 71.770 31.180 73.220 32.050 ;
        RECT 73.530 32.170 74.480 32.250 ;
        RECT 73.530 32.000 73.560 32.170 ;
        RECT 73.730 32.000 73.920 32.170 ;
        RECT 74.090 32.000 74.280 32.170 ;
        RECT 74.450 32.000 74.480 32.170 ;
        RECT 68.290 30.050 71.390 30.090 ;
      LAYER li1 ;
        RECT 67.940 29.870 68.110 30.040 ;
      LAYER li1 ;
        RECT 70.150 29.920 71.390 30.050 ;
        RECT 65.280 29.340 66.580 29.740 ;
        RECT 64.970 28.860 66.580 29.340 ;
        RECT 66.810 28.860 67.760 29.820 ;
      LAYER li1 ;
        RECT 67.940 29.700 69.750 29.870 ;
        RECT 67.940 28.990 68.190 29.700 ;
      LAYER li1 ;
        RECT 68.370 28.860 69.320 29.520 ;
      LAYER li1 ;
        RECT 69.500 28.990 69.750 29.700 ;
      LAYER li1 ;
        RECT 69.930 28.860 70.880 29.740 ;
        RECT 71.060 28.990 71.390 29.920 ;
        RECT 72.000 29.740 72.330 30.520 ;
        RECT 72.540 30.190 72.870 31.180 ;
        RECT 73.530 30.670 74.480 32.000 ;
      LAYER li1 ;
        RECT 74.660 30.570 74.910 32.250 ;
      LAYER li1 ;
        RECT 75.090 32.170 76.040 32.250 ;
        RECT 75.090 32.000 75.120 32.170 ;
        RECT 75.290 32.000 75.480 32.170 ;
        RECT 75.650 32.000 75.840 32.170 ;
        RECT 76.010 32.000 76.040 32.170 ;
        RECT 75.090 30.750 76.040 32.000 ;
      LAYER li1 ;
        RECT 76.220 30.570 76.550 32.250 ;
      LAYER li1 ;
        RECT 76.730 32.170 77.680 32.250 ;
        RECT 76.730 32.000 76.760 32.170 ;
        RECT 76.930 32.000 77.120 32.170 ;
        RECT 77.290 32.000 77.480 32.170 ;
        RECT 77.650 32.000 77.680 32.170 ;
        RECT 76.730 30.790 77.680 32.000 ;
      LAYER li1 ;
        RECT 74.660 30.400 76.550 30.570 ;
        RECT 74.660 30.270 74.830 30.400 ;
        RECT 77.330 30.270 77.660 30.610 ;
        RECT 73.570 30.040 74.830 30.270 ;
      LAYER li1 ;
        RECT 75.010 30.090 77.040 30.220 ;
        RECT 77.860 30.090 78.110 32.250 ;
        RECT 78.490 32.220 79.940 32.250 ;
        RECT 78.490 32.050 78.740 32.220 ;
        RECT 78.910 32.050 79.100 32.220 ;
        RECT 79.270 32.050 79.540 32.220 ;
        RECT 79.710 32.050 79.940 32.220 ;
        RECT 78.490 31.180 79.940 32.050 ;
        RECT 80.250 32.170 81.510 32.250 ;
        RECT 80.250 32.000 80.260 32.170 ;
        RECT 80.430 32.000 80.620 32.170 ;
        RECT 80.790 32.000 80.980 32.170 ;
        RECT 81.150 32.000 81.340 32.170 ;
        RECT 75.010 30.050 78.110 30.090 ;
      LAYER li1 ;
        RECT 74.660 29.870 74.830 30.040 ;
      LAYER li1 ;
        RECT 76.870 29.920 78.110 30.050 ;
        RECT 72.000 29.340 73.300 29.740 ;
        RECT 71.690 28.860 73.300 29.340 ;
        RECT 73.530 28.860 74.480 29.820 ;
      LAYER li1 ;
        RECT 74.660 29.700 76.470 29.870 ;
        RECT 74.660 28.990 74.910 29.700 ;
      LAYER li1 ;
        RECT 75.090 28.860 76.040 29.520 ;
      LAYER li1 ;
        RECT 76.220 28.990 76.470 29.700 ;
      LAYER li1 ;
        RECT 76.650 28.860 77.600 29.740 ;
        RECT 77.780 28.990 78.110 29.920 ;
        RECT 78.720 29.740 79.050 30.520 ;
        RECT 79.260 30.190 79.590 31.180 ;
        RECT 80.250 30.770 81.510 32.000 ;
      LAYER li1 ;
        RECT 82.040 31.750 82.210 32.250 ;
        RECT 81.690 30.670 82.210 31.750 ;
      LAYER li1 ;
        RECT 82.470 32.170 83.780 32.250 ;
        RECT 82.470 32.000 82.500 32.170 ;
        RECT 82.670 32.000 82.860 32.170 ;
        RECT 83.030 32.000 83.220 32.170 ;
        RECT 83.390 32.000 83.580 32.170 ;
        RECT 83.750 32.000 83.780 32.170 ;
        RECT 82.470 30.790 83.780 32.000 ;
        RECT 84.250 32.220 85.700 32.250 ;
        RECT 84.250 32.050 84.500 32.220 ;
        RECT 84.670 32.050 84.860 32.220 ;
        RECT 85.030 32.050 85.300 32.220 ;
        RECT 85.470 32.050 85.700 32.220 ;
        RECT 84.250 31.180 85.700 32.050 ;
        RECT 86.010 32.170 87.270 32.250 ;
        RECT 86.010 32.000 86.020 32.170 ;
        RECT 86.190 32.000 86.380 32.170 ;
        RECT 86.550 32.000 86.740 32.170 ;
        RECT 86.910 32.000 87.100 32.170 ;
      LAYER li1 ;
        RECT 81.690 30.590 81.960 30.670 ;
        RECT 80.900 30.420 81.960 30.590 ;
        RECT 80.290 30.030 80.710 30.360 ;
        RECT 80.900 29.850 81.070 30.420 ;
        RECT 82.410 30.300 82.920 30.610 ;
        RECT 83.170 30.300 83.880 30.610 ;
        RECT 81.250 30.030 81.760 30.240 ;
      LAYER li1 ;
        RECT 81.960 29.950 83.830 30.120 ;
        RECT 78.720 29.340 80.020 29.740 ;
        RECT 78.410 28.860 80.020 29.340 ;
        RECT 80.320 28.930 80.650 29.850 ;
      LAYER li1 ;
        RECT 80.900 29.500 81.430 29.850 ;
        RECT 80.900 29.330 81.440 29.500 ;
        RECT 80.900 29.110 81.430 29.330 ;
      LAYER li1 ;
        RECT 81.960 28.930 82.130 29.950 ;
        RECT 80.320 28.760 82.130 28.930 ;
        RECT 82.310 28.860 83.410 29.770 ;
        RECT 83.580 29.020 83.830 29.950 ;
        RECT 84.480 29.740 84.810 30.520 ;
        RECT 85.020 30.190 85.350 31.180 ;
        RECT 86.010 30.770 87.270 32.000 ;
      LAYER li1 ;
        RECT 87.800 31.750 87.970 32.250 ;
        RECT 87.450 30.670 87.970 31.750 ;
      LAYER li1 ;
        RECT 88.230 32.170 89.540 32.250 ;
        RECT 88.230 32.000 88.260 32.170 ;
        RECT 88.430 32.000 88.620 32.170 ;
        RECT 88.790 32.000 88.980 32.170 ;
        RECT 89.150 32.000 89.340 32.170 ;
        RECT 89.510 32.000 89.540 32.170 ;
        RECT 88.230 30.790 89.540 32.000 ;
        RECT 90.010 32.220 91.460 32.250 ;
        RECT 90.010 32.050 90.260 32.220 ;
        RECT 90.430 32.050 90.620 32.220 ;
        RECT 90.790 32.050 91.060 32.220 ;
        RECT 91.230 32.050 91.460 32.220 ;
        RECT 90.010 31.180 91.460 32.050 ;
      LAYER li1 ;
        RECT 87.450 30.590 87.720 30.670 ;
        RECT 86.660 30.420 87.720 30.590 ;
        RECT 86.050 30.030 86.470 30.360 ;
        RECT 86.660 29.850 86.830 30.420 ;
        RECT 88.170 30.300 88.680 30.610 ;
        RECT 88.930 30.300 89.640 30.610 ;
        RECT 87.010 30.030 87.520 30.240 ;
      LAYER li1 ;
        RECT 87.720 29.950 89.590 30.120 ;
        RECT 84.480 29.340 85.780 29.740 ;
        RECT 84.170 28.860 85.780 29.340 ;
        RECT 86.080 28.930 86.410 29.850 ;
      LAYER li1 ;
        RECT 86.660 29.500 87.190 29.850 ;
        RECT 86.660 29.330 87.200 29.500 ;
        RECT 86.660 29.110 87.190 29.330 ;
      LAYER li1 ;
        RECT 87.720 28.930 87.890 29.950 ;
        RECT 86.080 28.760 87.890 28.930 ;
        RECT 88.070 28.860 89.170 29.770 ;
        RECT 89.340 29.020 89.590 29.950 ;
        RECT 90.240 29.740 90.570 30.520 ;
        RECT 90.780 30.190 91.110 31.180 ;
        RECT 90.240 29.340 91.540 29.740 ;
        RECT 89.930 28.860 91.540 29.340 ;
      LAYER li1 ;
        RECT 91.810 28.990 92.060 32.250 ;
      LAYER li1 ;
        RECT 92.240 32.170 94.930 32.250 ;
        RECT 92.410 32.000 92.600 32.170 ;
        RECT 92.770 32.000 92.960 32.170 ;
        RECT 93.130 32.000 93.320 32.170 ;
        RECT 93.490 32.000 93.680 32.170 ;
        RECT 93.850 32.000 94.040 32.170 ;
        RECT 94.210 32.000 94.400 32.170 ;
        RECT 94.570 32.000 94.760 32.170 ;
        RECT 92.240 31.140 94.930 32.000 ;
        RECT 95.110 30.960 95.360 32.250 ;
        RECT 92.270 30.790 95.360 30.960 ;
        RECT 92.270 30.090 92.600 30.790 ;
        RECT 95.110 30.670 95.360 30.790 ;
        RECT 95.540 32.170 96.850 32.230 ;
        RECT 95.540 32.000 95.570 32.170 ;
        RECT 95.740 32.000 95.930 32.170 ;
        RECT 96.100 32.000 96.290 32.170 ;
        RECT 96.460 32.000 96.650 32.170 ;
        RECT 96.820 32.000 96.850 32.170 ;
        RECT 95.540 30.690 96.850 32.000 ;
        RECT 97.210 32.220 98.660 32.250 ;
        RECT 97.210 32.050 97.460 32.220 ;
        RECT 97.630 32.050 97.820 32.220 ;
        RECT 97.990 32.050 98.260 32.220 ;
        RECT 98.430 32.050 98.660 32.220 ;
        RECT 99.710 32.170 101.680 32.250 ;
        RECT 97.210 31.180 98.660 32.050 ;
        RECT 99.880 32.000 100.070 32.170 ;
        RECT 100.240 32.000 100.430 32.170 ;
        RECT 100.600 32.000 100.790 32.170 ;
        RECT 100.960 32.000 101.150 32.170 ;
        RECT 101.320 32.000 101.510 32.170 ;
      LAYER li1 ;
        RECT 93.100 30.270 93.830 30.550 ;
      LAYER li1 ;
        RECT 92.270 29.920 93.480 30.090 ;
        RECT 92.240 28.860 93.130 29.740 ;
        RECT 93.310 29.710 93.480 29.920 ;
      LAYER li1 ;
        RECT 93.660 30.060 93.830 30.270 ;
        RECT 94.010 30.240 94.440 30.610 ;
        RECT 94.640 30.070 94.930 30.610 ;
        RECT 95.170 30.070 95.880 30.400 ;
        RECT 96.230 30.240 96.560 30.510 ;
        RECT 96.150 30.070 96.560 30.240 ;
        RECT 93.660 29.890 94.460 30.060 ;
        RECT 96.230 29.890 96.560 30.070 ;
        RECT 94.290 29.720 96.560 29.890 ;
      LAYER li1 ;
        RECT 97.440 29.740 97.770 30.520 ;
        RECT 97.980 30.190 98.310 31.180 ;
        RECT 99.280 30.570 99.530 31.170 ;
        RECT 99.710 30.750 101.680 32.000 ;
        RECT 99.280 30.400 101.660 30.570 ;
        RECT 93.310 29.540 94.110 29.710 ;
      LAYER li1 ;
        RECT 94.720 29.700 95.390 29.720 ;
      LAYER li1 ;
        RECT 93.940 29.370 94.540 29.540 ;
        RECT 93.430 28.930 93.760 29.360 ;
        RECT 94.210 29.110 94.540 29.370 ;
        RECT 95.030 28.930 95.360 29.520 ;
        RECT 93.430 28.760 95.360 28.930 ;
        RECT 95.570 28.860 96.870 29.540 ;
        RECT 97.440 29.340 98.740 29.740 ;
      LAYER li1 ;
        RECT 99.490 29.670 99.820 30.220 ;
      LAYER li1 ;
        RECT 100.060 29.490 100.230 30.400 ;
        RECT 101.330 30.220 101.660 30.400 ;
      LAYER li1 ;
        RECT 100.410 29.670 100.740 30.220 ;
      LAYER li1 ;
        RECT 97.130 28.860 98.740 29.340 ;
        RECT 98.970 28.860 99.880 29.490 ;
        RECT 100.060 28.990 100.390 29.490 ;
        RECT 100.920 28.860 101.510 29.820 ;
      LAYER li1 ;
        RECT 101.860 28.990 102.120 32.250 ;
      LAYER li1 ;
        RECT 102.490 32.220 103.940 32.250 ;
        RECT 102.490 32.050 102.740 32.220 ;
        RECT 102.910 32.050 103.100 32.220 ;
        RECT 103.270 32.050 103.540 32.220 ;
        RECT 103.710 32.050 103.940 32.220 ;
        RECT 102.490 31.180 103.940 32.050 ;
        RECT 104.730 32.170 105.990 32.250 ;
        RECT 104.730 32.000 104.740 32.170 ;
        RECT 104.910 32.000 105.100 32.170 ;
        RECT 105.270 32.000 105.460 32.170 ;
        RECT 105.630 32.000 105.820 32.170 ;
        RECT 102.720 29.740 103.050 30.520 ;
        RECT 103.260 30.190 103.590 31.180 ;
        RECT 104.730 30.770 105.990 32.000 ;
      LAYER li1 ;
        RECT 106.520 31.750 106.690 32.250 ;
        RECT 106.170 30.670 106.690 31.750 ;
      LAYER li1 ;
        RECT 106.950 32.170 108.260 32.250 ;
        RECT 106.950 32.000 106.980 32.170 ;
        RECT 107.150 32.000 107.340 32.170 ;
        RECT 107.510 32.000 107.700 32.170 ;
        RECT 107.870 32.000 108.060 32.170 ;
        RECT 108.230 32.000 108.260 32.170 ;
        RECT 106.950 30.790 108.260 32.000 ;
        RECT 108.730 32.220 110.180 32.250 ;
        RECT 108.730 32.050 108.980 32.220 ;
        RECT 109.150 32.050 109.340 32.220 ;
        RECT 109.510 32.050 109.780 32.220 ;
        RECT 109.950 32.050 110.180 32.220 ;
        RECT 108.730 31.180 110.180 32.050 ;
      LAYER li1 ;
        RECT 106.170 30.590 106.440 30.670 ;
        RECT 105.380 30.420 106.440 30.590 ;
        RECT 104.770 30.030 105.190 30.360 ;
        RECT 105.380 29.850 105.550 30.420 ;
        RECT 106.890 30.300 107.400 30.610 ;
        RECT 107.650 30.300 108.360 30.610 ;
        RECT 105.730 30.030 106.240 30.240 ;
      LAYER li1 ;
        RECT 106.440 29.950 108.310 30.120 ;
        RECT 102.720 29.340 104.020 29.740 ;
        RECT 102.410 28.860 104.020 29.340 ;
        RECT 104.800 28.930 105.130 29.850 ;
      LAYER li1 ;
        RECT 105.380 29.500 105.910 29.850 ;
        RECT 105.380 29.330 105.920 29.500 ;
        RECT 105.380 29.110 105.910 29.330 ;
      LAYER li1 ;
        RECT 106.440 28.930 106.610 29.950 ;
        RECT 104.800 28.760 106.610 28.930 ;
        RECT 106.790 28.860 107.890 29.770 ;
        RECT 108.060 29.020 108.310 29.950 ;
        RECT 108.960 29.740 109.290 30.520 ;
        RECT 109.500 30.190 109.830 31.180 ;
        RECT 108.960 29.340 110.260 29.740 ;
        RECT 108.650 28.860 110.260 29.340 ;
      LAYER li1 ;
        RECT 110.530 28.990 110.780 32.250 ;
      LAYER li1 ;
        RECT 110.960 32.170 113.650 32.250 ;
        RECT 111.130 32.000 111.320 32.170 ;
        RECT 111.490 32.000 111.680 32.170 ;
        RECT 111.850 32.000 112.040 32.170 ;
        RECT 112.210 32.000 112.400 32.170 ;
        RECT 112.570 32.000 112.760 32.170 ;
        RECT 112.930 32.000 113.120 32.170 ;
        RECT 113.290 32.000 113.480 32.170 ;
        RECT 110.960 31.140 113.650 32.000 ;
        RECT 113.830 30.960 114.080 32.250 ;
        RECT 110.990 30.790 114.080 30.960 ;
        RECT 110.990 30.090 111.320 30.790 ;
        RECT 113.830 30.670 114.080 30.790 ;
        RECT 114.260 32.170 115.570 32.230 ;
        RECT 114.260 32.000 114.290 32.170 ;
        RECT 114.460 32.000 114.650 32.170 ;
        RECT 114.820 32.000 115.010 32.170 ;
        RECT 115.180 32.000 115.370 32.170 ;
        RECT 115.540 32.000 115.570 32.170 ;
        RECT 114.260 30.690 115.570 32.000 ;
        RECT 116.180 32.220 118.920 32.240 ;
        RECT 116.180 32.050 116.390 32.220 ;
        RECT 116.560 32.050 116.830 32.220 ;
        RECT 117.000 32.050 117.240 32.220 ;
        RECT 117.410 32.050 117.670 32.220 ;
        RECT 117.840 32.050 118.110 32.220 ;
        RECT 118.280 32.050 118.520 32.220 ;
        RECT 118.690 32.050 118.920 32.220 ;
        RECT 116.180 31.170 118.920 32.050 ;
        RECT 120.090 32.170 121.350 32.250 ;
        RECT 120.090 32.000 120.100 32.170 ;
        RECT 120.270 32.000 120.460 32.170 ;
        RECT 120.630 32.000 120.820 32.170 ;
        RECT 120.990 32.000 121.180 32.170 ;
      LAYER li1 ;
        RECT 111.820 30.270 112.550 30.550 ;
      LAYER li1 ;
        RECT 110.990 29.920 112.200 30.090 ;
        RECT 110.960 28.860 111.850 29.740 ;
        RECT 112.030 29.710 112.200 29.920 ;
      LAYER li1 ;
        RECT 112.380 30.060 112.550 30.270 ;
        RECT 112.730 30.240 113.160 30.610 ;
        RECT 113.360 30.070 113.650 30.610 ;
        RECT 113.890 30.070 114.600 30.400 ;
        RECT 112.380 29.890 113.180 30.060 ;
        RECT 114.950 29.890 115.280 30.510 ;
        RECT 113.010 29.720 115.280 29.890 ;
      LAYER li1 ;
        RECT 116.420 29.850 116.750 30.520 ;
        RECT 117.150 30.190 117.480 31.170 ;
        RECT 117.700 29.850 118.030 30.520 ;
        RECT 118.430 30.190 118.760 31.170 ;
        RECT 120.090 30.770 121.350 32.000 ;
      LAYER li1 ;
        RECT 121.880 31.750 122.050 32.250 ;
        RECT 121.530 30.670 122.050 31.750 ;
      LAYER li1 ;
        RECT 122.310 32.170 123.620 32.250 ;
        RECT 122.310 32.000 122.340 32.170 ;
        RECT 122.510 32.000 122.700 32.170 ;
        RECT 122.870 32.000 123.060 32.170 ;
        RECT 123.230 32.000 123.420 32.170 ;
        RECT 123.590 32.000 123.620 32.170 ;
        RECT 122.310 30.790 123.620 32.000 ;
        RECT 124.090 32.220 125.540 32.250 ;
        RECT 124.090 32.050 124.340 32.220 ;
        RECT 124.510 32.050 124.700 32.220 ;
        RECT 124.870 32.050 125.140 32.220 ;
        RECT 125.310 32.050 125.540 32.220 ;
        RECT 124.090 31.180 125.540 32.050 ;
        RECT 125.850 32.170 126.800 32.250 ;
        RECT 125.850 32.000 125.880 32.170 ;
        RECT 126.050 32.000 126.240 32.170 ;
        RECT 126.410 32.000 126.600 32.170 ;
        RECT 126.770 32.000 126.800 32.170 ;
      LAYER li1 ;
        RECT 121.530 30.590 121.800 30.670 ;
        RECT 120.740 30.420 121.800 30.590 ;
        RECT 120.130 30.030 120.550 30.360 ;
        RECT 120.740 29.850 120.910 30.420 ;
        RECT 122.250 30.300 122.760 30.610 ;
        RECT 123.010 30.300 123.720 30.610 ;
        RECT 121.090 30.030 121.600 30.240 ;
      LAYER li1 ;
        RECT 121.800 29.950 123.670 30.120 ;
        RECT 112.030 29.540 112.830 29.710 ;
      LAYER li1 ;
        RECT 113.440 29.700 114.110 29.720 ;
      LAYER li1 ;
        RECT 112.660 29.370 113.260 29.540 ;
        RECT 112.150 28.930 112.480 29.360 ;
        RECT 112.930 29.110 113.260 29.370 ;
        RECT 113.750 28.930 114.080 29.520 ;
        RECT 112.150 28.760 114.080 28.930 ;
        RECT 114.290 28.860 115.590 29.540 ;
        RECT 116.260 28.850 118.990 29.850 ;
        RECT 120.160 28.930 120.490 29.850 ;
      LAYER li1 ;
        RECT 120.740 29.500 121.270 29.850 ;
        RECT 120.740 29.330 121.280 29.500 ;
        RECT 120.740 29.110 121.270 29.330 ;
      LAYER li1 ;
        RECT 121.800 28.930 121.970 29.950 ;
        RECT 120.160 28.760 121.970 28.930 ;
        RECT 122.150 28.860 123.250 29.770 ;
        RECT 123.420 29.020 123.670 29.950 ;
        RECT 124.320 29.740 124.650 30.520 ;
        RECT 124.860 30.190 125.190 31.180 ;
        RECT 125.850 30.670 126.800 32.000 ;
      LAYER li1 ;
        RECT 125.890 30.040 126.780 30.430 ;
        RECT 126.980 30.190 127.230 32.250 ;
      LAYER li1 ;
        RECT 127.420 32.170 128.010 32.250 ;
        RECT 127.420 32.000 127.450 32.170 ;
        RECT 127.620 32.000 127.810 32.170 ;
        RECT 127.980 32.000 128.010 32.170 ;
        RECT 127.420 30.670 128.010 32.000 ;
        RECT 128.660 32.220 131.400 32.240 ;
        RECT 128.660 32.050 128.870 32.220 ;
        RECT 129.040 32.050 129.310 32.220 ;
        RECT 129.480 32.050 129.720 32.220 ;
        RECT 129.890 32.050 130.150 32.220 ;
        RECT 130.320 32.050 130.590 32.220 ;
        RECT 130.760 32.050 131.000 32.220 ;
        RECT 131.170 32.050 131.400 32.220 ;
        RECT 128.660 31.170 131.400 32.050 ;
        RECT 132.570 32.170 133.160 32.250 ;
        RECT 132.570 32.000 132.600 32.170 ;
        RECT 132.770 32.000 132.960 32.170 ;
        RECT 133.130 32.000 133.160 32.170 ;
      LAYER li1 ;
        RECT 126.980 30.020 127.560 30.190 ;
        RECT 127.740 30.020 128.040 30.350 ;
        RECT 127.340 29.840 127.560 30.020 ;
      LAYER li1 ;
        RECT 128.900 29.850 129.230 30.520 ;
        RECT 129.630 30.190 129.960 31.170 ;
        RECT 130.180 29.850 130.510 30.520 ;
        RECT 130.910 30.190 131.240 31.170 ;
        RECT 132.570 30.670 133.160 32.000 ;
      LAYER li1 ;
        RECT 133.440 30.670 133.830 32.250 ;
      LAYER li1 ;
        RECT 134.420 32.220 137.160 32.240 ;
        RECT 134.420 32.050 134.630 32.220 ;
        RECT 134.800 32.050 135.070 32.220 ;
        RECT 135.240 32.050 135.480 32.220 ;
        RECT 135.650 32.050 135.910 32.220 ;
        RECT 136.080 32.050 136.350 32.220 ;
        RECT 136.520 32.050 136.760 32.220 ;
        RECT 136.930 32.050 137.160 32.220 ;
        RECT 134.420 31.170 137.160 32.050 ;
        RECT 138.260 32.220 141.000 32.240 ;
        RECT 138.260 32.050 138.470 32.220 ;
        RECT 138.640 32.050 138.910 32.220 ;
        RECT 139.080 32.050 139.320 32.220 ;
        RECT 139.490 32.050 139.750 32.220 ;
        RECT 139.920 32.050 140.190 32.220 ;
        RECT 140.360 32.050 140.600 32.220 ;
        RECT 140.770 32.050 141.000 32.220 ;
        RECT 138.260 31.170 141.000 32.050 ;
      LAYER li1 ;
        RECT 132.610 30.040 133.320 30.430 ;
      LAYER li1 ;
        RECT 124.320 29.340 125.620 29.740 ;
        RECT 124.010 28.860 125.620 29.340 ;
        RECT 125.850 28.860 127.160 29.840 ;
      LAYER li1 ;
        RECT 127.340 29.670 127.940 29.840 ;
        RECT 127.610 29.010 127.940 29.670 ;
      LAYER li1 ;
        RECT 128.740 28.850 131.470 29.850 ;
        RECT 132.570 28.860 133.160 29.820 ;
      LAYER li1 ;
        RECT 133.500 28.990 133.830 30.670 ;
      LAYER li1 ;
        RECT 134.660 29.850 134.990 30.520 ;
        RECT 135.390 30.190 135.720 31.170 ;
        RECT 135.940 29.850 136.270 30.520 ;
        RECT 136.670 30.190 137.000 31.170 ;
        RECT 138.500 29.850 138.830 30.520 ;
        RECT 139.230 30.190 139.560 31.170 ;
        RECT 139.780 29.850 140.110 30.520 ;
        RECT 140.510 30.190 140.840 31.170 ;
        RECT 134.500 28.850 137.230 29.850 ;
        RECT 138.340 28.850 141.070 29.850 ;
        RECT 5.760 28.400 5.920 28.580 ;
        RECT 6.090 28.400 6.400 28.580 ;
        RECT 6.570 28.400 6.880 28.580 ;
        RECT 7.050 28.400 7.360 28.580 ;
        RECT 7.530 28.400 7.840 28.580 ;
        RECT 8.010 28.400 8.320 28.580 ;
        RECT 8.490 28.400 8.800 28.580 ;
        RECT 8.970 28.400 9.280 28.580 ;
        RECT 9.450 28.400 9.760 28.580 ;
        RECT 9.930 28.400 10.240 28.580 ;
        RECT 10.410 28.400 10.720 28.580 ;
        RECT 10.890 28.400 11.200 28.580 ;
        RECT 11.370 28.400 11.680 28.580 ;
        RECT 11.850 28.400 12.160 28.580 ;
        RECT 12.330 28.400 12.640 28.580 ;
        RECT 12.810 28.400 13.120 28.580 ;
        RECT 13.290 28.400 13.600 28.580 ;
        RECT 13.770 28.400 14.080 28.580 ;
        RECT 14.250 28.400 14.560 28.580 ;
        RECT 14.730 28.400 15.040 28.580 ;
        RECT 15.210 28.400 15.520 28.580 ;
        RECT 15.690 28.400 16.000 28.580 ;
        RECT 16.170 28.400 16.480 28.580 ;
        RECT 16.650 28.400 16.960 28.580 ;
        RECT 17.130 28.400 17.440 28.580 ;
        RECT 17.610 28.400 17.920 28.580 ;
        RECT 18.090 28.400 18.400 28.580 ;
        RECT 18.570 28.400 18.880 28.580 ;
        RECT 19.050 28.400 19.360 28.580 ;
        RECT 19.530 28.400 19.840 28.580 ;
        RECT 20.010 28.400 20.320 28.580 ;
        RECT 20.490 28.400 20.800 28.580 ;
        RECT 20.970 28.400 21.280 28.580 ;
        RECT 21.450 28.400 21.760 28.580 ;
        RECT 21.930 28.400 22.240 28.580 ;
        RECT 22.410 28.400 22.720 28.580 ;
        RECT 22.890 28.400 23.200 28.580 ;
        RECT 23.370 28.400 23.680 28.580 ;
        RECT 23.850 28.400 24.160 28.580 ;
        RECT 24.330 28.400 24.640 28.580 ;
        RECT 24.810 28.400 25.120 28.580 ;
        RECT 25.290 28.400 25.600 28.580 ;
        RECT 25.770 28.400 26.080 28.580 ;
        RECT 26.250 28.400 26.560 28.580 ;
        RECT 26.730 28.400 27.040 28.580 ;
        RECT 27.210 28.400 27.520 28.580 ;
        RECT 27.690 28.400 28.000 28.580 ;
        RECT 28.170 28.400 28.480 28.580 ;
        RECT 28.650 28.400 28.960 28.580 ;
        RECT 29.130 28.400 29.440 28.580 ;
        RECT 29.610 28.400 29.920 28.580 ;
        RECT 30.090 28.400 30.400 28.580 ;
        RECT 30.570 28.400 30.880 28.580 ;
        RECT 31.050 28.400 31.360 28.580 ;
        RECT 31.530 28.400 31.840 28.580 ;
        RECT 32.010 28.400 32.320 28.580 ;
        RECT 32.490 28.400 32.800 28.580 ;
        RECT 32.970 28.400 33.280 28.580 ;
        RECT 33.450 28.400 33.760 28.580 ;
        RECT 33.930 28.400 34.240 28.580 ;
        RECT 34.410 28.400 34.720 28.580 ;
        RECT 34.890 28.400 35.200 28.580 ;
        RECT 35.370 28.400 35.680 28.580 ;
        RECT 35.850 28.400 36.160 28.580 ;
        RECT 36.330 28.400 36.640 28.580 ;
        RECT 36.810 28.400 37.120 28.580 ;
        RECT 37.290 28.400 37.600 28.580 ;
        RECT 37.770 28.400 38.080 28.580 ;
        RECT 38.250 28.400 38.560 28.580 ;
        RECT 38.730 28.400 39.040 28.580 ;
        RECT 39.210 28.400 39.520 28.580 ;
        RECT 39.690 28.400 40.000 28.580 ;
        RECT 40.170 28.400 40.480 28.580 ;
        RECT 40.650 28.400 40.960 28.580 ;
        RECT 41.130 28.400 41.440 28.580 ;
        RECT 41.610 28.400 41.920 28.580 ;
        RECT 42.090 28.400 42.400 28.580 ;
        RECT 42.570 28.400 42.880 28.580 ;
        RECT 43.050 28.400 43.360 28.580 ;
        RECT 43.530 28.400 43.840 28.580 ;
        RECT 44.010 28.400 44.320 28.580 ;
        RECT 44.490 28.400 44.800 28.580 ;
        RECT 44.970 28.400 45.280 28.580 ;
        RECT 45.450 28.400 45.760 28.580 ;
        RECT 45.930 28.400 46.240 28.580 ;
        RECT 46.410 28.400 46.720 28.580 ;
        RECT 46.890 28.400 47.200 28.580 ;
        RECT 47.370 28.400 47.680 28.580 ;
        RECT 47.850 28.400 48.160 28.580 ;
        RECT 48.330 28.400 48.640 28.580 ;
        RECT 48.810 28.400 49.120 28.580 ;
        RECT 49.290 28.400 49.600 28.580 ;
        RECT 49.770 28.400 50.080 28.580 ;
        RECT 50.250 28.400 50.560 28.580 ;
        RECT 50.730 28.400 51.040 28.580 ;
        RECT 51.210 28.400 51.520 28.580 ;
        RECT 51.690 28.400 52.000 28.580 ;
        RECT 52.170 28.400 52.480 28.580 ;
        RECT 52.650 28.400 52.960 28.580 ;
        RECT 53.130 28.400 53.440 28.580 ;
        RECT 53.610 28.400 53.920 28.580 ;
        RECT 54.090 28.400 54.400 28.580 ;
        RECT 54.570 28.400 54.880 28.580 ;
        RECT 55.050 28.400 55.360 28.580 ;
        RECT 55.530 28.400 55.840 28.580 ;
        RECT 56.010 28.400 56.320 28.580 ;
        RECT 56.490 28.400 56.800 28.580 ;
        RECT 56.970 28.400 57.280 28.580 ;
        RECT 57.450 28.400 57.760 28.580 ;
        RECT 57.930 28.400 58.240 28.580 ;
        RECT 58.410 28.400 58.720 28.580 ;
        RECT 58.890 28.400 59.200 28.580 ;
        RECT 59.370 28.400 59.680 28.580 ;
        RECT 59.850 28.400 60.160 28.580 ;
        RECT 60.330 28.400 60.640 28.580 ;
        RECT 60.810 28.400 61.120 28.580 ;
        RECT 61.290 28.400 61.600 28.580 ;
        RECT 61.770 28.400 62.080 28.580 ;
        RECT 62.250 28.400 62.560 28.580 ;
        RECT 62.730 28.400 63.040 28.580 ;
        RECT 63.210 28.400 63.520 28.580 ;
        RECT 63.690 28.400 64.000 28.580 ;
        RECT 64.170 28.400 64.480 28.580 ;
        RECT 64.650 28.400 64.960 28.580 ;
        RECT 65.130 28.400 65.440 28.580 ;
        RECT 65.610 28.400 65.920 28.580 ;
        RECT 66.090 28.400 66.400 28.580 ;
        RECT 66.570 28.400 66.880 28.580 ;
        RECT 67.050 28.400 67.360 28.580 ;
        RECT 67.530 28.400 67.840 28.580 ;
        RECT 68.010 28.400 68.320 28.580 ;
        RECT 68.490 28.400 68.800 28.580 ;
        RECT 68.970 28.400 69.280 28.580 ;
        RECT 69.450 28.400 69.760 28.580 ;
        RECT 69.930 28.400 70.240 28.580 ;
        RECT 70.410 28.400 70.720 28.580 ;
        RECT 70.890 28.400 71.200 28.580 ;
        RECT 71.370 28.400 71.680 28.580 ;
        RECT 71.850 28.400 72.160 28.580 ;
        RECT 72.330 28.400 72.640 28.580 ;
        RECT 72.810 28.400 73.120 28.580 ;
        RECT 73.290 28.400 73.600 28.580 ;
        RECT 73.770 28.400 74.080 28.580 ;
        RECT 74.250 28.400 74.560 28.580 ;
        RECT 74.730 28.400 75.040 28.580 ;
        RECT 75.210 28.400 75.520 28.580 ;
        RECT 75.690 28.400 76.000 28.580 ;
        RECT 76.170 28.400 76.480 28.580 ;
        RECT 76.650 28.400 76.960 28.580 ;
        RECT 77.130 28.400 77.440 28.580 ;
        RECT 77.610 28.400 77.920 28.580 ;
        RECT 78.090 28.400 78.400 28.580 ;
        RECT 78.570 28.400 78.880 28.580 ;
        RECT 79.050 28.400 79.360 28.580 ;
        RECT 79.530 28.400 79.840 28.580 ;
        RECT 80.010 28.400 80.320 28.580 ;
        RECT 80.490 28.400 80.800 28.580 ;
        RECT 80.970 28.400 81.280 28.580 ;
        RECT 81.450 28.400 81.760 28.580 ;
        RECT 81.930 28.400 82.240 28.580 ;
        RECT 82.410 28.400 82.720 28.580 ;
        RECT 82.890 28.400 83.200 28.580 ;
        RECT 83.370 28.400 83.680 28.580 ;
        RECT 83.850 28.400 84.160 28.580 ;
        RECT 84.330 28.400 84.640 28.580 ;
        RECT 84.810 28.400 85.120 28.580 ;
        RECT 85.290 28.400 85.600 28.580 ;
        RECT 85.770 28.400 86.080 28.580 ;
        RECT 86.250 28.400 86.560 28.580 ;
        RECT 86.730 28.400 87.040 28.580 ;
        RECT 87.210 28.400 87.520 28.580 ;
        RECT 87.690 28.400 88.000 28.580 ;
        RECT 88.170 28.400 88.480 28.580 ;
        RECT 88.650 28.400 88.960 28.580 ;
        RECT 89.130 28.400 89.440 28.580 ;
        RECT 89.610 28.400 89.920 28.580 ;
        RECT 90.090 28.400 90.400 28.580 ;
        RECT 90.570 28.400 90.880 28.580 ;
        RECT 91.050 28.400 91.360 28.580 ;
        RECT 91.530 28.400 91.840 28.580 ;
        RECT 92.010 28.400 92.320 28.580 ;
        RECT 92.490 28.400 92.800 28.580 ;
        RECT 92.970 28.400 93.280 28.580 ;
        RECT 93.450 28.400 93.760 28.580 ;
        RECT 93.930 28.400 94.240 28.580 ;
        RECT 94.410 28.400 94.720 28.580 ;
        RECT 94.890 28.400 95.200 28.580 ;
        RECT 95.370 28.400 95.680 28.580 ;
        RECT 95.850 28.400 96.160 28.580 ;
        RECT 96.330 28.400 96.640 28.580 ;
        RECT 96.810 28.400 97.120 28.580 ;
        RECT 97.290 28.400 97.600 28.580 ;
        RECT 97.770 28.400 98.080 28.580 ;
        RECT 98.250 28.400 98.560 28.580 ;
        RECT 98.730 28.400 99.040 28.580 ;
        RECT 99.210 28.400 99.520 28.580 ;
        RECT 99.690 28.400 100.000 28.580 ;
        RECT 100.170 28.400 100.480 28.580 ;
        RECT 100.650 28.400 100.960 28.580 ;
        RECT 101.130 28.400 101.440 28.580 ;
        RECT 101.610 28.400 101.920 28.580 ;
        RECT 102.090 28.400 102.400 28.580 ;
        RECT 102.570 28.400 102.880 28.580 ;
        RECT 103.050 28.400 103.360 28.580 ;
        RECT 103.530 28.400 103.840 28.580 ;
        RECT 104.010 28.400 104.160 28.580 ;
        RECT 104.640 28.400 104.800 28.580 ;
        RECT 104.970 28.400 105.280 28.580 ;
        RECT 105.450 28.400 105.760 28.580 ;
        RECT 105.930 28.400 106.240 28.580 ;
        RECT 106.410 28.400 106.720 28.580 ;
        RECT 106.890 28.400 107.200 28.580 ;
        RECT 107.370 28.400 107.680 28.580 ;
        RECT 107.850 28.400 108.160 28.580 ;
        RECT 108.330 28.400 108.640 28.580 ;
        RECT 108.810 28.400 109.120 28.580 ;
        RECT 109.290 28.400 109.600 28.580 ;
        RECT 109.770 28.400 110.080 28.580 ;
        RECT 110.250 28.400 110.560 28.580 ;
        RECT 110.730 28.400 111.040 28.580 ;
        RECT 111.210 28.400 111.520 28.580 ;
        RECT 111.690 28.400 112.000 28.580 ;
        RECT 112.170 28.400 112.480 28.580 ;
        RECT 112.650 28.400 112.960 28.580 ;
        RECT 113.130 28.400 113.440 28.580 ;
        RECT 113.610 28.400 113.920 28.580 ;
        RECT 114.090 28.400 114.400 28.580 ;
        RECT 114.570 28.400 114.880 28.580 ;
        RECT 115.050 28.400 115.360 28.580 ;
        RECT 115.530 28.400 115.840 28.580 ;
        RECT 116.010 28.400 116.320 28.580 ;
        RECT 116.490 28.400 116.800 28.580 ;
        RECT 116.970 28.400 117.280 28.580 ;
        RECT 117.450 28.400 117.760 28.580 ;
        RECT 117.930 28.400 118.240 28.580 ;
        RECT 118.410 28.400 118.720 28.580 ;
        RECT 118.890 28.400 119.200 28.580 ;
        RECT 119.370 28.400 119.520 28.580 ;
        RECT 120.000 28.400 120.160 28.580 ;
        RECT 120.330 28.400 120.640 28.580 ;
        RECT 120.810 28.400 121.120 28.580 ;
        RECT 121.290 28.400 121.600 28.580 ;
        RECT 121.770 28.400 122.080 28.580 ;
        RECT 122.250 28.400 122.560 28.580 ;
        RECT 122.730 28.400 123.040 28.580 ;
        RECT 123.210 28.400 123.520 28.580 ;
        RECT 123.690 28.400 124.000 28.580 ;
        RECT 124.170 28.400 124.480 28.580 ;
        RECT 124.650 28.400 124.960 28.580 ;
        RECT 125.130 28.400 125.440 28.580 ;
        RECT 125.610 28.400 125.920 28.580 ;
        RECT 126.090 28.400 126.400 28.580 ;
        RECT 126.570 28.400 126.880 28.580 ;
        RECT 127.050 28.400 127.360 28.580 ;
        RECT 127.530 28.400 127.840 28.580 ;
        RECT 128.010 28.400 128.320 28.580 ;
        RECT 128.490 28.400 128.800 28.580 ;
        RECT 128.970 28.400 129.280 28.580 ;
        RECT 129.450 28.400 129.760 28.580 ;
        RECT 129.930 28.400 130.240 28.580 ;
        RECT 130.410 28.400 130.720 28.580 ;
        RECT 130.890 28.400 131.200 28.580 ;
        RECT 131.370 28.400 131.680 28.580 ;
        RECT 131.850 28.400 132.000 28.580 ;
        RECT 132.480 28.400 132.640 28.580 ;
        RECT 132.810 28.400 133.120 28.580 ;
        RECT 133.290 28.400 133.600 28.580 ;
        RECT 133.770 28.400 134.080 28.580 ;
        RECT 134.250 28.400 134.560 28.580 ;
        RECT 134.730 28.400 135.040 28.580 ;
        RECT 135.210 28.400 135.520 28.580 ;
        RECT 135.690 28.400 136.000 28.580 ;
        RECT 136.170 28.400 136.480 28.580 ;
        RECT 136.650 28.400 136.960 28.580 ;
        RECT 137.130 28.400 137.440 28.580 ;
        RECT 137.610 28.400 137.920 28.580 ;
        RECT 138.090 28.400 138.400 28.580 ;
        RECT 138.570 28.400 138.880 28.580 ;
        RECT 139.050 28.400 139.360 28.580 ;
        RECT 139.530 28.400 139.840 28.580 ;
        RECT 140.010 28.400 140.320 28.580 ;
        RECT 140.490 28.400 140.800 28.580 ;
        RECT 140.970 28.400 141.280 28.580 ;
        RECT 141.450 28.400 141.600 28.580 ;
        RECT 6.340 28.100 9.070 28.130 ;
        RECT 6.340 27.930 6.510 28.100 ;
        RECT 6.680 27.930 6.950 28.100 ;
        RECT 7.120 27.930 7.360 28.100 ;
        RECT 7.530 27.930 7.790 28.100 ;
        RECT 7.960 27.930 8.230 28.100 ;
        RECT 8.400 27.930 8.640 28.100 ;
        RECT 8.810 27.930 9.070 28.100 ;
        RECT 6.340 27.130 9.070 27.930 ;
        RECT 10.180 28.100 12.910 28.130 ;
        RECT 10.180 27.930 10.350 28.100 ;
        RECT 10.520 27.930 10.790 28.100 ;
        RECT 10.960 27.930 11.200 28.100 ;
        RECT 11.370 27.930 11.630 28.100 ;
        RECT 11.800 27.930 12.070 28.100 ;
        RECT 12.240 27.930 12.480 28.100 ;
        RECT 12.650 27.930 12.910 28.100 ;
        RECT 10.180 27.130 12.910 27.930 ;
        RECT 14.970 28.090 15.560 28.120 ;
        RECT 14.970 27.920 15.000 28.090 ;
        RECT 15.170 27.920 15.360 28.090 ;
        RECT 15.530 27.920 15.560 28.090 ;
        RECT 16.490 28.090 18.100 28.120 ;
        RECT 14.970 27.160 15.560 27.920 ;
        RECT 6.500 26.460 6.830 27.130 ;
        RECT 7.230 25.810 7.560 26.790 ;
        RECT 7.780 26.460 8.110 27.130 ;
        RECT 8.510 25.810 8.840 26.790 ;
        RECT 10.340 26.460 10.670 27.130 ;
        RECT 11.070 25.810 11.400 26.790 ;
        RECT 11.620 26.460 11.950 27.130 ;
        RECT 12.350 25.810 12.680 26.790 ;
      LAYER li1 ;
        RECT 15.010 26.550 15.720 26.940 ;
        RECT 15.900 26.310 16.230 27.990 ;
      LAYER li1 ;
        RECT 16.490 27.920 16.540 28.090 ;
        RECT 16.710 27.920 16.980 28.090 ;
        RECT 17.150 27.920 17.420 28.090 ;
        RECT 17.590 27.920 17.830 28.090 ;
        RECT 18.000 27.920 18.100 28.090 ;
        RECT 16.490 27.640 18.100 27.920 ;
        RECT 16.800 27.240 18.100 27.640 ;
        RECT 18.330 28.090 19.260 28.120 ;
        RECT 18.330 27.920 18.350 28.090 ;
        RECT 18.520 27.920 18.710 28.090 ;
        RECT 18.880 27.920 19.070 28.090 ;
        RECT 19.240 27.920 19.260 28.090 ;
        RECT 19.960 28.090 20.550 28.120 ;
        RECT 16.800 26.460 17.130 27.240 ;
        RECT 18.330 27.160 19.260 27.920 ;
      LAYER li1 ;
        RECT 19.440 27.060 19.770 27.990 ;
      LAYER li1 ;
        RECT 19.960 27.920 19.990 28.090 ;
        RECT 20.160 27.920 20.350 28.090 ;
        RECT 20.520 27.920 20.550 28.090 ;
        RECT 19.960 27.240 20.550 27.920 ;
        RECT 20.810 28.090 22.420 28.120 ;
        RECT 23.110 28.090 24.360 28.120 ;
        RECT 25.130 28.090 26.740 28.120 ;
        RECT 20.810 27.920 20.860 28.090 ;
        RECT 21.030 27.920 21.300 28.090 ;
        RECT 21.470 27.920 21.740 28.090 ;
        RECT 21.910 27.920 22.150 28.090 ;
        RECT 22.320 27.920 22.420 28.090 ;
        RECT 20.810 27.640 22.420 27.920 ;
        RECT 21.120 27.240 22.420 27.640 ;
      LAYER li1 ;
        RECT 19.440 26.890 20.520 27.060 ;
      LAYER li1 ;
        RECT 6.260 24.930 9.000 25.810 ;
        RECT 6.260 24.760 6.470 24.930 ;
        RECT 6.640 24.760 6.910 24.930 ;
        RECT 7.080 24.760 7.320 24.930 ;
        RECT 7.490 24.760 7.750 24.930 ;
        RECT 7.920 24.760 8.190 24.930 ;
        RECT 8.360 24.760 8.600 24.930 ;
        RECT 8.770 24.760 9.000 24.930 ;
        RECT 6.260 24.740 9.000 24.760 ;
        RECT 10.100 24.930 12.840 25.810 ;
        RECT 10.100 24.760 10.310 24.930 ;
        RECT 10.480 24.760 10.750 24.930 ;
        RECT 10.920 24.760 11.160 24.930 ;
        RECT 11.330 24.760 11.590 24.930 ;
        RECT 11.760 24.760 12.030 24.930 ;
        RECT 12.200 24.760 12.440 24.930 ;
        RECT 12.610 24.760 12.840 24.930 ;
        RECT 10.100 24.740 12.840 24.760 ;
        RECT 14.970 24.980 15.560 26.310 ;
        RECT 14.970 24.810 15.000 24.980 ;
        RECT 15.170 24.810 15.360 24.980 ;
        RECT 15.530 24.810 15.560 24.980 ;
        RECT 14.970 24.730 15.560 24.810 ;
      LAYER li1 ;
        RECT 15.840 24.730 16.230 26.310 ;
      LAYER li1 ;
        RECT 17.340 25.800 17.670 26.790 ;
      LAYER li1 ;
        RECT 18.370 26.370 19.560 26.710 ;
        RECT 19.740 26.370 20.070 26.710 ;
      LAYER li1 ;
        RECT 16.570 24.930 18.020 25.800 ;
        RECT 16.570 24.760 16.820 24.930 ;
        RECT 16.990 24.760 17.180 24.930 ;
        RECT 17.350 24.760 17.620 24.930 ;
        RECT 17.790 24.760 18.020 24.930 ;
        RECT 16.570 24.730 18.020 24.760 ;
        RECT 18.330 24.980 20.000 26.190 ;
        RECT 18.330 24.810 18.360 24.980 ;
        RECT 18.530 24.810 18.720 24.980 ;
        RECT 18.890 24.810 19.080 24.980 ;
        RECT 19.250 24.810 19.440 24.980 ;
        RECT 19.610 24.810 19.800 24.980 ;
        RECT 19.970 24.810 20.000 24.980 ;
        RECT 18.330 24.730 20.000 24.810 ;
      LAYER li1 ;
        RECT 20.260 24.730 20.520 26.890 ;
      LAYER li1 ;
        RECT 21.120 26.460 21.450 27.240 ;
        RECT 21.660 25.800 21.990 26.790 ;
      LAYER li1 ;
        RECT 22.680 26.310 22.930 27.990 ;
      LAYER li1 ;
        RECT 23.280 27.920 23.470 28.090 ;
        RECT 23.640 27.920 23.830 28.090 ;
        RECT 24.000 27.920 24.190 28.090 ;
        RECT 23.110 27.550 24.360 27.920 ;
        RECT 24.540 27.370 24.790 27.990 ;
        RECT 25.130 27.920 25.180 28.090 ;
        RECT 25.350 27.920 25.620 28.090 ;
        RECT 25.790 27.920 26.060 28.090 ;
        RECT 26.230 27.920 26.470 28.090 ;
        RECT 26.640 27.920 26.740 28.090 ;
        RECT 25.130 27.640 26.740 27.920 ;
        RECT 23.240 27.200 24.790 27.370 ;
        RECT 23.240 26.740 23.570 27.200 ;
        RECT 20.890 24.930 22.340 25.800 ;
        RECT 20.890 24.760 21.140 24.930 ;
        RECT 21.310 24.760 21.500 24.930 ;
        RECT 21.670 24.760 21.940 24.930 ;
        RECT 22.110 24.760 22.340 24.930 ;
        RECT 20.890 24.730 22.340 24.760 ;
      LAYER li1 ;
        RECT 22.680 24.730 23.110 26.310 ;
      LAYER li1 ;
        RECT 23.290 24.980 23.850 26.310 ;
      LAYER li1 ;
        RECT 24.030 25.230 24.360 27.020 ;
      LAYER li1 ;
        RECT 24.540 25.480 24.790 27.200 ;
        RECT 25.440 27.240 26.740 27.640 ;
        RECT 26.970 28.090 27.900 28.120 ;
        RECT 26.970 27.920 26.990 28.090 ;
        RECT 27.160 27.920 27.350 28.090 ;
        RECT 27.520 27.920 27.710 28.090 ;
        RECT 27.880 27.920 27.900 28.090 ;
        RECT 28.600 28.090 29.190 28.120 ;
        RECT 25.440 26.460 25.770 27.240 ;
        RECT 26.970 27.160 27.900 27.920 ;
      LAYER li1 ;
        RECT 28.080 27.060 28.410 27.990 ;
      LAYER li1 ;
        RECT 28.600 27.920 28.630 28.090 ;
        RECT 28.800 27.920 28.990 28.090 ;
        RECT 29.160 27.920 29.190 28.090 ;
        RECT 28.600 27.240 29.190 27.920 ;
        RECT 29.450 28.090 31.060 28.120 ;
        RECT 29.450 27.920 29.500 28.090 ;
        RECT 29.670 27.920 29.940 28.090 ;
        RECT 30.110 27.920 30.380 28.090 ;
        RECT 30.550 27.920 30.790 28.090 ;
        RECT 30.960 27.920 31.060 28.090 ;
        RECT 29.450 27.640 31.060 27.920 ;
        RECT 29.760 27.240 31.060 27.640 ;
        RECT 31.290 28.090 32.910 28.120 ;
        RECT 35.140 28.100 37.870 28.130 ;
        RECT 31.290 27.920 31.300 28.090 ;
        RECT 31.470 27.920 31.660 28.090 ;
        RECT 31.830 27.920 32.020 28.090 ;
        RECT 32.190 27.920 32.380 28.090 ;
        RECT 32.550 27.920 32.740 28.090 ;
      LAYER li1 ;
        RECT 28.080 26.890 29.160 27.060 ;
      LAYER li1 ;
        RECT 25.980 25.800 26.310 26.790 ;
      LAYER li1 ;
        RECT 27.010 26.370 28.200 26.710 ;
        RECT 28.380 26.370 28.710 26.710 ;
      LAYER li1 ;
        RECT 23.290 24.810 23.300 24.980 ;
        RECT 23.470 24.810 23.660 24.980 ;
        RECT 23.830 24.810 23.850 24.980 ;
        RECT 23.290 24.730 23.850 24.810 ;
        RECT 25.210 24.930 26.660 25.800 ;
        RECT 25.210 24.760 25.460 24.930 ;
        RECT 25.630 24.760 25.820 24.930 ;
        RECT 25.990 24.760 26.260 24.930 ;
        RECT 26.430 24.760 26.660 24.930 ;
        RECT 25.210 24.730 26.660 24.760 ;
        RECT 26.970 24.980 28.640 26.190 ;
        RECT 26.970 24.810 27.000 24.980 ;
        RECT 27.170 24.810 27.360 24.980 ;
        RECT 27.530 24.810 27.720 24.980 ;
        RECT 27.890 24.810 28.080 24.980 ;
        RECT 28.250 24.810 28.440 24.980 ;
        RECT 28.610 24.810 28.640 24.980 ;
        RECT 26.970 24.730 28.640 24.810 ;
      LAYER li1 ;
        RECT 28.900 24.730 29.160 26.890 ;
      LAYER li1 ;
        RECT 29.760 26.460 30.090 27.240 ;
        RECT 31.290 27.160 32.910 27.920 ;
        RECT 30.300 25.800 30.630 26.790 ;
      LAYER li1 ;
        RECT 31.330 26.650 32.200 26.980 ;
        RECT 33.090 26.760 33.480 27.680 ;
        RECT 33.660 26.760 33.930 27.680 ;
        RECT 34.110 27.160 34.440 27.990 ;
        RECT 34.180 26.580 34.440 27.160 ;
      LAYER li1 ;
        RECT 35.140 27.930 35.310 28.100 ;
        RECT 35.480 27.930 35.750 28.100 ;
        RECT 35.920 27.930 36.160 28.100 ;
        RECT 36.330 27.930 36.590 28.100 ;
        RECT 36.760 27.930 37.030 28.100 ;
        RECT 37.200 27.930 37.440 28.100 ;
        RECT 37.610 27.930 37.870 28.100 ;
        RECT 35.140 27.130 37.870 27.930 ;
        RECT 39.450 28.090 40.040 28.120 ;
        RECT 39.450 27.920 39.480 28.090 ;
        RECT 39.650 27.920 39.840 28.090 ;
        RECT 40.010 27.920 40.040 28.090 ;
        RECT 40.720 28.090 41.670 28.120 ;
        RECT 39.450 27.160 40.040 27.920 ;
      LAYER li1 ;
        RECT 32.400 26.410 34.440 26.580 ;
      LAYER li1 ;
        RECT 35.300 26.460 35.630 27.130 ;
        RECT 29.530 24.930 30.980 25.800 ;
        RECT 29.530 24.760 29.780 24.930 ;
        RECT 29.950 24.760 30.140 24.930 ;
        RECT 30.310 24.760 30.580 24.930 ;
        RECT 30.750 24.760 30.980 24.930 ;
        RECT 29.530 24.730 30.980 24.760 ;
        RECT 31.290 24.980 32.220 26.310 ;
        RECT 31.290 24.810 31.310 24.980 ;
        RECT 31.480 24.810 31.670 24.980 ;
        RECT 31.840 24.810 32.030 24.980 ;
        RECT 32.200 24.810 32.220 24.980 ;
        RECT 31.290 24.730 32.220 24.810 ;
      LAYER li1 ;
        RECT 32.400 24.730 32.570 26.410 ;
      LAYER li1 ;
        RECT 32.750 24.980 34.000 26.230 ;
        RECT 32.920 24.810 33.110 24.980 ;
        RECT 33.280 24.810 33.470 24.980 ;
        RECT 33.640 24.810 33.830 24.980 ;
        RECT 32.750 24.730 34.000 24.810 ;
      LAYER li1 ;
        RECT 34.180 24.730 34.440 26.410 ;
      LAYER li1 ;
        RECT 36.030 25.810 36.360 26.790 ;
        RECT 36.580 26.460 36.910 27.130 ;
      LAYER li1 ;
        RECT 40.290 27.060 40.540 27.990 ;
      LAYER li1 ;
        RECT 40.720 27.920 40.750 28.090 ;
        RECT 40.920 27.920 41.110 28.090 ;
        RECT 41.280 27.920 41.470 28.090 ;
        RECT 41.640 27.920 41.670 28.090 ;
        RECT 42.890 28.090 44.500 28.120 ;
        RECT 40.720 27.240 41.670 27.920 ;
      LAYER li1 ;
        RECT 41.850 27.060 42.120 27.990 ;
      LAYER li1 ;
        RECT 42.890 27.920 42.940 28.090 ;
        RECT 43.110 27.920 43.380 28.090 ;
        RECT 43.550 27.920 43.820 28.090 ;
        RECT 43.990 27.920 44.230 28.090 ;
        RECT 44.400 27.920 44.500 28.090 ;
        RECT 45.170 28.090 46.030 28.120 ;
        RECT 42.890 27.640 44.500 27.920 ;
        RECT 37.310 25.810 37.640 26.790 ;
        RECT 35.060 24.930 37.800 25.810 ;
      LAYER li1 ;
        RECT 38.070 25.260 38.240 26.910 ;
        RECT 39.490 26.370 39.790 26.960 ;
        RECT 40.290 26.890 42.120 27.060 ;
        RECT 39.970 26.370 41.160 26.710 ;
      LAYER li1 ;
        RECT 35.060 24.760 35.270 24.930 ;
        RECT 35.440 24.760 35.710 24.930 ;
        RECT 35.880 24.760 36.120 24.930 ;
        RECT 36.290 24.760 36.550 24.930 ;
        RECT 36.720 24.760 36.990 24.930 ;
        RECT 37.160 24.760 37.400 24.930 ;
        RECT 37.570 24.760 37.800 24.930 ;
        RECT 35.060 24.740 37.800 24.760 ;
        RECT 39.450 24.980 41.120 26.190 ;
      LAYER li1 ;
        RECT 41.340 25.230 41.670 26.710 ;
      LAYER li1 ;
        RECT 39.450 24.810 39.480 24.980 ;
        RECT 39.650 24.810 39.840 24.980 ;
        RECT 40.010 24.810 40.200 24.980 ;
        RECT 40.370 24.810 40.560 24.980 ;
        RECT 40.730 24.810 40.920 24.980 ;
        RECT 41.090 24.810 41.120 24.980 ;
        RECT 39.450 24.730 41.120 24.810 ;
      LAYER li1 ;
        RECT 41.850 24.730 42.120 26.890 ;
      LAYER li1 ;
        RECT 43.200 27.240 44.500 27.640 ;
        RECT 43.200 26.460 43.530 27.240 ;
        RECT 44.790 26.930 45.000 27.990 ;
        RECT 45.170 27.920 45.220 28.090 ;
        RECT 45.390 27.920 45.810 28.090 ;
        RECT 45.980 27.920 46.030 28.090 ;
        RECT 47.260 28.090 47.930 28.120 ;
        RECT 45.170 27.580 46.030 27.920 ;
        RECT 46.210 27.580 46.610 27.990 ;
        RECT 47.260 27.920 47.330 28.090 ;
        RECT 47.500 27.920 47.690 28.090 ;
        RECT 47.860 27.920 47.930 28.090 ;
        RECT 49.060 28.100 51.790 28.130 ;
      LAYER li1 ;
        RECT 45.170 27.100 45.960 27.410 ;
      LAYER li1 ;
        RECT 46.210 26.930 46.380 27.580 ;
      LAYER li1 ;
        RECT 46.560 27.100 47.090 27.410 ;
      LAYER li1 ;
        RECT 47.260 27.160 47.930 27.920 ;
        RECT 43.740 25.800 44.070 26.790 ;
        RECT 44.790 26.760 47.900 26.930 ;
        RECT 42.970 24.930 44.420 25.800 ;
        RECT 44.790 25.710 45.040 26.760 ;
      LAYER li1 ;
        RECT 45.250 25.230 46.180 26.580 ;
      LAYER li1 ;
        RECT 47.570 26.550 47.900 26.760 ;
        RECT 46.350 25.060 47.920 26.310 ;
        RECT 42.970 24.760 43.220 24.930 ;
        RECT 43.390 24.760 43.580 24.930 ;
        RECT 43.750 24.760 44.020 24.930 ;
        RECT 44.190 24.760 44.420 24.930 ;
        RECT 42.970 24.730 44.420 24.760 ;
        RECT 46.260 24.980 47.920 25.060 ;
        RECT 46.260 24.810 46.310 24.980 ;
        RECT 46.480 24.810 46.670 24.980 ;
        RECT 46.840 24.810 47.030 24.980 ;
        RECT 47.200 24.810 47.390 24.980 ;
        RECT 47.560 24.810 47.750 24.980 ;
        RECT 46.260 24.730 47.920 24.810 ;
      LAYER li1 ;
        RECT 48.100 24.730 48.360 27.990 ;
      LAYER li1 ;
        RECT 49.060 27.930 49.230 28.100 ;
        RECT 49.400 27.930 49.670 28.100 ;
        RECT 49.840 27.930 50.080 28.100 ;
        RECT 50.250 27.930 50.510 28.100 ;
        RECT 50.680 27.930 50.950 28.100 ;
        RECT 51.120 27.930 51.360 28.100 ;
        RECT 51.530 27.930 51.790 28.100 ;
        RECT 49.060 27.130 51.790 27.930 ;
        RECT 52.890 28.090 53.840 28.120 ;
        RECT 52.890 27.920 52.920 28.090 ;
        RECT 53.090 27.920 53.280 28.090 ;
        RECT 53.450 27.920 53.640 28.090 ;
        RECT 53.810 27.920 53.840 28.090 ;
        RECT 54.450 28.090 55.400 28.120 ;
        RECT 52.890 27.160 53.840 27.920 ;
      LAYER li1 ;
        RECT 54.020 27.280 54.270 27.990 ;
      LAYER li1 ;
        RECT 54.450 27.920 54.480 28.090 ;
        RECT 54.650 27.920 54.840 28.090 ;
        RECT 55.010 27.920 55.200 28.090 ;
        RECT 55.370 27.920 55.400 28.090 ;
        RECT 56.010 28.090 56.960 28.120 ;
        RECT 54.450 27.460 55.400 27.920 ;
      LAYER li1 ;
        RECT 55.580 27.280 55.830 27.990 ;
      LAYER li1 ;
        RECT 49.220 26.460 49.550 27.130 ;
        RECT 49.950 25.810 50.280 26.790 ;
        RECT 50.500 26.460 50.830 27.130 ;
      LAYER li1 ;
        RECT 54.020 27.110 55.830 27.280 ;
      LAYER li1 ;
        RECT 56.010 27.920 56.040 28.090 ;
        RECT 56.210 27.920 56.400 28.090 ;
        RECT 56.570 27.920 56.760 28.090 ;
        RECT 56.930 27.920 56.960 28.090 ;
        RECT 57.770 28.090 59.380 28.120 ;
        RECT 56.010 27.240 56.960 27.920 ;
      LAYER li1 ;
        RECT 54.020 26.940 54.190 27.110 ;
      LAYER li1 ;
        RECT 57.140 27.060 57.470 27.990 ;
        RECT 57.770 27.920 57.820 28.090 ;
        RECT 57.990 27.920 58.260 28.090 ;
        RECT 58.430 27.920 58.700 28.090 ;
        RECT 58.870 27.920 59.110 28.090 ;
        RECT 59.280 27.920 59.380 28.090 ;
        RECT 57.770 27.640 59.380 27.920 ;
        RECT 51.230 25.810 51.560 26.790 ;
      LAYER li1 ;
        RECT 52.930 26.710 54.190 26.940 ;
      LAYER li1 ;
        RECT 56.230 26.930 57.470 27.060 ;
        RECT 54.370 26.890 57.470 26.930 ;
        RECT 54.370 26.760 56.400 26.890 ;
      LAYER li1 ;
        RECT 54.020 26.580 54.190 26.710 ;
        RECT 54.020 26.410 55.910 26.580 ;
      LAYER li1 ;
        RECT 48.980 24.930 51.720 25.810 ;
        RECT 48.980 24.760 49.190 24.930 ;
        RECT 49.360 24.760 49.630 24.930 ;
        RECT 49.800 24.760 50.040 24.930 ;
        RECT 50.210 24.760 50.470 24.930 ;
        RECT 50.640 24.760 50.910 24.930 ;
        RECT 51.080 24.760 51.320 24.930 ;
        RECT 51.490 24.760 51.720 24.930 ;
        RECT 48.980 24.740 51.720 24.760 ;
        RECT 52.890 24.980 53.840 26.310 ;
        RECT 52.890 24.810 52.920 24.980 ;
        RECT 53.090 24.810 53.280 24.980 ;
        RECT 53.450 24.810 53.640 24.980 ;
        RECT 53.810 24.810 53.840 24.980 ;
        RECT 52.890 24.730 53.840 24.810 ;
      LAYER li1 ;
        RECT 54.020 24.730 54.270 26.410 ;
      LAYER li1 ;
        RECT 54.450 24.980 55.400 26.230 ;
        RECT 54.450 24.810 54.480 24.980 ;
        RECT 54.650 24.810 54.840 24.980 ;
        RECT 55.010 24.810 55.200 24.980 ;
        RECT 55.370 24.810 55.400 24.980 ;
        RECT 54.450 24.730 55.400 24.810 ;
      LAYER li1 ;
        RECT 55.580 24.730 55.910 26.410 ;
        RECT 56.690 26.370 57.020 26.710 ;
      LAYER li1 ;
        RECT 56.090 24.980 57.040 26.190 ;
        RECT 56.090 24.810 56.120 24.980 ;
        RECT 56.290 24.810 56.480 24.980 ;
        RECT 56.650 24.810 56.840 24.980 ;
        RECT 57.010 24.810 57.040 24.980 ;
        RECT 56.090 24.730 57.040 24.810 ;
        RECT 57.220 24.730 57.470 26.890 ;
        RECT 58.080 27.240 59.380 27.640 ;
        RECT 59.610 28.090 60.560 28.120 ;
        RECT 59.610 27.920 59.640 28.090 ;
        RECT 59.810 27.920 60.000 28.090 ;
        RECT 60.170 27.920 60.360 28.090 ;
        RECT 60.530 27.920 60.560 28.090 ;
        RECT 61.170 28.090 62.120 28.120 ;
        RECT 58.080 26.460 58.410 27.240 ;
        RECT 59.610 27.160 60.560 27.920 ;
      LAYER li1 ;
        RECT 60.740 27.280 60.990 27.990 ;
      LAYER li1 ;
        RECT 61.170 27.920 61.200 28.090 ;
        RECT 61.370 27.920 61.560 28.090 ;
        RECT 61.730 27.920 61.920 28.090 ;
        RECT 62.090 27.920 62.120 28.090 ;
        RECT 62.730 28.090 63.680 28.120 ;
        RECT 61.170 27.460 62.120 27.920 ;
      LAYER li1 ;
        RECT 62.300 27.280 62.550 27.990 ;
        RECT 60.740 27.110 62.550 27.280 ;
      LAYER li1 ;
        RECT 62.730 27.920 62.760 28.090 ;
        RECT 62.930 27.920 63.120 28.090 ;
        RECT 63.290 27.920 63.480 28.090 ;
        RECT 63.650 27.920 63.680 28.090 ;
        RECT 64.490 28.090 66.100 28.120 ;
        RECT 62.730 27.240 63.680 27.920 ;
      LAYER li1 ;
        RECT 60.740 26.940 60.910 27.110 ;
      LAYER li1 ;
        RECT 63.860 27.060 64.190 27.990 ;
        RECT 64.490 27.920 64.540 28.090 ;
        RECT 64.710 27.920 64.980 28.090 ;
        RECT 65.150 27.920 65.420 28.090 ;
        RECT 65.590 27.920 65.830 28.090 ;
        RECT 66.000 27.920 66.100 28.090 ;
        RECT 64.490 27.640 66.100 27.920 ;
        RECT 58.620 25.800 58.950 26.790 ;
      LAYER li1 ;
        RECT 59.650 26.710 60.910 26.940 ;
      LAYER li1 ;
        RECT 62.950 26.930 64.190 27.060 ;
        RECT 61.090 26.890 64.190 26.930 ;
        RECT 61.090 26.760 63.120 26.890 ;
      LAYER li1 ;
        RECT 60.740 26.580 60.910 26.710 ;
        RECT 60.740 26.410 62.630 26.580 ;
      LAYER li1 ;
        RECT 57.850 24.930 59.300 25.800 ;
        RECT 57.850 24.760 58.100 24.930 ;
        RECT 58.270 24.760 58.460 24.930 ;
        RECT 58.630 24.760 58.900 24.930 ;
        RECT 59.070 24.760 59.300 24.930 ;
        RECT 57.850 24.730 59.300 24.760 ;
        RECT 59.610 24.980 60.560 26.310 ;
        RECT 59.610 24.810 59.640 24.980 ;
        RECT 59.810 24.810 60.000 24.980 ;
        RECT 60.170 24.810 60.360 24.980 ;
        RECT 60.530 24.810 60.560 24.980 ;
        RECT 59.610 24.730 60.560 24.810 ;
      LAYER li1 ;
        RECT 60.740 24.730 60.990 26.410 ;
      LAYER li1 ;
        RECT 61.170 24.980 62.120 26.230 ;
        RECT 61.170 24.810 61.200 24.980 ;
        RECT 61.370 24.810 61.560 24.980 ;
        RECT 61.730 24.810 61.920 24.980 ;
        RECT 62.090 24.810 62.120 24.980 ;
        RECT 61.170 24.730 62.120 24.810 ;
      LAYER li1 ;
        RECT 62.300 24.730 62.630 26.410 ;
        RECT 63.410 26.370 63.740 26.710 ;
      LAYER li1 ;
        RECT 62.810 24.980 63.760 26.190 ;
        RECT 62.810 24.810 62.840 24.980 ;
        RECT 63.010 24.810 63.200 24.980 ;
        RECT 63.370 24.810 63.560 24.980 ;
        RECT 63.730 24.810 63.760 24.980 ;
        RECT 62.810 24.730 63.760 24.810 ;
        RECT 63.940 24.730 64.190 26.890 ;
        RECT 64.800 27.240 66.100 27.640 ;
        RECT 66.330 28.090 67.280 28.120 ;
        RECT 66.330 27.920 66.360 28.090 ;
        RECT 66.530 27.920 66.720 28.090 ;
        RECT 66.890 27.920 67.080 28.090 ;
        RECT 67.250 27.920 67.280 28.090 ;
        RECT 67.890 28.090 68.840 28.120 ;
        RECT 64.800 26.460 65.130 27.240 ;
        RECT 66.330 27.160 67.280 27.920 ;
      LAYER li1 ;
        RECT 67.460 27.280 67.710 27.990 ;
      LAYER li1 ;
        RECT 67.890 27.920 67.920 28.090 ;
        RECT 68.090 27.920 68.280 28.090 ;
        RECT 68.450 27.920 68.640 28.090 ;
        RECT 68.810 27.920 68.840 28.090 ;
        RECT 69.450 28.090 70.400 28.120 ;
        RECT 67.890 27.460 68.840 27.920 ;
      LAYER li1 ;
        RECT 69.020 27.280 69.270 27.990 ;
        RECT 67.460 27.110 69.270 27.280 ;
      LAYER li1 ;
        RECT 69.450 27.920 69.480 28.090 ;
        RECT 69.650 27.920 69.840 28.090 ;
        RECT 70.010 27.920 70.200 28.090 ;
        RECT 70.370 27.920 70.400 28.090 ;
        RECT 71.210 28.090 72.820 28.120 ;
        RECT 69.450 27.240 70.400 27.920 ;
      LAYER li1 ;
        RECT 67.460 26.940 67.630 27.110 ;
      LAYER li1 ;
        RECT 70.580 27.060 70.910 27.990 ;
        RECT 71.210 27.920 71.260 28.090 ;
        RECT 71.430 27.920 71.700 28.090 ;
        RECT 71.870 27.920 72.140 28.090 ;
        RECT 72.310 27.920 72.550 28.090 ;
        RECT 72.720 27.920 72.820 28.090 ;
        RECT 71.210 27.640 72.820 27.920 ;
        RECT 65.340 25.800 65.670 26.790 ;
      LAYER li1 ;
        RECT 66.370 26.710 67.630 26.940 ;
      LAYER li1 ;
        RECT 69.670 26.930 70.910 27.060 ;
        RECT 67.810 26.890 70.910 26.930 ;
        RECT 67.810 26.760 69.840 26.890 ;
      LAYER li1 ;
        RECT 67.460 26.580 67.630 26.710 ;
        RECT 67.460 26.410 69.350 26.580 ;
      LAYER li1 ;
        RECT 64.570 24.930 66.020 25.800 ;
        RECT 64.570 24.760 64.820 24.930 ;
        RECT 64.990 24.760 65.180 24.930 ;
        RECT 65.350 24.760 65.620 24.930 ;
        RECT 65.790 24.760 66.020 24.930 ;
        RECT 64.570 24.730 66.020 24.760 ;
        RECT 66.330 24.980 67.280 26.310 ;
        RECT 66.330 24.810 66.360 24.980 ;
        RECT 66.530 24.810 66.720 24.980 ;
        RECT 66.890 24.810 67.080 24.980 ;
        RECT 67.250 24.810 67.280 24.980 ;
        RECT 66.330 24.730 67.280 24.810 ;
      LAYER li1 ;
        RECT 67.460 24.730 67.710 26.410 ;
      LAYER li1 ;
        RECT 67.890 24.980 68.840 26.230 ;
        RECT 67.890 24.810 67.920 24.980 ;
        RECT 68.090 24.810 68.280 24.980 ;
        RECT 68.450 24.810 68.640 24.980 ;
        RECT 68.810 24.810 68.840 24.980 ;
        RECT 67.890 24.730 68.840 24.810 ;
      LAYER li1 ;
        RECT 69.020 24.730 69.350 26.410 ;
        RECT 70.130 26.370 70.460 26.710 ;
      LAYER li1 ;
        RECT 69.530 24.980 70.480 26.190 ;
        RECT 69.530 24.810 69.560 24.980 ;
        RECT 69.730 24.810 69.920 24.980 ;
        RECT 70.090 24.810 70.280 24.980 ;
        RECT 70.450 24.810 70.480 24.980 ;
        RECT 69.530 24.730 70.480 24.810 ;
        RECT 70.660 24.730 70.910 26.890 ;
        RECT 71.520 27.240 72.820 27.640 ;
        RECT 73.050 28.090 74.000 28.120 ;
        RECT 73.050 27.920 73.080 28.090 ;
        RECT 73.250 27.920 73.440 28.090 ;
        RECT 73.610 27.920 73.800 28.090 ;
        RECT 73.970 27.920 74.000 28.090 ;
        RECT 74.610 28.090 75.560 28.120 ;
        RECT 71.520 26.460 71.850 27.240 ;
        RECT 73.050 27.160 74.000 27.920 ;
      LAYER li1 ;
        RECT 74.180 27.280 74.430 27.990 ;
      LAYER li1 ;
        RECT 74.610 27.920 74.640 28.090 ;
        RECT 74.810 27.920 75.000 28.090 ;
        RECT 75.170 27.920 75.360 28.090 ;
        RECT 75.530 27.920 75.560 28.090 ;
        RECT 76.170 28.090 77.120 28.120 ;
        RECT 74.610 27.460 75.560 27.920 ;
      LAYER li1 ;
        RECT 75.740 27.280 75.990 27.990 ;
        RECT 74.180 27.110 75.990 27.280 ;
      LAYER li1 ;
        RECT 76.170 27.920 76.200 28.090 ;
        RECT 76.370 27.920 76.560 28.090 ;
        RECT 76.730 27.920 76.920 28.090 ;
        RECT 77.090 27.920 77.120 28.090 ;
        RECT 78.340 28.100 81.070 28.130 ;
        RECT 76.170 27.240 77.120 27.920 ;
      LAYER li1 ;
        RECT 74.180 26.940 74.350 27.110 ;
      LAYER li1 ;
        RECT 77.300 27.060 77.630 27.990 ;
        RECT 78.340 27.930 78.510 28.100 ;
        RECT 78.680 27.930 78.950 28.100 ;
        RECT 79.120 27.930 79.360 28.100 ;
        RECT 79.530 27.930 79.790 28.100 ;
        RECT 79.960 27.930 80.230 28.100 ;
        RECT 80.400 27.930 80.640 28.100 ;
        RECT 80.810 27.930 81.070 28.100 ;
        RECT 82.630 28.090 83.880 28.120 ;
        RECT 85.060 28.100 87.790 28.130 ;
        RECT 78.340 27.130 81.070 27.930 ;
        RECT 72.060 25.800 72.390 26.790 ;
      LAYER li1 ;
        RECT 73.090 26.710 74.350 26.940 ;
      LAYER li1 ;
        RECT 76.390 26.930 77.630 27.060 ;
        RECT 74.530 26.890 77.630 26.930 ;
        RECT 74.530 26.760 76.560 26.890 ;
      LAYER li1 ;
        RECT 74.180 26.580 74.350 26.710 ;
        RECT 74.180 26.410 76.070 26.580 ;
      LAYER li1 ;
        RECT 71.290 24.930 72.740 25.800 ;
        RECT 71.290 24.760 71.540 24.930 ;
        RECT 71.710 24.760 71.900 24.930 ;
        RECT 72.070 24.760 72.340 24.930 ;
        RECT 72.510 24.760 72.740 24.930 ;
        RECT 71.290 24.730 72.740 24.760 ;
        RECT 73.050 24.980 74.000 26.310 ;
        RECT 73.050 24.810 73.080 24.980 ;
        RECT 73.250 24.810 73.440 24.980 ;
        RECT 73.610 24.810 73.800 24.980 ;
        RECT 73.970 24.810 74.000 24.980 ;
        RECT 73.050 24.730 74.000 24.810 ;
      LAYER li1 ;
        RECT 74.180 24.730 74.430 26.410 ;
      LAYER li1 ;
        RECT 74.610 24.980 75.560 26.230 ;
        RECT 74.610 24.810 74.640 24.980 ;
        RECT 74.810 24.810 75.000 24.980 ;
        RECT 75.170 24.810 75.360 24.980 ;
        RECT 75.530 24.810 75.560 24.980 ;
        RECT 74.610 24.730 75.560 24.810 ;
      LAYER li1 ;
        RECT 75.740 24.730 76.070 26.410 ;
        RECT 76.850 26.370 77.180 26.710 ;
      LAYER li1 ;
        RECT 76.250 24.980 77.200 26.190 ;
        RECT 76.250 24.810 76.280 24.980 ;
        RECT 76.450 24.810 76.640 24.980 ;
        RECT 76.810 24.810 77.000 24.980 ;
        RECT 77.170 24.810 77.200 24.980 ;
        RECT 76.250 24.730 77.200 24.810 ;
        RECT 77.380 24.730 77.630 26.890 ;
        RECT 78.500 26.460 78.830 27.130 ;
        RECT 79.230 25.810 79.560 26.790 ;
        RECT 79.780 26.460 80.110 27.130 ;
        RECT 80.510 25.810 80.840 26.790 ;
      LAYER li1 ;
        RECT 82.200 26.310 82.450 27.990 ;
      LAYER li1 ;
        RECT 82.800 27.920 82.990 28.090 ;
        RECT 83.160 27.920 83.350 28.090 ;
        RECT 83.520 27.920 83.710 28.090 ;
        RECT 82.630 27.550 83.880 27.920 ;
        RECT 84.060 27.370 84.310 27.990 ;
        RECT 82.760 27.200 84.310 27.370 ;
        RECT 82.760 26.740 83.090 27.200 ;
        RECT 78.260 24.930 81.000 25.810 ;
        RECT 78.260 24.760 78.470 24.930 ;
        RECT 78.640 24.760 78.910 24.930 ;
        RECT 79.080 24.760 79.320 24.930 ;
        RECT 79.490 24.760 79.750 24.930 ;
        RECT 79.920 24.760 80.190 24.930 ;
        RECT 80.360 24.760 80.600 24.930 ;
        RECT 80.770 24.760 81.000 24.930 ;
        RECT 78.260 24.740 81.000 24.760 ;
      LAYER li1 ;
        RECT 82.200 24.730 82.630 26.310 ;
      LAYER li1 ;
        RECT 82.810 24.980 83.370 26.310 ;
      LAYER li1 ;
        RECT 83.550 25.230 83.880 27.020 ;
      LAYER li1 ;
        RECT 84.060 25.480 84.310 27.200 ;
        RECT 85.060 27.930 85.230 28.100 ;
        RECT 85.400 27.930 85.670 28.100 ;
        RECT 85.840 27.930 86.080 28.100 ;
        RECT 86.250 27.930 86.510 28.100 ;
        RECT 86.680 27.930 86.950 28.100 ;
        RECT 87.120 27.930 87.360 28.100 ;
        RECT 87.530 27.930 87.790 28.100 ;
        RECT 85.060 27.130 87.790 27.930 ;
        RECT 88.890 28.090 89.820 28.120 ;
        RECT 88.890 27.920 88.910 28.090 ;
        RECT 89.080 27.920 89.270 28.090 ;
        RECT 89.440 27.920 89.630 28.090 ;
        RECT 89.800 27.920 89.820 28.090 ;
        RECT 90.520 28.090 91.110 28.120 ;
        RECT 88.890 27.160 89.820 27.920 ;
        RECT 85.220 26.460 85.550 27.130 ;
        RECT 85.950 25.810 86.280 26.790 ;
        RECT 86.500 26.460 86.830 27.130 ;
      LAYER li1 ;
        RECT 90.000 27.060 90.330 27.990 ;
      LAYER li1 ;
        RECT 90.520 27.920 90.550 28.090 ;
        RECT 90.720 27.920 90.910 28.090 ;
        RECT 91.080 27.920 91.110 28.090 ;
        RECT 90.520 27.240 91.110 27.920 ;
        RECT 91.370 28.090 92.980 28.120 ;
        RECT 91.370 27.920 91.420 28.090 ;
        RECT 91.590 27.920 91.860 28.090 ;
        RECT 92.030 27.920 92.300 28.090 ;
        RECT 92.470 27.920 92.710 28.090 ;
        RECT 92.880 27.920 92.980 28.090 ;
        RECT 91.370 27.640 92.980 27.920 ;
        RECT 91.680 27.240 92.980 27.640 ;
        RECT 94.650 28.090 95.960 28.120 ;
        RECT 94.650 27.920 94.680 28.090 ;
        RECT 94.850 27.920 95.040 28.090 ;
        RECT 95.210 27.920 95.400 28.090 ;
        RECT 95.570 27.920 95.760 28.090 ;
        RECT 95.930 27.920 95.960 28.090 ;
        RECT 97.130 28.090 98.740 28.120 ;
      LAYER li1 ;
        RECT 90.000 26.890 91.080 27.060 ;
      LAYER li1 ;
        RECT 87.230 25.810 87.560 26.790 ;
      LAYER li1 ;
        RECT 88.930 26.370 90.120 26.710 ;
        RECT 90.300 26.370 90.630 26.710 ;
      LAYER li1 ;
        RECT 82.810 24.810 82.820 24.980 ;
        RECT 82.990 24.810 83.180 24.980 ;
        RECT 83.350 24.810 83.370 24.980 ;
        RECT 82.810 24.730 83.370 24.810 ;
        RECT 84.980 24.930 87.720 25.810 ;
        RECT 84.980 24.760 85.190 24.930 ;
        RECT 85.360 24.760 85.630 24.930 ;
        RECT 85.800 24.760 86.040 24.930 ;
        RECT 86.210 24.760 86.470 24.930 ;
        RECT 86.640 24.760 86.910 24.930 ;
        RECT 87.080 24.760 87.320 24.930 ;
        RECT 87.490 24.760 87.720 24.930 ;
        RECT 84.980 24.740 87.720 24.760 ;
        RECT 88.890 24.980 90.560 26.190 ;
        RECT 88.890 24.810 88.920 24.980 ;
        RECT 89.090 24.810 89.280 24.980 ;
        RECT 89.450 24.810 89.640 24.980 ;
        RECT 89.810 24.810 90.000 24.980 ;
        RECT 90.170 24.810 90.360 24.980 ;
        RECT 90.530 24.810 90.560 24.980 ;
        RECT 88.890 24.730 90.560 24.810 ;
      LAYER li1 ;
        RECT 90.820 24.730 91.080 26.890 ;
      LAYER li1 ;
        RECT 91.680 26.460 92.010 27.240 ;
        RECT 94.650 27.140 95.960 27.920 ;
      LAYER li1 ;
        RECT 96.410 27.310 96.740 27.970 ;
      LAYER li1 ;
        RECT 97.130 27.920 97.180 28.090 ;
        RECT 97.350 27.920 97.620 28.090 ;
        RECT 97.790 27.920 98.060 28.090 ;
        RECT 98.230 27.920 98.470 28.090 ;
        RECT 98.640 27.920 98.740 28.090 ;
        RECT 97.130 27.640 98.740 27.920 ;
      LAYER li1 ;
        RECT 96.140 27.140 96.740 27.310 ;
      LAYER li1 ;
        RECT 97.440 27.240 98.740 27.640 ;
        RECT 98.970 28.090 99.560 28.120 ;
        RECT 98.970 27.920 99.000 28.090 ;
        RECT 99.170 27.920 99.360 28.090 ;
        RECT 99.530 27.920 99.560 28.090 ;
        RECT 100.490 28.090 102.100 28.120 ;
        RECT 102.790 28.090 104.040 28.120 ;
        RECT 104.810 28.090 106.420 28.120 ;
        RECT 107.110 28.090 108.360 28.120 ;
        RECT 109.130 28.090 110.740 28.120 ;
      LAYER li1 ;
        RECT 96.140 26.960 96.360 27.140 ;
      LAYER li1 ;
        RECT 92.220 25.800 92.550 26.790 ;
      LAYER li1 ;
        RECT 94.690 26.550 95.580 26.940 ;
        RECT 95.780 26.790 96.360 26.960 ;
      LAYER li1 ;
        RECT 91.450 24.930 92.900 25.800 ;
        RECT 91.450 24.760 91.700 24.930 ;
        RECT 91.870 24.760 92.060 24.930 ;
        RECT 92.230 24.760 92.500 24.930 ;
        RECT 92.670 24.760 92.900 24.930 ;
        RECT 91.450 24.730 92.900 24.760 ;
        RECT 94.650 24.980 95.600 26.310 ;
        RECT 94.650 24.810 94.680 24.980 ;
        RECT 94.850 24.810 95.040 24.980 ;
        RECT 95.210 24.810 95.400 24.980 ;
        RECT 95.570 24.810 95.600 24.980 ;
        RECT 94.650 24.730 95.600 24.810 ;
      LAYER li1 ;
        RECT 95.780 24.730 96.030 26.790 ;
        RECT 96.540 26.630 96.840 26.960 ;
      LAYER li1 ;
        RECT 97.440 26.460 97.770 27.240 ;
        RECT 98.970 27.160 99.560 27.920 ;
        RECT 96.220 24.980 96.810 26.310 ;
        RECT 97.980 25.800 98.310 26.790 ;
      LAYER li1 ;
        RECT 99.010 26.550 99.720 26.940 ;
        RECT 99.900 26.310 100.230 27.990 ;
      LAYER li1 ;
        RECT 100.490 27.920 100.540 28.090 ;
        RECT 100.710 27.920 100.980 28.090 ;
        RECT 101.150 27.920 101.420 28.090 ;
        RECT 101.590 27.920 101.830 28.090 ;
        RECT 102.000 27.920 102.100 28.090 ;
        RECT 100.490 27.640 102.100 27.920 ;
        RECT 100.800 27.240 102.100 27.640 ;
        RECT 100.800 26.460 101.130 27.240 ;
        RECT 96.220 24.810 96.250 24.980 ;
        RECT 96.420 24.810 96.610 24.980 ;
        RECT 96.780 24.810 96.810 24.980 ;
        RECT 96.220 24.730 96.810 24.810 ;
        RECT 97.210 24.930 98.660 25.800 ;
        RECT 97.210 24.760 97.460 24.930 ;
        RECT 97.630 24.760 97.820 24.930 ;
        RECT 97.990 24.760 98.260 24.930 ;
        RECT 98.430 24.760 98.660 24.930 ;
        RECT 97.210 24.730 98.660 24.760 ;
        RECT 98.970 24.980 99.560 26.310 ;
        RECT 98.970 24.810 99.000 24.980 ;
        RECT 99.170 24.810 99.360 24.980 ;
        RECT 99.530 24.810 99.560 24.980 ;
        RECT 98.970 24.730 99.560 24.810 ;
      LAYER li1 ;
        RECT 99.840 24.730 100.230 26.310 ;
      LAYER li1 ;
        RECT 101.340 25.800 101.670 26.790 ;
      LAYER li1 ;
        RECT 102.360 26.310 102.610 27.990 ;
      LAYER li1 ;
        RECT 102.960 27.920 103.150 28.090 ;
        RECT 103.320 27.920 103.510 28.090 ;
        RECT 103.680 27.920 103.870 28.090 ;
        RECT 102.790 27.550 104.040 27.920 ;
        RECT 104.220 27.370 104.470 27.990 ;
        RECT 104.810 27.920 104.860 28.090 ;
        RECT 105.030 27.920 105.300 28.090 ;
        RECT 105.470 27.920 105.740 28.090 ;
        RECT 105.910 27.920 106.150 28.090 ;
        RECT 106.320 27.920 106.420 28.090 ;
        RECT 104.810 27.640 106.420 27.920 ;
        RECT 102.920 27.200 104.470 27.370 ;
        RECT 102.920 26.740 103.250 27.200 ;
        RECT 100.570 24.930 102.020 25.800 ;
        RECT 100.570 24.760 100.820 24.930 ;
        RECT 100.990 24.760 101.180 24.930 ;
        RECT 101.350 24.760 101.620 24.930 ;
        RECT 101.790 24.760 102.020 24.930 ;
        RECT 100.570 24.730 102.020 24.760 ;
      LAYER li1 ;
        RECT 102.360 24.730 102.790 26.310 ;
      LAYER li1 ;
        RECT 102.970 24.980 103.530 26.310 ;
      LAYER li1 ;
        RECT 103.710 25.230 104.040 27.020 ;
      LAYER li1 ;
        RECT 104.220 25.480 104.470 27.200 ;
        RECT 105.120 27.240 106.420 27.640 ;
        RECT 105.120 26.460 105.450 27.240 ;
        RECT 105.660 25.800 105.990 26.790 ;
      LAYER li1 ;
        RECT 106.680 26.310 106.930 27.990 ;
      LAYER li1 ;
        RECT 107.280 27.920 107.470 28.090 ;
        RECT 107.640 27.920 107.830 28.090 ;
        RECT 108.000 27.920 108.190 28.090 ;
        RECT 107.110 27.550 108.360 27.920 ;
        RECT 108.540 27.370 108.790 27.990 ;
        RECT 109.130 27.920 109.180 28.090 ;
        RECT 109.350 27.920 109.620 28.090 ;
        RECT 109.790 27.920 110.060 28.090 ;
        RECT 110.230 27.920 110.470 28.090 ;
        RECT 110.640 27.920 110.740 28.090 ;
        RECT 109.130 27.640 110.740 27.920 ;
        RECT 107.240 27.200 108.790 27.370 ;
        RECT 107.240 26.740 107.570 27.200 ;
        RECT 102.970 24.810 102.980 24.980 ;
        RECT 103.150 24.810 103.340 24.980 ;
        RECT 103.510 24.810 103.530 24.980 ;
        RECT 102.970 24.730 103.530 24.810 ;
        RECT 104.890 24.930 106.340 25.800 ;
        RECT 104.890 24.760 105.140 24.930 ;
        RECT 105.310 24.760 105.500 24.930 ;
        RECT 105.670 24.760 105.940 24.930 ;
        RECT 106.110 24.760 106.340 24.930 ;
        RECT 104.890 24.730 106.340 24.760 ;
      LAYER li1 ;
        RECT 106.680 24.730 107.110 26.310 ;
      LAYER li1 ;
        RECT 107.290 24.980 107.850 26.310 ;
      LAYER li1 ;
        RECT 108.030 25.230 108.360 27.020 ;
      LAYER li1 ;
        RECT 108.540 25.480 108.790 27.200 ;
        RECT 109.440 27.240 110.740 27.640 ;
        RECT 110.970 28.090 112.280 28.120 ;
        RECT 110.970 27.920 111.000 28.090 ;
        RECT 111.170 27.920 111.360 28.090 ;
        RECT 111.530 27.920 111.720 28.090 ;
        RECT 111.890 27.920 112.080 28.090 ;
        RECT 112.250 27.920 112.280 28.090 ;
        RECT 113.450 28.090 115.060 28.120 ;
        RECT 109.440 26.460 109.770 27.240 ;
        RECT 110.970 27.140 112.280 27.920 ;
      LAYER li1 ;
        RECT 112.730 27.310 113.060 27.970 ;
      LAYER li1 ;
        RECT 113.450 27.920 113.500 28.090 ;
        RECT 113.670 27.920 113.940 28.090 ;
        RECT 114.110 27.920 114.380 28.090 ;
        RECT 114.550 27.920 114.790 28.090 ;
        RECT 114.960 27.920 115.060 28.090 ;
        RECT 113.450 27.640 115.060 27.920 ;
      LAYER li1 ;
        RECT 112.460 27.140 113.060 27.310 ;
      LAYER li1 ;
        RECT 113.760 27.240 115.060 27.640 ;
        RECT 115.290 28.090 115.880 28.120 ;
        RECT 115.290 27.920 115.320 28.090 ;
        RECT 115.490 27.920 115.680 28.090 ;
        RECT 115.850 27.920 115.880 28.090 ;
        RECT 116.560 28.090 117.510 28.120 ;
      LAYER li1 ;
        RECT 112.460 26.960 112.680 27.140 ;
      LAYER li1 ;
        RECT 109.980 25.800 110.310 26.790 ;
      LAYER li1 ;
        RECT 111.010 26.550 111.900 26.940 ;
        RECT 112.100 26.790 112.680 26.960 ;
      LAYER li1 ;
        RECT 107.290 24.810 107.300 24.980 ;
        RECT 107.470 24.810 107.660 24.980 ;
        RECT 107.830 24.810 107.850 24.980 ;
        RECT 107.290 24.730 107.850 24.810 ;
        RECT 109.210 24.930 110.660 25.800 ;
        RECT 109.210 24.760 109.460 24.930 ;
        RECT 109.630 24.760 109.820 24.930 ;
        RECT 109.990 24.760 110.260 24.930 ;
        RECT 110.430 24.760 110.660 24.930 ;
        RECT 109.210 24.730 110.660 24.760 ;
        RECT 110.970 24.980 111.920 26.310 ;
        RECT 110.970 24.810 111.000 24.980 ;
        RECT 111.170 24.810 111.360 24.980 ;
        RECT 111.530 24.810 111.720 24.980 ;
        RECT 111.890 24.810 111.920 24.980 ;
        RECT 110.970 24.730 111.920 24.810 ;
      LAYER li1 ;
        RECT 112.100 24.730 112.350 26.790 ;
        RECT 112.860 26.630 113.160 26.960 ;
      LAYER li1 ;
        RECT 113.760 26.460 114.090 27.240 ;
        RECT 115.290 27.160 115.880 27.920 ;
      LAYER li1 ;
        RECT 116.130 27.060 116.380 27.990 ;
      LAYER li1 ;
        RECT 116.560 27.920 116.590 28.090 ;
        RECT 116.760 27.920 116.950 28.090 ;
        RECT 117.120 27.920 117.310 28.090 ;
        RECT 117.480 27.920 117.510 28.090 ;
        RECT 118.730 28.090 120.340 28.120 ;
        RECT 116.560 27.240 117.510 27.920 ;
      LAYER li1 ;
        RECT 117.690 27.060 117.960 27.990 ;
      LAYER li1 ;
        RECT 118.730 27.920 118.780 28.090 ;
        RECT 118.950 27.920 119.220 28.090 ;
        RECT 119.390 27.920 119.660 28.090 ;
        RECT 119.830 27.920 120.070 28.090 ;
        RECT 120.240 27.920 120.340 28.090 ;
        RECT 118.730 27.640 120.340 27.920 ;
        RECT 112.540 24.980 113.130 26.310 ;
        RECT 114.300 25.800 114.630 26.790 ;
      LAYER li1 ;
        RECT 115.330 26.370 115.630 26.960 ;
        RECT 116.130 26.890 117.960 27.060 ;
        RECT 115.810 26.370 117.000 26.710 ;
      LAYER li1 ;
        RECT 112.540 24.810 112.570 24.980 ;
        RECT 112.740 24.810 112.930 24.980 ;
        RECT 113.100 24.810 113.130 24.980 ;
        RECT 112.540 24.730 113.130 24.810 ;
        RECT 113.530 24.930 114.980 25.800 ;
        RECT 113.530 24.760 113.780 24.930 ;
        RECT 113.950 24.760 114.140 24.930 ;
        RECT 114.310 24.760 114.580 24.930 ;
        RECT 114.750 24.760 114.980 24.930 ;
        RECT 113.530 24.730 114.980 24.760 ;
        RECT 115.290 24.980 116.960 26.190 ;
      LAYER li1 ;
        RECT 117.180 25.230 117.510 26.710 ;
      LAYER li1 ;
        RECT 115.290 24.810 115.320 24.980 ;
        RECT 115.490 24.810 115.680 24.980 ;
        RECT 115.850 24.810 116.040 24.980 ;
        RECT 116.210 24.810 116.400 24.980 ;
        RECT 116.570 24.810 116.760 24.980 ;
        RECT 116.930 24.810 116.960 24.980 ;
        RECT 115.290 24.730 116.960 24.810 ;
      LAYER li1 ;
        RECT 117.690 24.730 117.960 26.890 ;
      LAYER li1 ;
        RECT 119.040 27.240 120.340 27.640 ;
        RECT 120.810 28.090 122.520 28.120 ;
        RECT 120.810 27.920 120.860 28.090 ;
        RECT 121.030 27.920 121.220 28.090 ;
        RECT 121.390 27.920 121.580 28.090 ;
        RECT 121.750 27.920 121.940 28.090 ;
        RECT 122.110 27.920 122.300 28.090 ;
        RECT 122.470 27.920 122.520 28.090 ;
        RECT 123.160 28.090 123.750 28.120 ;
        RECT 119.040 26.460 119.370 27.240 ;
        RECT 120.810 27.160 122.520 27.920 ;
      LAYER li1 ;
        RECT 122.700 27.030 122.950 27.990 ;
      LAYER li1 ;
        RECT 123.160 27.920 123.190 28.090 ;
        RECT 123.360 27.920 123.550 28.090 ;
        RECT 123.720 27.920 123.750 28.090 ;
        RECT 123.160 27.210 123.750 27.920 ;
        RECT 124.010 28.090 125.620 28.120 ;
        RECT 124.010 27.920 124.060 28.090 ;
        RECT 124.230 27.920 124.500 28.090 ;
        RECT 124.670 27.920 124.940 28.090 ;
        RECT 125.110 27.920 125.350 28.090 ;
        RECT 125.520 27.920 125.620 28.090 ;
        RECT 124.010 27.640 125.620 27.920 ;
        RECT 124.320 27.240 125.620 27.640 ;
        RECT 125.850 28.090 126.440 28.120 ;
        RECT 125.850 27.920 125.880 28.090 ;
        RECT 126.050 27.920 126.240 28.090 ;
        RECT 126.410 27.920 126.440 28.090 ;
        RECT 127.370 28.090 128.980 28.120 ;
        RECT 129.670 28.090 130.920 28.120 ;
        RECT 131.690 28.090 133.300 28.120 ;
        RECT 119.580 25.800 119.910 26.790 ;
      LAYER li1 ;
        RECT 120.610 26.740 121.800 26.980 ;
        RECT 122.050 26.740 122.400 26.980 ;
        RECT 122.700 26.860 123.720 27.030 ;
      LAYER li1 ;
        RECT 120.740 26.390 122.770 26.560 ;
        RECT 118.810 24.930 120.260 25.800 ;
        RECT 118.810 24.760 119.060 24.930 ;
        RECT 119.230 24.760 119.420 24.930 ;
        RECT 119.590 24.760 119.860 24.930 ;
        RECT 120.030 24.760 120.260 24.930 ;
        RECT 118.810 24.730 120.260 24.760 ;
        RECT 120.740 24.730 120.990 26.390 ;
        RECT 121.170 24.980 122.420 26.210 ;
        RECT 121.340 24.810 121.530 24.980 ;
        RECT 121.700 24.810 121.890 24.980 ;
        RECT 122.060 24.810 122.250 24.980 ;
        RECT 121.170 24.730 122.420 24.810 ;
        RECT 122.600 24.730 122.770 26.390 ;
      LAYER li1 ;
        RECT 122.950 25.230 123.280 26.680 ;
        RECT 123.460 24.730 123.720 26.860 ;
      LAYER li1 ;
        RECT 124.320 26.460 124.650 27.240 ;
        RECT 125.850 27.160 126.440 27.920 ;
        RECT 124.860 25.800 125.190 26.790 ;
      LAYER li1 ;
        RECT 125.890 26.550 126.600 26.940 ;
        RECT 126.780 26.310 127.110 27.990 ;
      LAYER li1 ;
        RECT 127.370 27.920 127.420 28.090 ;
        RECT 127.590 27.920 127.860 28.090 ;
        RECT 128.030 27.920 128.300 28.090 ;
        RECT 128.470 27.920 128.710 28.090 ;
        RECT 128.880 27.920 128.980 28.090 ;
        RECT 127.370 27.640 128.980 27.920 ;
        RECT 127.680 27.240 128.980 27.640 ;
        RECT 127.680 26.460 128.010 27.240 ;
        RECT 124.090 24.930 125.540 25.800 ;
        RECT 124.090 24.760 124.340 24.930 ;
        RECT 124.510 24.760 124.700 24.930 ;
        RECT 124.870 24.760 125.140 24.930 ;
        RECT 125.310 24.760 125.540 24.930 ;
        RECT 124.090 24.730 125.540 24.760 ;
        RECT 125.850 24.980 126.440 26.310 ;
        RECT 125.850 24.810 125.880 24.980 ;
        RECT 126.050 24.810 126.240 24.980 ;
        RECT 126.410 24.810 126.440 24.980 ;
        RECT 125.850 24.730 126.440 24.810 ;
      LAYER li1 ;
        RECT 126.720 24.730 127.110 26.310 ;
      LAYER li1 ;
        RECT 128.220 25.800 128.550 26.790 ;
      LAYER li1 ;
        RECT 129.240 26.310 129.490 27.990 ;
      LAYER li1 ;
        RECT 129.840 27.920 130.030 28.090 ;
        RECT 130.200 27.920 130.390 28.090 ;
        RECT 130.560 27.920 130.750 28.090 ;
        RECT 129.670 27.550 130.920 27.920 ;
        RECT 131.100 27.370 131.350 27.990 ;
        RECT 131.690 27.920 131.740 28.090 ;
        RECT 131.910 27.920 132.180 28.090 ;
        RECT 132.350 27.920 132.620 28.090 ;
        RECT 132.790 27.920 133.030 28.090 ;
        RECT 133.200 27.920 133.300 28.090 ;
        RECT 135.940 28.090 136.590 28.200 ;
        RECT 131.690 27.640 133.300 27.920 ;
        RECT 129.800 27.200 131.350 27.370 ;
        RECT 129.800 26.740 130.130 27.200 ;
        RECT 127.450 24.930 128.900 25.800 ;
        RECT 127.450 24.760 127.700 24.930 ;
        RECT 127.870 24.760 128.060 24.930 ;
        RECT 128.230 24.760 128.500 24.930 ;
        RECT 128.670 24.760 128.900 24.930 ;
        RECT 127.450 24.730 128.900 24.760 ;
      LAYER li1 ;
        RECT 129.240 24.730 129.670 26.310 ;
      LAYER li1 ;
        RECT 129.850 24.980 130.410 26.310 ;
      LAYER li1 ;
        RECT 130.590 25.230 130.920 27.020 ;
      LAYER li1 ;
        RECT 131.100 25.480 131.350 27.200 ;
        RECT 132.000 27.240 133.300 27.640 ;
      LAYER li1 ;
        RECT 134.690 27.420 135.270 28.060 ;
      LAYER li1 ;
        RECT 135.940 27.920 136.000 28.090 ;
        RECT 136.170 27.920 136.360 28.090 ;
        RECT 136.530 27.920 136.590 28.090 ;
        RECT 135.940 27.860 136.590 27.920 ;
        RECT 136.180 27.420 136.590 27.860 ;
        RECT 137.380 28.100 140.110 28.130 ;
        RECT 137.380 27.930 137.550 28.100 ;
        RECT 137.720 27.930 137.990 28.100 ;
        RECT 138.160 27.930 138.400 28.100 ;
        RECT 138.570 27.930 138.830 28.100 ;
        RECT 139.000 27.930 139.270 28.100 ;
        RECT 139.440 27.930 139.680 28.100 ;
        RECT 139.850 27.930 140.110 28.100 ;
        RECT 132.000 26.460 132.330 27.240 ;
        RECT 132.540 25.800 132.870 26.790 ;
      LAYER li1 ;
        RECT 135.020 26.550 135.270 27.420 ;
      LAYER li1 ;
        RECT 137.380 27.130 140.110 27.930 ;
      LAYER li1 ;
        RECT 135.020 26.300 135.730 26.550 ;
      LAYER li1 ;
        RECT 137.540 26.460 137.870 27.130 ;
        RECT 129.850 24.810 129.860 24.980 ;
        RECT 130.030 24.810 130.220 24.980 ;
        RECT 130.390 24.810 130.410 24.980 ;
        RECT 129.850 24.730 130.410 24.810 ;
        RECT 131.770 24.930 133.220 25.800 ;
        RECT 131.770 24.760 132.020 24.930 ;
        RECT 132.190 24.760 132.380 24.930 ;
        RECT 132.550 24.760 132.820 24.930 ;
        RECT 132.990 24.760 133.220 24.930 ;
        RECT 131.770 24.730 133.220 24.760 ;
        RECT 134.620 25.040 135.020 25.310 ;
        RECT 134.620 24.980 135.270 25.040 ;
        RECT 134.620 24.810 134.680 24.980 ;
        RECT 134.850 24.810 135.040 24.980 ;
        RECT 135.210 24.810 135.270 24.980 ;
      LAYER li1 ;
        RECT 135.480 24.960 135.730 26.300 ;
      LAYER li1 ;
        RECT 138.270 25.810 138.600 26.790 ;
        RECT 138.820 26.460 139.150 27.130 ;
        RECT 139.550 25.810 139.880 26.790 ;
        RECT 134.620 24.700 135.270 24.810 ;
        RECT 137.300 24.930 140.040 25.810 ;
        RECT 137.300 24.760 137.510 24.930 ;
        RECT 137.680 24.760 137.950 24.930 ;
        RECT 138.120 24.760 138.360 24.930 ;
        RECT 138.530 24.760 138.790 24.930 ;
        RECT 138.960 24.760 139.230 24.930 ;
        RECT 139.400 24.760 139.640 24.930 ;
        RECT 139.810 24.760 140.040 24.930 ;
        RECT 137.300 24.740 140.040 24.760 ;
        RECT 5.760 24.330 5.920 24.510 ;
        RECT 6.090 24.330 6.400 24.510 ;
        RECT 6.570 24.330 6.880 24.510 ;
        RECT 7.050 24.330 7.360 24.510 ;
        RECT 7.530 24.330 7.840 24.510 ;
        RECT 8.010 24.330 8.320 24.510 ;
        RECT 8.490 24.330 8.800 24.510 ;
        RECT 8.970 24.330 9.280 24.510 ;
        RECT 9.450 24.330 9.760 24.510 ;
        RECT 9.930 24.330 10.240 24.510 ;
        RECT 10.410 24.330 10.720 24.510 ;
        RECT 10.890 24.330 11.200 24.510 ;
        RECT 11.370 24.330 11.680 24.510 ;
        RECT 11.850 24.330 12.160 24.510 ;
        RECT 12.330 24.330 12.640 24.510 ;
        RECT 12.810 24.330 13.120 24.510 ;
        RECT 13.290 24.330 13.600 24.510 ;
        RECT 13.770 24.330 14.080 24.510 ;
        RECT 14.250 24.500 14.560 24.510 ;
        RECT 14.730 24.500 15.040 24.510 ;
        RECT 14.250 24.330 14.400 24.500 ;
        RECT 14.880 24.330 15.040 24.500 ;
        RECT 15.210 24.330 15.520 24.510 ;
        RECT 15.690 24.330 16.000 24.510 ;
        RECT 16.170 24.330 16.480 24.510 ;
        RECT 16.650 24.500 16.800 24.510 ;
        RECT 17.280 24.500 17.440 24.510 ;
        RECT 16.650 24.330 16.960 24.500 ;
        RECT 17.130 24.330 17.440 24.500 ;
        RECT 17.610 24.330 17.920 24.510 ;
        RECT 18.090 24.330 18.400 24.510 ;
        RECT 18.570 24.330 18.880 24.510 ;
        RECT 19.050 24.330 19.360 24.510 ;
        RECT 19.530 24.330 19.840 24.510 ;
        RECT 20.010 24.330 20.320 24.510 ;
        RECT 20.490 24.330 20.800 24.510 ;
        RECT 20.970 24.330 21.280 24.510 ;
        RECT 21.450 24.330 21.760 24.510 ;
        RECT 21.930 24.330 22.240 24.510 ;
        RECT 22.410 24.330 22.720 24.510 ;
        RECT 22.890 24.330 23.200 24.510 ;
        RECT 23.370 24.330 23.680 24.510 ;
        RECT 23.850 24.330 24.160 24.510 ;
        RECT 24.330 24.330 24.640 24.510 ;
        RECT 24.810 24.330 25.120 24.510 ;
        RECT 25.290 24.330 25.600 24.510 ;
        RECT 25.770 24.330 26.080 24.510 ;
        RECT 26.250 24.330 26.560 24.510 ;
        RECT 26.730 24.330 27.040 24.510 ;
        RECT 27.210 24.330 27.520 24.510 ;
        RECT 27.690 24.330 28.000 24.510 ;
        RECT 28.170 24.330 28.480 24.510 ;
        RECT 28.650 24.330 28.960 24.510 ;
        RECT 29.130 24.330 29.440 24.510 ;
        RECT 29.610 24.330 29.920 24.510 ;
        RECT 30.090 24.330 30.400 24.510 ;
        RECT 30.570 24.330 30.880 24.510 ;
        RECT 31.050 24.330 31.360 24.510 ;
        RECT 31.530 24.330 31.840 24.510 ;
        RECT 32.010 24.330 32.320 24.510 ;
        RECT 32.490 24.330 32.800 24.510 ;
        RECT 32.970 24.330 33.280 24.510 ;
        RECT 33.450 24.330 33.760 24.510 ;
        RECT 33.930 24.330 34.240 24.510 ;
        RECT 34.410 24.330 34.720 24.510 ;
        RECT 34.890 24.330 35.200 24.510 ;
        RECT 35.370 24.330 35.680 24.510 ;
        RECT 35.850 24.330 36.160 24.510 ;
        RECT 36.330 24.330 36.640 24.510 ;
        RECT 36.810 24.330 37.120 24.510 ;
        RECT 37.290 24.330 37.600 24.510 ;
        RECT 37.770 24.330 38.080 24.510 ;
        RECT 38.250 24.330 38.560 24.510 ;
        RECT 38.730 24.330 39.040 24.510 ;
        RECT 39.210 24.330 39.520 24.510 ;
        RECT 39.690 24.330 40.000 24.510 ;
        RECT 40.170 24.330 40.480 24.510 ;
        RECT 40.650 24.330 40.960 24.510 ;
        RECT 41.130 24.330 41.440 24.510 ;
        RECT 41.610 24.330 41.920 24.510 ;
        RECT 42.090 24.330 42.400 24.510 ;
        RECT 42.570 24.330 42.880 24.510 ;
        RECT 43.050 24.330 43.360 24.510 ;
        RECT 43.530 24.330 43.840 24.510 ;
        RECT 44.010 24.330 44.320 24.510 ;
        RECT 44.490 24.330 44.800 24.510 ;
        RECT 44.970 24.330 45.280 24.510 ;
        RECT 45.450 24.330 45.760 24.510 ;
        RECT 45.930 24.330 46.240 24.510 ;
        RECT 46.410 24.330 46.720 24.510 ;
        RECT 46.890 24.330 47.200 24.510 ;
        RECT 47.370 24.330 47.680 24.510 ;
        RECT 47.850 24.330 48.160 24.510 ;
        RECT 48.330 24.330 48.640 24.510 ;
        RECT 48.810 24.330 49.120 24.510 ;
        RECT 49.290 24.330 49.600 24.510 ;
        RECT 49.770 24.330 50.080 24.510 ;
        RECT 50.250 24.330 50.560 24.510 ;
        RECT 50.730 24.330 51.040 24.510 ;
        RECT 51.210 24.330 51.520 24.510 ;
        RECT 51.690 24.330 52.000 24.510 ;
        RECT 52.170 24.500 52.480 24.510 ;
        RECT 52.650 24.500 52.960 24.510 ;
        RECT 52.170 24.330 52.320 24.500 ;
        RECT 52.800 24.330 52.960 24.500 ;
        RECT 53.130 24.330 53.440 24.510 ;
        RECT 53.610 24.330 53.920 24.510 ;
        RECT 54.090 24.330 54.400 24.510 ;
        RECT 54.570 24.330 54.880 24.510 ;
        RECT 55.050 24.330 55.360 24.510 ;
        RECT 55.530 24.330 55.840 24.510 ;
        RECT 56.010 24.330 56.320 24.510 ;
        RECT 56.490 24.330 56.800 24.510 ;
        RECT 56.970 24.330 57.280 24.510 ;
        RECT 57.450 24.330 57.760 24.510 ;
        RECT 57.930 24.330 58.240 24.510 ;
        RECT 58.410 24.330 58.720 24.510 ;
        RECT 58.890 24.330 59.200 24.510 ;
        RECT 59.370 24.330 59.680 24.510 ;
        RECT 59.850 24.330 60.160 24.510 ;
        RECT 60.330 24.330 60.640 24.510 ;
        RECT 60.810 24.330 61.120 24.510 ;
        RECT 61.290 24.330 61.600 24.510 ;
        RECT 61.770 24.330 62.080 24.510 ;
        RECT 62.250 24.330 62.560 24.510 ;
        RECT 62.730 24.330 63.040 24.510 ;
        RECT 63.210 24.330 63.520 24.510 ;
        RECT 63.690 24.330 64.000 24.510 ;
        RECT 64.170 24.330 64.480 24.510 ;
        RECT 64.650 24.330 64.960 24.510 ;
        RECT 65.130 24.330 65.440 24.510 ;
        RECT 65.610 24.330 65.920 24.510 ;
        RECT 66.090 24.330 66.400 24.510 ;
        RECT 66.570 24.330 66.880 24.510 ;
        RECT 67.050 24.330 67.360 24.510 ;
        RECT 67.530 24.330 67.840 24.510 ;
        RECT 68.010 24.330 68.320 24.510 ;
        RECT 68.490 24.330 68.800 24.510 ;
        RECT 68.970 24.330 69.280 24.510 ;
        RECT 69.450 24.330 69.760 24.510 ;
        RECT 69.930 24.330 70.240 24.510 ;
        RECT 70.410 24.330 70.720 24.510 ;
        RECT 70.890 24.330 71.200 24.510 ;
        RECT 71.370 24.330 71.680 24.510 ;
        RECT 71.850 24.330 72.160 24.510 ;
        RECT 72.330 24.330 72.640 24.510 ;
        RECT 72.810 24.330 73.120 24.510 ;
        RECT 73.290 24.330 73.600 24.510 ;
        RECT 73.770 24.330 74.080 24.510 ;
        RECT 74.250 24.330 74.560 24.510 ;
        RECT 74.730 24.330 75.040 24.510 ;
        RECT 75.210 24.330 75.520 24.510 ;
        RECT 75.690 24.330 76.000 24.510 ;
        RECT 76.170 24.330 76.480 24.510 ;
        RECT 76.650 24.330 76.960 24.510 ;
        RECT 77.130 24.330 77.440 24.510 ;
        RECT 77.610 24.330 77.920 24.510 ;
        RECT 78.090 24.330 78.400 24.510 ;
        RECT 78.570 24.330 78.880 24.510 ;
        RECT 79.050 24.330 79.360 24.510 ;
        RECT 79.530 24.330 79.840 24.510 ;
        RECT 80.010 24.330 80.320 24.510 ;
        RECT 80.490 24.330 80.800 24.510 ;
        RECT 80.970 24.330 81.280 24.510 ;
        RECT 81.450 24.500 81.760 24.510 ;
        RECT 81.930 24.500 82.240 24.510 ;
        RECT 81.450 24.330 81.600 24.500 ;
        RECT 82.080 24.330 82.240 24.500 ;
        RECT 82.410 24.330 82.720 24.510 ;
        RECT 82.890 24.330 83.200 24.510 ;
        RECT 83.370 24.330 83.680 24.510 ;
        RECT 83.850 24.330 84.160 24.510 ;
        RECT 84.330 24.330 84.640 24.510 ;
        RECT 84.810 24.330 85.120 24.510 ;
        RECT 85.290 24.330 85.600 24.510 ;
        RECT 85.770 24.330 86.080 24.510 ;
        RECT 86.250 24.330 86.560 24.510 ;
        RECT 86.730 24.330 87.040 24.510 ;
        RECT 87.210 24.330 87.520 24.510 ;
        RECT 87.690 24.330 88.000 24.510 ;
        RECT 88.170 24.500 88.480 24.510 ;
        RECT 88.650 24.500 88.960 24.510 ;
        RECT 88.170 24.330 88.320 24.500 ;
        RECT 88.800 24.330 88.960 24.500 ;
        RECT 89.130 24.330 89.440 24.510 ;
        RECT 89.610 24.330 89.920 24.510 ;
        RECT 90.090 24.330 90.400 24.510 ;
        RECT 90.570 24.330 90.880 24.510 ;
        RECT 91.050 24.330 91.360 24.510 ;
        RECT 91.530 24.330 91.840 24.510 ;
        RECT 92.010 24.330 92.320 24.510 ;
        RECT 92.490 24.330 92.800 24.510 ;
        RECT 92.970 24.330 93.280 24.510 ;
        RECT 93.450 24.330 93.760 24.510 ;
        RECT 93.930 24.500 94.240 24.510 ;
        RECT 94.410 24.500 94.720 24.510 ;
        RECT 93.930 24.330 94.080 24.500 ;
        RECT 94.560 24.330 94.720 24.500 ;
        RECT 94.890 24.330 95.200 24.510 ;
        RECT 95.370 24.330 95.680 24.510 ;
        RECT 95.850 24.330 96.160 24.510 ;
        RECT 96.330 24.330 96.640 24.510 ;
        RECT 96.810 24.330 97.120 24.510 ;
        RECT 97.290 24.330 97.600 24.510 ;
        RECT 97.770 24.330 98.080 24.510 ;
        RECT 98.250 24.330 98.560 24.510 ;
        RECT 98.730 24.330 99.040 24.510 ;
        RECT 99.210 24.330 99.520 24.510 ;
        RECT 99.690 24.330 100.000 24.510 ;
        RECT 100.170 24.330 100.480 24.510 ;
        RECT 100.650 24.330 100.960 24.510 ;
        RECT 101.130 24.330 101.440 24.510 ;
        RECT 101.610 24.330 101.920 24.510 ;
        RECT 102.090 24.330 102.400 24.510 ;
        RECT 102.570 24.330 102.880 24.510 ;
        RECT 103.050 24.330 103.360 24.510 ;
        RECT 103.530 24.330 103.840 24.510 ;
        RECT 104.010 24.330 104.320 24.510 ;
        RECT 104.490 24.330 104.800 24.510 ;
        RECT 104.970 24.330 105.280 24.510 ;
        RECT 105.450 24.330 105.760 24.510 ;
        RECT 105.930 24.330 106.240 24.510 ;
        RECT 106.410 24.330 106.720 24.510 ;
        RECT 106.890 24.330 107.200 24.510 ;
        RECT 107.370 24.330 107.680 24.510 ;
        RECT 107.850 24.330 108.160 24.510 ;
        RECT 108.330 24.330 108.640 24.510 ;
        RECT 108.810 24.330 109.120 24.510 ;
        RECT 109.290 24.330 109.600 24.510 ;
        RECT 109.770 24.330 110.080 24.510 ;
        RECT 110.250 24.330 110.560 24.510 ;
        RECT 110.730 24.330 111.040 24.510 ;
        RECT 111.210 24.330 111.520 24.510 ;
        RECT 111.690 24.330 112.000 24.510 ;
        RECT 112.170 24.330 112.480 24.510 ;
        RECT 112.650 24.330 112.960 24.510 ;
        RECT 113.130 24.330 113.440 24.510 ;
        RECT 113.610 24.330 113.920 24.510 ;
        RECT 114.090 24.330 114.400 24.510 ;
        RECT 114.570 24.330 114.880 24.510 ;
        RECT 115.050 24.330 115.360 24.510 ;
        RECT 115.530 24.330 115.840 24.510 ;
        RECT 116.010 24.330 116.320 24.510 ;
        RECT 116.490 24.330 116.800 24.510 ;
        RECT 116.970 24.330 117.280 24.510 ;
        RECT 117.450 24.330 117.760 24.510 ;
        RECT 117.930 24.330 118.240 24.510 ;
        RECT 118.410 24.330 118.720 24.510 ;
        RECT 118.890 24.330 119.200 24.510 ;
        RECT 119.370 24.330 119.680 24.510 ;
        RECT 119.850 24.330 120.160 24.510 ;
        RECT 120.330 24.330 120.640 24.510 ;
        RECT 120.810 24.330 121.120 24.510 ;
        RECT 121.290 24.330 121.600 24.510 ;
        RECT 121.770 24.330 122.080 24.510 ;
        RECT 122.250 24.330 122.560 24.510 ;
        RECT 122.730 24.330 123.040 24.510 ;
        RECT 123.210 24.330 123.520 24.510 ;
        RECT 123.690 24.330 124.000 24.510 ;
        RECT 124.170 24.330 124.480 24.510 ;
        RECT 124.650 24.330 124.960 24.510 ;
        RECT 125.130 24.330 125.440 24.510 ;
        RECT 125.610 24.330 125.920 24.510 ;
        RECT 126.090 24.330 126.400 24.510 ;
        RECT 126.570 24.330 126.880 24.510 ;
        RECT 127.050 24.330 127.360 24.510 ;
        RECT 127.530 24.330 127.840 24.510 ;
        RECT 128.010 24.330 128.320 24.510 ;
        RECT 128.490 24.330 128.800 24.510 ;
        RECT 128.970 24.330 129.280 24.510 ;
        RECT 129.450 24.330 129.760 24.510 ;
        RECT 129.930 24.330 130.240 24.510 ;
        RECT 130.410 24.330 130.720 24.510 ;
        RECT 130.890 24.330 131.200 24.510 ;
        RECT 131.370 24.330 131.680 24.510 ;
        RECT 131.850 24.330 132.160 24.510 ;
        RECT 132.330 24.330 132.640 24.510 ;
        RECT 132.810 24.330 133.120 24.510 ;
        RECT 133.290 24.330 133.600 24.510 ;
        RECT 133.770 24.330 134.080 24.510 ;
        RECT 134.250 24.330 134.560 24.510 ;
        RECT 134.730 24.330 135.040 24.510 ;
        RECT 135.210 24.330 135.520 24.510 ;
        RECT 135.690 24.330 136.000 24.510 ;
        RECT 136.170 24.330 136.480 24.510 ;
        RECT 136.650 24.330 136.960 24.510 ;
        RECT 137.130 24.330 137.440 24.510 ;
        RECT 137.610 24.330 137.920 24.510 ;
        RECT 138.090 24.330 138.400 24.510 ;
        RECT 138.570 24.330 138.880 24.510 ;
        RECT 139.050 24.330 139.360 24.510 ;
        RECT 139.530 24.330 139.840 24.510 ;
        RECT 140.010 24.330 140.320 24.510 ;
        RECT 140.490 24.330 140.800 24.510 ;
        RECT 140.970 24.330 141.280 24.510 ;
        RECT 141.450 24.500 141.760 24.510 ;
        RECT 141.930 24.500 142.080 24.510 ;
        RECT 141.450 24.330 141.600 24.500 ;
        RECT 6.260 24.080 9.000 24.100 ;
        RECT 6.260 23.910 6.470 24.080 ;
        RECT 6.640 23.910 6.910 24.080 ;
        RECT 7.080 23.910 7.320 24.080 ;
        RECT 7.490 23.910 7.750 24.080 ;
        RECT 7.920 23.910 8.190 24.080 ;
        RECT 8.360 23.910 8.600 24.080 ;
        RECT 8.770 23.910 9.000 24.080 ;
        RECT 6.260 23.030 9.000 23.910 ;
        RECT 10.780 24.030 11.430 24.140 ;
        RECT 10.780 23.860 10.840 24.030 ;
        RECT 11.010 23.860 11.200 24.030 ;
        RECT 11.370 23.860 11.430 24.030 ;
        RECT 13.460 24.080 16.200 24.100 ;
        RECT 13.460 23.910 13.670 24.080 ;
        RECT 13.840 23.910 14.110 24.080 ;
        RECT 14.280 23.910 14.520 24.080 ;
        RECT 14.690 23.910 14.950 24.080 ;
        RECT 15.120 23.910 15.390 24.080 ;
        RECT 15.560 23.910 15.800 24.080 ;
        RECT 15.970 23.910 16.200 24.080 ;
        RECT 10.780 23.800 11.430 23.860 ;
        RECT 10.780 23.530 11.180 23.800 ;
        RECT 6.500 21.710 6.830 22.380 ;
        RECT 7.230 22.050 7.560 23.030 ;
        RECT 7.780 21.710 8.110 22.380 ;
        RECT 8.510 22.050 8.840 23.030 ;
      LAYER li1 ;
        RECT 11.640 22.540 11.890 23.880 ;
      LAYER li1 ;
        RECT 13.460 23.030 16.200 23.910 ;
        RECT 17.500 24.030 18.150 24.140 ;
        RECT 17.500 23.860 17.560 24.030 ;
        RECT 17.730 23.860 17.920 24.030 ;
        RECT 18.090 23.860 18.150 24.030 ;
        RECT 19.930 24.080 21.380 24.110 ;
        RECT 19.930 23.910 20.180 24.080 ;
        RECT 20.350 23.910 20.540 24.080 ;
        RECT 20.710 23.910 20.980 24.080 ;
        RECT 21.150 23.910 21.380 24.080 ;
        RECT 17.500 23.800 18.150 23.860 ;
        RECT 17.500 23.530 17.900 23.800 ;
      LAYER li1 ;
        RECT 11.180 22.290 11.890 22.540 ;
      LAYER li1 ;
        RECT 6.340 20.710 9.070 21.710 ;
      LAYER li1 ;
        RECT 11.180 21.420 11.430 22.290 ;
      LAYER li1 ;
        RECT 13.700 21.710 14.030 22.380 ;
        RECT 14.430 22.050 14.760 23.030 ;
        RECT 14.980 21.710 15.310 22.380 ;
        RECT 15.710 22.050 16.040 23.030 ;
      LAYER li1 ;
        RECT 18.360 22.540 18.610 23.880 ;
      LAYER li1 ;
        RECT 19.930 23.040 21.380 23.910 ;
        RECT 21.820 24.030 22.470 24.140 ;
        RECT 21.820 23.860 21.880 24.030 ;
        RECT 22.050 23.860 22.240 24.030 ;
        RECT 22.410 23.860 22.470 24.030 ;
        RECT 21.820 23.800 22.470 23.860 ;
        RECT 21.820 23.530 22.220 23.800 ;
      LAYER li1 ;
        RECT 23.130 23.530 23.710 24.170 ;
      LAYER li1 ;
        RECT 24.250 24.080 25.700 24.110 ;
        RECT 24.250 23.910 24.500 24.080 ;
        RECT 24.670 23.910 24.860 24.080 ;
        RECT 25.030 23.910 25.300 24.080 ;
        RECT 25.470 23.910 25.700 24.080 ;
      LAYER li1 ;
        RECT 17.900 22.290 18.610 22.540 ;
        RECT 10.850 20.780 11.430 21.420 ;
      LAYER li1 ;
        RECT 12.340 20.980 12.750 21.420 ;
        RECT 12.100 20.640 12.750 20.980 ;
        RECT 13.540 20.710 16.270 21.710 ;
      LAYER li1 ;
        RECT 17.900 21.420 18.150 22.290 ;
      LAYER li1 ;
        RECT 20.160 21.600 20.490 22.380 ;
        RECT 20.700 22.050 21.030 23.040 ;
      LAYER li1 ;
        RECT 23.130 22.120 23.400 23.530 ;
      LAYER li1 ;
        RECT 24.250 23.040 25.700 23.910 ;
        RECT 26.550 24.030 27.140 24.060 ;
        RECT 26.550 23.860 26.580 24.030 ;
        RECT 26.750 23.860 26.940 24.030 ;
        RECT 27.110 23.860 27.140 24.030 ;
      LAYER li1 ;
        RECT 22.640 21.850 23.400 22.120 ;
        RECT 17.570 20.780 18.150 21.420 ;
      LAYER li1 ;
        RECT 19.060 20.980 19.470 21.420 ;
        RECT 20.160 21.200 21.460 21.600 ;
        RECT 18.820 20.640 19.470 20.980 ;
        RECT 19.850 20.720 21.460 21.200 ;
      LAYER li1 ;
        RECT 22.640 20.850 22.970 21.850 ;
      LAYER li1 ;
        RECT 24.480 21.600 24.810 22.380 ;
        RECT 25.020 22.050 25.350 23.040 ;
        RECT 26.030 22.880 26.360 23.810 ;
        RECT 26.550 23.080 27.140 23.860 ;
        RECT 27.320 23.990 28.760 24.160 ;
        RECT 27.320 22.880 27.490 23.990 ;
        RECT 26.030 22.710 27.490 22.880 ;
        RECT 23.380 20.980 23.790 21.420 ;
        RECT 24.480 21.200 25.780 21.600 ;
        RECT 23.140 20.640 23.790 20.980 ;
        RECT 24.170 20.720 25.780 21.200 ;
        RECT 26.030 20.850 26.300 22.710 ;
        RECT 27.160 22.210 27.490 22.710 ;
        RECT 27.670 22.500 27.920 23.810 ;
        RECT 28.160 23.190 28.410 23.810 ;
        RECT 28.590 23.540 28.760 23.990 ;
        RECT 28.940 24.030 29.270 24.060 ;
        RECT 28.940 23.860 28.970 24.030 ;
        RECT 29.140 23.860 29.270 24.030 ;
        RECT 28.940 23.720 29.270 23.860 ;
        RECT 29.450 23.990 31.190 24.160 ;
        RECT 29.450 23.540 29.620 23.990 ;
        RECT 28.590 23.370 29.620 23.540 ;
        RECT 29.800 23.190 29.970 23.810 ;
        RECT 30.500 23.550 30.830 23.810 ;
        RECT 28.160 23.020 29.970 23.190 ;
        RECT 30.150 23.020 30.370 23.350 ;
        RECT 29.800 22.840 29.970 23.020 ;
        RECT 27.670 22.270 28.200 22.500 ;
        RECT 27.670 21.350 27.940 22.270 ;
      LAYER li1 ;
        RECT 28.620 21.970 29.160 22.840 ;
      LAYER li1 ;
        RECT 29.800 22.670 30.020 22.840 ;
        RECT 26.480 20.720 27.430 21.350 ;
        RECT 27.610 20.850 27.940 21.350 ;
        RECT 28.120 20.720 28.710 21.600 ;
      LAYER li1 ;
        RECT 28.990 21.360 29.160 21.970 ;
        RECT 28.950 21.190 29.160 21.360 ;
        RECT 28.990 20.980 29.160 21.190 ;
        RECT 29.340 21.160 29.670 22.460 ;
      LAYER li1 ;
        RECT 29.850 21.680 30.020 22.670 ;
        RECT 30.200 22.500 30.370 23.020 ;
        RECT 30.550 22.850 30.720 23.550 ;
        RECT 31.020 23.400 31.190 23.990 ;
        RECT 31.370 24.030 32.320 24.060 ;
        RECT 31.370 23.860 31.400 24.030 ;
        RECT 31.570 23.860 31.760 24.030 ;
        RECT 31.930 23.860 32.120 24.030 ;
        RECT 32.290 23.860 32.320 24.030 ;
        RECT 31.370 23.580 32.320 23.860 ;
        RECT 32.500 23.990 33.530 24.160 ;
        RECT 32.500 23.400 32.670 23.990 ;
        RECT 31.020 23.350 32.670 23.400 ;
        RECT 30.900 23.230 32.670 23.350 ;
        RECT 30.900 23.030 31.230 23.230 ;
        RECT 32.850 23.050 33.180 23.810 ;
        RECT 33.360 23.630 33.530 23.990 ;
        RECT 33.710 24.030 34.660 24.110 ;
        RECT 33.710 23.860 33.740 24.030 ;
        RECT 33.910 23.860 34.100 24.030 ;
        RECT 34.270 23.860 34.460 24.030 ;
        RECT 34.630 23.860 34.660 24.030 ;
        RECT 33.710 23.810 34.660 23.860 ;
        RECT 33.360 23.460 35.170 23.630 ;
        RECT 31.410 22.880 33.180 23.050 ;
        RECT 31.410 22.850 31.580 22.880 ;
        RECT 30.550 22.680 31.580 22.850 ;
        RECT 34.490 22.700 34.820 23.280 ;
        RECT 30.200 22.270 31.230 22.500 ;
        RECT 30.900 21.780 31.230 22.270 ;
        RECT 31.410 22.000 31.580 22.680 ;
        RECT 31.760 22.530 34.820 22.700 ;
        RECT 31.760 22.180 32.090 22.530 ;
      LAYER li1 ;
        RECT 32.530 22.180 34.380 22.350 ;
      LAYER li1 ;
        RECT 31.410 21.830 34.030 22.000 ;
        RECT 29.850 21.180 30.120 21.680 ;
        RECT 31.410 21.600 31.580 21.830 ;
      LAYER li1 ;
        RECT 34.210 21.650 34.380 22.180 ;
      LAYER li1 ;
        RECT 30.570 21.430 31.580 21.600 ;
      LAYER li1 ;
        RECT 31.760 21.480 34.380 21.650 ;
      LAYER li1 ;
        RECT 30.570 21.180 30.900 21.430 ;
      LAYER li1 ;
        RECT 31.760 20.980 31.930 21.480 ;
        RECT 28.990 20.810 31.930 20.980 ;
      LAYER li1 ;
        RECT 33.080 20.720 34.030 21.300 ;
      LAYER li1 ;
        RECT 34.210 20.790 34.380 21.480 ;
      LAYER li1 ;
        RECT 34.560 21.680 34.820 22.530 ;
        RECT 35.000 22.110 35.170 23.460 ;
        RECT 35.350 23.200 35.600 24.110 ;
        RECT 36.410 24.030 37.360 24.060 ;
        RECT 38.190 24.030 39.090 24.060 ;
        RECT 36.410 23.860 36.440 24.030 ;
        RECT 36.610 23.860 36.800 24.030 ;
        RECT 36.970 23.860 37.160 24.030 ;
        RECT 37.330 23.860 37.360 24.030 ;
        RECT 38.360 23.860 38.550 24.030 ;
        RECT 38.720 23.860 38.910 24.030 ;
        RECT 39.080 23.860 39.090 24.030 ;
        RECT 35.350 23.030 36.230 23.200 ;
        RECT 36.410 23.030 37.360 23.860 ;
        RECT 37.760 23.060 38.010 23.530 ;
        RECT 38.190 23.240 39.090 23.860 ;
        RECT 39.700 24.030 40.640 24.090 ;
        RECT 39.700 23.860 39.720 24.030 ;
        RECT 39.890 23.860 40.080 24.030 ;
        RECT 40.250 23.860 40.440 24.030 ;
        RECT 40.610 23.860 40.640 24.030 ;
        RECT 35.550 22.290 35.880 22.790 ;
        RECT 36.060 22.710 36.230 23.030 ;
        RECT 37.760 22.890 38.770 23.060 ;
        RECT 36.060 22.540 38.420 22.710 ;
        RECT 35.000 21.940 36.170 22.110 ;
        RECT 34.560 20.970 34.890 21.680 ;
        RECT 35.350 21.140 35.680 21.680 ;
        RECT 35.890 21.440 36.170 21.940 ;
        RECT 36.350 21.140 36.520 22.540 ;
        RECT 38.600 22.360 38.770 22.890 ;
        RECT 36.730 22.190 38.770 22.360 ;
        RECT 36.730 21.800 37.060 22.190 ;
      LAYER li1 ;
        RECT 37.380 21.620 37.710 22.010 ;
      LAYER li1 ;
        RECT 35.350 20.970 36.520 21.140 ;
      LAYER li1 ;
        RECT 36.700 21.450 37.710 21.620 ;
        RECT 36.700 20.790 36.870 21.450 ;
      LAYER li1 ;
        RECT 38.540 21.350 38.770 22.190 ;
        RECT 39.270 22.360 39.520 23.360 ;
        RECT 39.700 22.550 40.640 23.860 ;
        RECT 39.270 22.030 40.640 22.360 ;
        RECT 39.270 21.850 39.480 22.030 ;
        RECT 39.150 21.350 39.480 21.850 ;
      LAYER li1 ;
        RECT 34.210 20.620 36.870 20.790 ;
      LAYER li1 ;
        RECT 37.050 20.720 38.000 21.270 ;
        RECT 38.540 20.850 38.870 21.350 ;
        RECT 39.660 20.720 40.610 21.850 ;
      LAYER li1 ;
        RECT 40.820 21.020 41.160 24.090 ;
      LAYER li1 ;
        RECT 41.780 24.080 44.520 24.100 ;
        RECT 41.780 23.910 41.990 24.080 ;
        RECT 42.160 23.910 42.430 24.080 ;
        RECT 42.600 23.910 42.840 24.080 ;
        RECT 43.010 23.910 43.270 24.080 ;
        RECT 43.440 23.910 43.710 24.080 ;
        RECT 43.880 23.910 44.120 24.080 ;
        RECT 44.290 23.910 44.520 24.080 ;
        RECT 41.780 23.030 44.520 23.910 ;
        RECT 42.020 21.710 42.350 22.380 ;
        RECT 42.750 22.050 43.080 23.030 ;
        RECT 43.300 21.710 43.630 22.380 ;
        RECT 44.030 22.050 44.360 23.030 ;
        RECT 45.240 21.820 45.490 24.090 ;
        RECT 45.670 24.030 46.620 24.110 ;
        RECT 45.670 23.860 45.700 24.030 ;
        RECT 45.870 23.860 46.060 24.030 ;
        RECT 46.230 23.860 46.420 24.030 ;
        RECT 46.590 23.860 46.620 24.030 ;
        RECT 45.670 23.280 46.620 23.860 ;
        RECT 46.800 23.300 47.130 24.090 ;
        RECT 46.810 22.800 47.130 23.300 ;
        RECT 47.360 24.030 47.610 24.060 ;
        RECT 47.360 23.860 47.390 24.030 ;
        RECT 47.560 23.860 47.610 24.030 ;
        RECT 47.360 22.980 47.610 23.860 ;
        RECT 47.790 22.800 47.960 24.110 ;
        RECT 50.730 24.030 51.060 24.060 ;
        RECT 46.810 22.630 47.960 22.800 ;
        RECT 48.140 23.640 50.130 23.970 ;
        RECT 46.300 21.820 46.630 22.250 ;
        RECT 41.860 20.710 44.590 21.710 ;
        RECT 45.240 21.650 46.630 21.820 ;
        RECT 45.240 20.970 45.500 21.650 ;
        RECT 45.690 20.720 46.280 21.470 ;
        RECT 46.460 20.790 46.630 21.650 ;
        RECT 46.810 20.970 47.060 22.630 ;
      LAYER li1 ;
        RECT 47.630 21.880 47.960 22.450 ;
      LAYER li1 ;
        RECT 48.140 21.700 48.310 23.640 ;
        RECT 47.240 21.530 48.310 21.700 ;
        RECT 47.240 20.790 47.410 21.530 ;
        RECT 48.490 21.350 48.660 23.460 ;
        RECT 48.840 21.440 49.010 23.640 ;
        RECT 49.190 22.960 49.520 23.460 ;
        RECT 49.190 21.490 49.360 22.960 ;
        RECT 49.960 22.680 50.130 23.640 ;
        RECT 50.310 23.030 50.550 23.910 ;
        RECT 50.730 23.860 50.760 24.030 ;
        RECT 50.930 23.860 51.060 24.030 ;
        RECT 50.730 23.210 51.060 23.860 ;
        RECT 52.200 24.030 53.150 24.060 ;
        RECT 52.200 23.860 52.230 24.030 ;
        RECT 52.400 23.860 52.590 24.030 ;
        RECT 52.760 23.860 52.950 24.030 ;
        RECT 53.120 23.860 53.150 24.030 ;
        RECT 51.690 23.200 52.020 23.460 ;
        RECT 51.240 23.030 52.020 23.200 ;
        RECT 52.200 23.030 53.150 23.860 ;
        RECT 53.820 23.950 54.950 24.160 ;
        RECT 55.130 24.030 56.080 24.060 ;
        RECT 53.820 23.200 53.990 23.950 ;
        RECT 55.130 23.860 55.160 24.030 ;
        RECT 55.330 23.860 55.520 24.030 ;
        RECT 55.690 23.860 55.880 24.030 ;
        RECT 56.050 23.860 56.080 24.030 ;
        RECT 54.170 23.380 54.780 23.770 ;
        RECT 53.820 23.030 54.430 23.200 ;
        RECT 50.310 22.860 51.410 23.030 ;
        RECT 51.590 22.680 54.080 22.850 ;
        RECT 49.540 22.330 49.780 22.520 ;
        RECT 49.960 22.510 51.760 22.680 ;
        RECT 51.940 22.330 53.570 22.500 ;
        RECT 53.750 22.440 54.080 22.680 ;
        RECT 49.540 22.160 52.110 22.330 ;
        RECT 53.400 22.230 53.570 22.330 ;
        RECT 54.260 22.230 54.430 23.030 ;
        RECT 49.540 21.850 49.780 22.160 ;
        RECT 50.260 21.670 50.990 21.980 ;
      LAYER li1 ;
        RECT 52.290 21.910 53.220 22.150 ;
      LAYER li1 ;
        RECT 46.460 20.620 47.410 20.790 ;
        RECT 47.590 20.720 48.130 21.350 ;
        RECT 48.310 20.850 48.660 21.350 ;
        RECT 49.190 21.320 51.440 21.490 ;
        RECT 49.190 20.850 49.440 21.320 ;
        RECT 49.980 20.720 50.930 21.140 ;
        RECT 51.110 20.620 51.440 21.320 ;
        RECT 51.920 20.720 52.870 21.730 ;
      LAYER li1 ;
        RECT 53.050 21.360 53.220 21.910 ;
      LAYER li1 ;
        RECT 53.400 22.060 54.430 22.230 ;
        RECT 54.610 22.840 54.780 23.380 ;
        RECT 55.130 23.020 56.080 23.860 ;
        RECT 56.420 23.610 56.670 24.110 ;
        RECT 56.850 24.030 57.800 24.090 ;
        RECT 60.500 24.080 63.240 24.100 ;
        RECT 56.850 23.860 56.880 24.030 ;
        RECT 57.050 23.860 57.240 24.030 ;
        RECT 57.410 23.860 57.600 24.030 ;
        RECT 57.770 23.860 57.800 24.030 ;
        RECT 56.850 23.710 57.800 23.860 ;
        RECT 58.420 24.030 59.360 24.060 ;
        RECT 58.420 23.860 58.440 24.030 ;
        RECT 58.610 23.860 58.800 24.030 ;
        RECT 58.970 23.860 59.160 24.030 ;
        RECT 59.330 23.860 59.360 24.030 ;
        RECT 56.500 23.530 56.670 23.610 ;
        RECT 56.500 23.360 57.680 23.530 ;
        RECT 56.530 23.030 56.860 23.180 ;
        RECT 56.530 22.840 57.330 23.030 ;
        RECT 54.610 22.670 57.330 22.840 ;
        RECT 53.400 21.900 53.910 22.060 ;
        RECT 54.610 21.830 54.780 22.670 ;
        RECT 55.430 22.180 55.760 22.490 ;
        RECT 57.000 22.360 57.330 22.670 ;
        RECT 57.510 22.180 57.680 23.360 ;
        RECT 55.430 22.010 57.680 22.180 ;
        RECT 57.990 22.750 58.240 23.720 ;
        RECT 58.420 22.930 59.360 23.860 ;
        RECT 57.990 22.580 59.360 22.750 ;
        RECT 55.430 21.900 55.760 22.010 ;
        RECT 54.150 21.540 54.780 21.830 ;
      LAYER li1 ;
        RECT 56.010 21.360 56.280 21.390 ;
        RECT 53.050 21.190 56.280 21.360 ;
        RECT 53.410 20.910 56.280 21.190 ;
      LAYER li1 ;
        RECT 56.460 20.720 57.050 21.830 ;
        RECT 57.240 21.330 57.570 22.010 ;
        RECT 57.990 21.830 58.200 22.580 ;
        RECT 59.030 22.080 59.360 22.580 ;
        RECT 57.870 21.330 58.200 21.830 ;
        RECT 58.380 20.720 59.330 21.830 ;
      LAYER li1 ;
        RECT 59.540 21.000 59.890 23.970 ;
      LAYER li1 ;
        RECT 60.500 23.910 60.710 24.080 ;
        RECT 60.880 23.910 61.150 24.080 ;
        RECT 61.320 23.910 61.560 24.080 ;
        RECT 61.730 23.910 61.990 24.080 ;
        RECT 62.160 23.910 62.430 24.080 ;
        RECT 62.600 23.910 62.840 24.080 ;
        RECT 63.010 23.910 63.240 24.080 ;
        RECT 60.500 23.030 63.240 23.910 ;
        RECT 64.470 24.030 65.060 24.060 ;
        RECT 64.470 23.860 64.500 24.030 ;
        RECT 64.670 23.860 64.860 24.030 ;
        RECT 65.030 23.860 65.060 24.030 ;
        RECT 60.740 21.710 61.070 22.380 ;
        RECT 61.470 22.050 61.800 23.030 ;
        RECT 62.020 21.710 62.350 22.380 ;
        RECT 62.750 22.050 63.080 23.030 ;
        RECT 63.950 22.880 64.280 23.810 ;
        RECT 64.470 23.080 65.060 23.860 ;
        RECT 65.240 23.990 66.680 24.160 ;
        RECT 65.240 22.880 65.410 23.990 ;
        RECT 63.950 22.710 65.410 22.880 ;
        RECT 60.580 20.710 63.310 21.710 ;
        RECT 63.950 20.850 64.220 22.710 ;
        RECT 65.080 22.210 65.410 22.710 ;
        RECT 65.590 22.500 65.840 23.810 ;
        RECT 66.080 23.190 66.330 23.810 ;
        RECT 66.510 23.540 66.680 23.990 ;
        RECT 66.860 24.030 67.190 24.060 ;
        RECT 66.860 23.860 66.890 24.030 ;
        RECT 67.060 23.860 67.190 24.030 ;
        RECT 66.860 23.720 67.190 23.860 ;
        RECT 67.370 23.990 69.110 24.160 ;
        RECT 67.370 23.540 67.540 23.990 ;
        RECT 66.510 23.370 67.540 23.540 ;
        RECT 67.720 23.190 67.890 23.810 ;
        RECT 68.420 23.550 68.750 23.810 ;
        RECT 66.080 23.020 67.890 23.190 ;
        RECT 68.070 23.020 68.290 23.350 ;
        RECT 67.720 22.840 67.890 23.020 ;
        RECT 65.590 22.270 66.120 22.500 ;
        RECT 65.590 21.350 65.860 22.270 ;
      LAYER li1 ;
        RECT 66.540 21.970 67.080 22.840 ;
      LAYER li1 ;
        RECT 67.720 22.670 67.940 22.840 ;
        RECT 64.400 20.720 65.350 21.350 ;
        RECT 65.530 20.850 65.860 21.350 ;
        RECT 66.040 20.720 66.630 21.600 ;
      LAYER li1 ;
        RECT 66.910 21.360 67.080 21.970 ;
        RECT 66.870 21.190 67.080 21.360 ;
        RECT 66.910 20.980 67.080 21.190 ;
        RECT 67.260 21.160 67.590 22.460 ;
      LAYER li1 ;
        RECT 67.770 21.680 67.940 22.670 ;
        RECT 68.120 22.500 68.290 23.020 ;
        RECT 68.470 22.850 68.640 23.550 ;
        RECT 68.940 23.400 69.110 23.990 ;
        RECT 69.290 24.030 70.240 24.060 ;
        RECT 69.290 23.860 69.320 24.030 ;
        RECT 69.490 23.860 69.680 24.030 ;
        RECT 69.850 23.860 70.040 24.030 ;
        RECT 70.210 23.860 70.240 24.030 ;
        RECT 69.290 23.580 70.240 23.860 ;
        RECT 70.420 23.990 71.450 24.160 ;
        RECT 70.420 23.400 70.590 23.990 ;
        RECT 68.940 23.350 70.590 23.400 ;
        RECT 68.820 23.230 70.590 23.350 ;
        RECT 68.820 23.030 69.150 23.230 ;
        RECT 70.770 23.050 71.100 23.810 ;
        RECT 71.280 23.630 71.450 23.990 ;
        RECT 71.630 24.030 72.580 24.110 ;
        RECT 71.630 23.860 71.660 24.030 ;
        RECT 71.830 23.860 72.020 24.030 ;
        RECT 72.190 23.860 72.380 24.030 ;
        RECT 72.550 23.860 72.580 24.030 ;
        RECT 71.630 23.810 72.580 23.860 ;
        RECT 71.280 23.460 73.090 23.630 ;
        RECT 69.330 22.880 71.100 23.050 ;
        RECT 69.330 22.850 69.500 22.880 ;
        RECT 68.470 22.680 69.500 22.850 ;
        RECT 72.410 22.700 72.740 23.280 ;
        RECT 68.120 22.270 69.150 22.500 ;
        RECT 68.820 21.780 69.150 22.270 ;
        RECT 69.330 22.000 69.500 22.680 ;
        RECT 69.680 22.530 72.740 22.700 ;
        RECT 69.680 22.180 70.010 22.530 ;
      LAYER li1 ;
        RECT 70.450 22.180 72.300 22.350 ;
      LAYER li1 ;
        RECT 69.330 21.830 71.950 22.000 ;
        RECT 67.770 21.180 68.040 21.680 ;
        RECT 69.330 21.600 69.500 21.830 ;
      LAYER li1 ;
        RECT 72.130 21.650 72.300 22.180 ;
      LAYER li1 ;
        RECT 68.490 21.430 69.500 21.600 ;
      LAYER li1 ;
        RECT 69.680 21.480 72.300 21.650 ;
      LAYER li1 ;
        RECT 68.490 21.180 68.820 21.430 ;
      LAYER li1 ;
        RECT 69.680 20.980 69.850 21.480 ;
        RECT 66.910 20.810 69.850 20.980 ;
      LAYER li1 ;
        RECT 71.000 20.720 71.950 21.300 ;
      LAYER li1 ;
        RECT 72.130 20.790 72.300 21.480 ;
      LAYER li1 ;
        RECT 72.480 21.680 72.740 22.530 ;
        RECT 72.920 22.110 73.090 23.460 ;
        RECT 73.270 23.200 73.520 24.110 ;
        RECT 74.330 24.030 75.280 24.060 ;
        RECT 76.110 24.030 77.010 24.060 ;
        RECT 74.330 23.860 74.360 24.030 ;
        RECT 74.530 23.860 74.720 24.030 ;
        RECT 74.890 23.860 75.080 24.030 ;
        RECT 75.250 23.860 75.280 24.030 ;
        RECT 76.280 23.860 76.470 24.030 ;
        RECT 76.640 23.860 76.830 24.030 ;
        RECT 77.000 23.860 77.010 24.030 ;
        RECT 73.270 23.030 74.150 23.200 ;
        RECT 74.330 23.030 75.280 23.860 ;
        RECT 75.680 23.060 75.930 23.530 ;
        RECT 76.110 23.240 77.010 23.860 ;
        RECT 77.620 24.030 78.560 24.090 ;
        RECT 77.620 23.860 77.640 24.030 ;
        RECT 77.810 23.860 78.000 24.030 ;
        RECT 78.170 23.860 78.360 24.030 ;
        RECT 78.530 23.860 78.560 24.030 ;
        RECT 73.470 22.290 73.800 22.790 ;
        RECT 73.980 22.710 74.150 23.030 ;
        RECT 75.680 22.890 76.690 23.060 ;
        RECT 73.980 22.540 76.340 22.710 ;
        RECT 72.920 21.940 74.090 22.110 ;
        RECT 72.480 20.970 72.810 21.680 ;
        RECT 73.270 21.140 73.600 21.680 ;
        RECT 73.810 21.440 74.090 21.940 ;
        RECT 74.270 21.140 74.440 22.540 ;
        RECT 76.520 22.360 76.690 22.890 ;
        RECT 74.650 22.190 76.690 22.360 ;
        RECT 74.650 21.800 74.980 22.190 ;
      LAYER li1 ;
        RECT 75.300 21.620 75.630 22.010 ;
      LAYER li1 ;
        RECT 73.270 20.970 74.440 21.140 ;
      LAYER li1 ;
        RECT 74.620 21.450 75.630 21.620 ;
        RECT 74.620 20.790 74.790 21.450 ;
      LAYER li1 ;
        RECT 76.460 21.350 76.690 22.190 ;
        RECT 77.190 22.360 77.440 23.360 ;
        RECT 77.620 22.550 78.560 23.860 ;
        RECT 77.190 22.030 78.560 22.360 ;
        RECT 77.190 21.850 77.400 22.030 ;
        RECT 77.070 21.350 77.400 21.850 ;
      LAYER li1 ;
        RECT 72.130 20.620 74.790 20.790 ;
      LAYER li1 ;
        RECT 74.970 20.720 75.920 21.270 ;
        RECT 76.460 20.850 76.790 21.350 ;
        RECT 77.580 20.720 78.530 21.850 ;
      LAYER li1 ;
        RECT 78.740 21.020 79.080 24.090 ;
      LAYER li1 ;
        RECT 79.450 24.080 80.900 24.110 ;
        RECT 79.450 23.910 79.700 24.080 ;
        RECT 79.870 23.910 80.060 24.080 ;
        RECT 80.230 23.910 80.500 24.080 ;
        RECT 80.670 23.910 80.900 24.080 ;
        RECT 79.450 23.040 80.900 23.910 ;
        RECT 79.680 21.600 80.010 22.380 ;
        RECT 80.220 22.050 80.550 23.040 ;
      LAYER li1 ;
        RECT 81.240 22.530 81.670 24.110 ;
      LAYER li1 ;
        RECT 81.850 24.030 82.410 24.110 ;
        RECT 81.850 23.860 81.860 24.030 ;
        RECT 82.030 23.860 82.220 24.030 ;
        RECT 82.390 23.860 82.410 24.030 ;
        RECT 81.850 22.530 82.410 23.860 ;
        RECT 83.770 24.080 85.220 24.110 ;
        RECT 83.770 23.910 84.020 24.080 ;
        RECT 84.190 23.910 84.380 24.080 ;
        RECT 84.550 23.910 84.820 24.080 ;
        RECT 84.990 23.910 85.220 24.080 ;
        RECT 79.680 21.200 80.980 21.600 ;
        RECT 79.370 20.720 80.980 21.200 ;
      LAYER li1 ;
        RECT 81.240 20.850 81.490 22.530 ;
      LAYER li1 ;
        RECT 81.800 21.640 82.130 22.100 ;
      LAYER li1 ;
        RECT 82.590 21.820 82.920 23.610 ;
      LAYER li1 ;
        RECT 83.100 21.640 83.350 23.360 ;
        RECT 83.770 23.040 85.220 23.910 ;
        RECT 81.800 21.470 83.350 21.640 ;
        RECT 81.670 20.720 82.920 21.290 ;
        RECT 83.100 20.850 83.350 21.470 ;
        RECT 84.000 21.600 84.330 22.380 ;
        RECT 84.540 22.050 84.870 23.040 ;
      LAYER li1 ;
        RECT 85.560 22.530 85.990 24.110 ;
      LAYER li1 ;
        RECT 86.170 24.030 86.730 24.110 ;
        RECT 86.170 23.860 86.180 24.030 ;
        RECT 86.350 23.860 86.540 24.030 ;
        RECT 86.710 23.860 86.730 24.030 ;
        RECT 86.170 22.530 86.730 23.860 ;
        RECT 88.090 24.080 89.540 24.110 ;
        RECT 88.090 23.910 88.340 24.080 ;
        RECT 88.510 23.910 88.700 24.080 ;
        RECT 88.870 23.910 89.140 24.080 ;
        RECT 89.310 23.910 89.540 24.080 ;
        RECT 84.000 21.200 85.300 21.600 ;
        RECT 83.690 20.720 85.300 21.200 ;
      LAYER li1 ;
        RECT 85.560 20.850 85.810 22.530 ;
      LAYER li1 ;
        RECT 86.120 21.640 86.450 22.100 ;
      LAYER li1 ;
        RECT 86.910 21.820 87.240 23.610 ;
      LAYER li1 ;
        RECT 87.420 21.640 87.670 23.360 ;
        RECT 88.090 23.040 89.540 23.910 ;
        RECT 90.810 24.030 92.480 24.110 ;
        RECT 90.810 23.860 90.840 24.030 ;
        RECT 91.010 23.860 91.200 24.030 ;
        RECT 91.370 23.860 91.560 24.030 ;
        RECT 91.730 23.860 91.920 24.030 ;
        RECT 92.090 23.860 92.280 24.030 ;
        RECT 92.450 23.860 92.480 24.030 ;
        RECT 86.120 21.470 87.670 21.640 ;
        RECT 85.990 20.720 87.240 21.290 ;
        RECT 87.420 20.850 87.670 21.470 ;
        RECT 88.320 21.600 88.650 22.380 ;
        RECT 88.860 22.050 89.190 23.040 ;
        RECT 90.810 22.650 92.480 23.860 ;
      LAYER li1 ;
        RECT 90.850 22.130 92.040 22.470 ;
        RECT 92.220 22.130 92.550 22.470 ;
        RECT 92.740 21.950 93.000 24.110 ;
      LAYER li1 ;
        RECT 93.370 24.080 94.820 24.110 ;
        RECT 93.370 23.910 93.620 24.080 ;
        RECT 93.790 23.910 93.980 24.080 ;
        RECT 94.150 23.910 94.420 24.080 ;
        RECT 94.590 23.910 94.820 24.080 ;
        RECT 93.370 23.040 94.820 23.910 ;
      LAYER li1 ;
        RECT 91.920 21.780 93.000 21.950 ;
      LAYER li1 ;
        RECT 88.320 21.200 89.620 21.600 ;
        RECT 88.010 20.720 89.620 21.200 ;
        RECT 90.810 20.720 91.740 21.680 ;
      LAYER li1 ;
        RECT 91.920 20.850 92.250 21.780 ;
      LAYER li1 ;
        RECT 93.600 21.600 93.930 22.380 ;
        RECT 94.140 22.050 94.470 23.040 ;
      LAYER li1 ;
        RECT 95.160 22.530 95.590 24.110 ;
      LAYER li1 ;
        RECT 95.770 24.030 96.330 24.110 ;
        RECT 95.770 23.860 95.780 24.030 ;
        RECT 95.950 23.860 96.140 24.030 ;
        RECT 96.310 23.860 96.330 24.030 ;
        RECT 95.770 22.530 96.330 23.860 ;
        RECT 97.690 24.080 99.140 24.110 ;
        RECT 97.690 23.910 97.940 24.080 ;
        RECT 98.110 23.910 98.300 24.080 ;
        RECT 98.470 23.910 98.740 24.080 ;
        RECT 98.910 23.910 99.140 24.080 ;
        RECT 92.440 20.720 93.030 21.600 ;
        RECT 93.600 21.200 94.900 21.600 ;
        RECT 93.290 20.720 94.900 21.200 ;
      LAYER li1 ;
        RECT 95.160 20.850 95.410 22.530 ;
      LAYER li1 ;
        RECT 95.720 21.640 96.050 22.100 ;
      LAYER li1 ;
        RECT 96.510 21.820 96.840 23.610 ;
      LAYER li1 ;
        RECT 97.020 21.640 97.270 23.360 ;
        RECT 97.690 23.040 99.140 23.910 ;
        RECT 99.450 24.030 100.400 24.110 ;
        RECT 99.450 23.860 99.480 24.030 ;
        RECT 99.650 23.860 99.840 24.030 ;
        RECT 100.010 23.860 100.200 24.030 ;
        RECT 100.370 23.860 100.400 24.030 ;
        RECT 95.720 21.470 97.270 21.640 ;
        RECT 95.590 20.720 96.840 21.290 ;
        RECT 97.020 20.850 97.270 21.470 ;
        RECT 97.920 21.600 98.250 22.380 ;
        RECT 98.460 22.050 98.790 23.040 ;
      LAYER li1 ;
        RECT 99.030 21.930 99.200 22.840 ;
      LAYER li1 ;
        RECT 99.450 22.530 100.400 23.860 ;
      LAYER li1 ;
        RECT 99.490 21.900 100.380 22.290 ;
        RECT 100.580 22.050 100.830 24.110 ;
      LAYER li1 ;
        RECT 101.020 24.030 101.610 24.110 ;
        RECT 101.020 23.860 101.050 24.030 ;
        RECT 101.220 23.860 101.410 24.030 ;
        RECT 101.580 23.860 101.610 24.030 ;
        RECT 101.020 22.530 101.610 23.860 ;
        RECT 102.010 24.080 103.460 24.110 ;
        RECT 102.010 23.910 102.260 24.080 ;
        RECT 102.430 23.910 102.620 24.080 ;
        RECT 102.790 23.910 103.060 24.080 ;
        RECT 103.230 23.910 103.460 24.080 ;
        RECT 102.010 23.040 103.460 23.910 ;
        RECT 103.770 24.030 104.720 24.110 ;
        RECT 103.770 23.860 103.800 24.030 ;
        RECT 103.970 23.860 104.160 24.030 ;
        RECT 104.330 23.860 104.520 24.030 ;
        RECT 104.690 23.860 104.720 24.030 ;
      LAYER li1 ;
        RECT 100.580 21.880 101.160 22.050 ;
        RECT 101.340 21.880 101.640 22.210 ;
        RECT 100.940 21.700 101.160 21.880 ;
      LAYER li1 ;
        RECT 97.920 21.200 99.220 21.600 ;
        RECT 97.610 20.720 99.220 21.200 ;
        RECT 99.450 20.720 100.760 21.700 ;
      LAYER li1 ;
        RECT 100.940 21.530 101.540 21.700 ;
        RECT 101.210 20.870 101.540 21.530 ;
      LAYER li1 ;
        RECT 102.240 21.600 102.570 22.380 ;
        RECT 102.780 22.050 103.110 23.040 ;
        RECT 103.770 22.530 104.720 23.860 ;
      LAYER li1 ;
        RECT 103.810 21.900 104.700 22.290 ;
        RECT 104.900 22.050 105.150 24.110 ;
      LAYER li1 ;
        RECT 105.340 24.030 105.930 24.110 ;
        RECT 105.340 23.860 105.370 24.030 ;
        RECT 105.540 23.860 105.730 24.030 ;
        RECT 105.900 23.860 105.930 24.030 ;
        RECT 105.340 22.530 105.930 23.860 ;
        RECT 106.330 24.080 107.780 24.110 ;
        RECT 106.330 23.910 106.580 24.080 ;
        RECT 106.750 23.910 106.940 24.080 ;
        RECT 107.110 23.910 107.380 24.080 ;
        RECT 107.550 23.910 107.780 24.080 ;
        RECT 106.330 23.040 107.780 23.910 ;
      LAYER li1 ;
        RECT 104.900 21.880 105.480 22.050 ;
        RECT 105.660 21.880 105.960 22.210 ;
        RECT 105.260 21.700 105.480 21.880 ;
      LAYER li1 ;
        RECT 102.240 21.200 103.540 21.600 ;
        RECT 101.930 20.720 103.540 21.200 ;
        RECT 103.770 20.720 105.080 21.700 ;
      LAYER li1 ;
        RECT 105.260 21.530 105.860 21.700 ;
        RECT 105.530 20.870 105.860 21.530 ;
      LAYER li1 ;
        RECT 106.560 21.600 106.890 22.380 ;
        RECT 107.100 22.050 107.430 23.040 ;
      LAYER li1 ;
        RECT 108.630 21.930 108.800 22.840 ;
        RECT 109.080 22.530 109.510 24.110 ;
      LAYER li1 ;
        RECT 109.690 24.030 110.250 24.110 ;
        RECT 109.690 23.860 109.700 24.030 ;
        RECT 109.870 23.860 110.060 24.030 ;
        RECT 110.230 23.860 110.250 24.030 ;
        RECT 109.690 22.530 110.250 23.860 ;
        RECT 111.610 24.080 113.060 24.110 ;
        RECT 111.610 23.910 111.860 24.080 ;
        RECT 112.030 23.910 112.220 24.080 ;
        RECT 112.390 23.910 112.660 24.080 ;
        RECT 112.830 23.910 113.060 24.080 ;
        RECT 106.560 21.200 107.860 21.600 ;
        RECT 106.250 20.720 107.860 21.200 ;
      LAYER li1 ;
        RECT 109.080 20.850 109.330 22.530 ;
      LAYER li1 ;
        RECT 109.640 21.640 109.970 22.100 ;
      LAYER li1 ;
        RECT 110.430 21.820 110.760 23.610 ;
      LAYER li1 ;
        RECT 110.940 21.640 111.190 23.360 ;
        RECT 111.610 23.040 113.060 23.910 ;
        RECT 113.370 24.030 115.040 24.110 ;
        RECT 113.370 23.860 113.400 24.030 ;
        RECT 113.570 23.860 113.760 24.030 ;
        RECT 113.930 23.860 114.120 24.030 ;
        RECT 114.290 23.860 114.480 24.030 ;
        RECT 114.650 23.860 114.840 24.030 ;
        RECT 115.010 23.860 115.040 24.030 ;
        RECT 109.640 21.470 111.190 21.640 ;
        RECT 109.510 20.720 110.760 21.290 ;
        RECT 110.940 20.850 111.190 21.470 ;
        RECT 111.840 21.600 112.170 22.380 ;
        RECT 112.380 22.050 112.710 23.040 ;
        RECT 113.370 22.650 115.040 23.860 ;
      LAYER li1 ;
        RECT 113.410 22.130 114.600 22.470 ;
        RECT 114.780 22.130 115.110 22.470 ;
        RECT 115.300 21.950 115.560 24.110 ;
      LAYER li1 ;
        RECT 115.930 24.080 117.380 24.110 ;
        RECT 115.930 23.910 116.180 24.080 ;
        RECT 116.350 23.910 116.540 24.080 ;
        RECT 116.710 23.910 116.980 24.080 ;
        RECT 117.150 23.910 117.380 24.080 ;
        RECT 115.930 23.040 117.380 23.910 ;
        RECT 117.690 24.030 119.360 24.110 ;
        RECT 117.690 23.860 117.720 24.030 ;
        RECT 117.890 23.860 118.080 24.030 ;
        RECT 118.250 23.860 118.440 24.030 ;
        RECT 118.610 23.860 118.800 24.030 ;
        RECT 118.970 23.860 119.160 24.030 ;
        RECT 119.330 23.860 119.360 24.030 ;
      LAYER li1 ;
        RECT 114.480 21.780 115.560 21.950 ;
      LAYER li1 ;
        RECT 111.840 21.200 113.140 21.600 ;
        RECT 111.530 20.720 113.140 21.200 ;
        RECT 113.370 20.720 114.300 21.680 ;
      LAYER li1 ;
        RECT 114.480 20.850 114.810 21.780 ;
      LAYER li1 ;
        RECT 116.160 21.600 116.490 22.380 ;
        RECT 116.700 22.050 117.030 23.040 ;
        RECT 117.690 22.650 119.360 23.860 ;
      LAYER li1 ;
        RECT 117.730 22.130 118.920 22.470 ;
        RECT 119.100 22.130 119.430 22.470 ;
        RECT 119.620 21.950 119.880 24.110 ;
      LAYER li1 ;
        RECT 120.250 24.080 121.700 24.110 ;
        RECT 120.250 23.910 120.500 24.080 ;
        RECT 120.670 23.910 120.860 24.080 ;
        RECT 121.030 23.910 121.300 24.080 ;
        RECT 121.470 23.910 121.700 24.080 ;
        RECT 120.250 23.040 121.700 23.910 ;
        RECT 122.550 24.030 123.140 24.060 ;
        RECT 122.550 23.860 122.580 24.030 ;
        RECT 122.750 23.860 122.940 24.030 ;
        RECT 123.110 23.860 123.140 24.030 ;
      LAYER li1 ;
        RECT 118.800 21.780 119.880 21.950 ;
      LAYER li1 ;
        RECT 115.000 20.720 115.590 21.600 ;
        RECT 116.160 21.200 117.460 21.600 ;
        RECT 115.850 20.720 117.460 21.200 ;
        RECT 117.690 20.720 118.620 21.680 ;
      LAYER li1 ;
        RECT 118.800 20.850 119.130 21.780 ;
      LAYER li1 ;
        RECT 120.480 21.600 120.810 22.380 ;
        RECT 121.020 22.050 121.350 23.040 ;
        RECT 122.030 22.880 122.360 23.810 ;
        RECT 122.550 23.080 123.140 23.860 ;
        RECT 123.320 23.990 124.760 24.160 ;
        RECT 123.320 22.880 123.490 23.990 ;
        RECT 122.030 22.710 123.490 22.880 ;
        RECT 119.320 20.720 119.910 21.600 ;
        RECT 120.480 21.200 121.780 21.600 ;
        RECT 120.170 20.720 121.780 21.200 ;
        RECT 122.030 20.850 122.300 22.710 ;
        RECT 123.160 22.210 123.490 22.710 ;
        RECT 123.670 22.500 123.920 23.810 ;
        RECT 124.160 23.190 124.410 23.810 ;
        RECT 124.590 23.540 124.760 23.990 ;
        RECT 124.940 24.030 125.270 24.060 ;
        RECT 124.940 23.860 124.970 24.030 ;
        RECT 125.140 23.860 125.270 24.030 ;
        RECT 124.940 23.720 125.270 23.860 ;
        RECT 125.450 23.990 127.190 24.160 ;
        RECT 125.450 23.540 125.620 23.990 ;
        RECT 124.590 23.370 125.620 23.540 ;
        RECT 125.800 23.190 125.970 23.810 ;
        RECT 126.500 23.550 126.830 23.810 ;
        RECT 124.160 23.020 125.970 23.190 ;
        RECT 126.150 23.020 126.370 23.350 ;
        RECT 125.800 22.840 125.970 23.020 ;
        RECT 123.670 22.270 124.200 22.500 ;
        RECT 123.670 21.350 123.940 22.270 ;
      LAYER li1 ;
        RECT 124.620 21.970 125.160 22.840 ;
      LAYER li1 ;
        RECT 125.800 22.670 126.020 22.840 ;
        RECT 122.480 20.720 123.430 21.350 ;
        RECT 123.610 20.850 123.940 21.350 ;
        RECT 124.120 20.720 124.710 21.600 ;
      LAYER li1 ;
        RECT 124.990 20.980 125.160 21.970 ;
        RECT 125.340 21.160 125.670 22.460 ;
      LAYER li1 ;
        RECT 125.850 21.680 126.020 22.670 ;
        RECT 126.200 22.500 126.370 23.020 ;
        RECT 126.550 22.850 126.720 23.550 ;
        RECT 127.020 23.400 127.190 23.990 ;
        RECT 127.370 24.030 128.320 24.060 ;
        RECT 127.370 23.860 127.400 24.030 ;
        RECT 127.570 23.860 127.760 24.030 ;
        RECT 127.930 23.860 128.120 24.030 ;
        RECT 128.290 23.860 128.320 24.030 ;
        RECT 127.370 23.580 128.320 23.860 ;
        RECT 128.500 23.990 129.530 24.160 ;
        RECT 128.500 23.400 128.670 23.990 ;
        RECT 127.020 23.350 128.670 23.400 ;
        RECT 126.900 23.230 128.670 23.350 ;
        RECT 126.900 23.030 127.230 23.230 ;
        RECT 128.850 23.050 129.180 23.810 ;
        RECT 129.360 23.630 129.530 23.990 ;
        RECT 129.710 24.030 130.660 24.110 ;
        RECT 129.710 23.860 129.740 24.030 ;
        RECT 129.910 23.860 130.100 24.030 ;
        RECT 130.270 23.860 130.460 24.030 ;
        RECT 130.630 23.860 130.660 24.030 ;
        RECT 129.710 23.810 130.660 23.860 ;
        RECT 129.360 23.460 131.170 23.630 ;
        RECT 127.410 22.880 129.180 23.050 ;
        RECT 127.410 22.850 127.580 22.880 ;
        RECT 126.550 22.680 127.580 22.850 ;
        RECT 130.490 22.700 130.820 23.280 ;
        RECT 126.200 22.270 127.230 22.500 ;
        RECT 126.900 21.780 127.230 22.270 ;
        RECT 127.410 22.000 127.580 22.680 ;
        RECT 127.760 22.530 130.820 22.700 ;
        RECT 127.760 22.180 128.090 22.530 ;
      LAYER li1 ;
        RECT 128.530 22.180 130.380 22.350 ;
      LAYER li1 ;
        RECT 127.410 21.830 130.030 22.000 ;
        RECT 125.850 21.180 126.120 21.680 ;
        RECT 127.410 21.600 127.580 21.830 ;
      LAYER li1 ;
        RECT 130.210 21.650 130.380 22.180 ;
      LAYER li1 ;
        RECT 126.570 21.430 127.580 21.600 ;
      LAYER li1 ;
        RECT 127.760 21.480 130.380 21.650 ;
      LAYER li1 ;
        RECT 126.570 21.180 126.900 21.430 ;
      LAYER li1 ;
        RECT 127.760 20.980 127.930 21.480 ;
        RECT 124.990 20.810 127.930 20.980 ;
      LAYER li1 ;
        RECT 129.080 20.720 130.030 21.300 ;
      LAYER li1 ;
        RECT 130.210 20.790 130.380 21.480 ;
      LAYER li1 ;
        RECT 130.560 21.680 130.820 22.530 ;
        RECT 131.000 22.110 131.170 23.460 ;
        RECT 131.350 23.200 131.600 24.110 ;
        RECT 132.410 24.030 133.360 24.060 ;
        RECT 134.190 24.030 135.090 24.060 ;
        RECT 132.410 23.860 132.440 24.030 ;
        RECT 132.610 23.860 132.800 24.030 ;
        RECT 132.970 23.860 133.160 24.030 ;
        RECT 133.330 23.860 133.360 24.030 ;
        RECT 134.360 23.860 134.550 24.030 ;
        RECT 134.720 23.860 134.910 24.030 ;
        RECT 135.080 23.860 135.090 24.030 ;
        RECT 131.350 23.030 132.230 23.200 ;
        RECT 132.410 23.030 133.360 23.860 ;
        RECT 133.760 23.060 134.010 23.530 ;
        RECT 134.190 23.240 135.090 23.860 ;
        RECT 135.700 24.030 136.640 24.090 ;
        RECT 135.700 23.860 135.720 24.030 ;
        RECT 135.890 23.860 136.080 24.030 ;
        RECT 136.250 23.860 136.440 24.030 ;
        RECT 136.610 23.860 136.640 24.030 ;
        RECT 131.550 22.290 131.880 22.790 ;
        RECT 132.060 22.710 132.230 23.030 ;
        RECT 133.760 22.890 134.770 23.060 ;
        RECT 132.060 22.540 134.420 22.710 ;
        RECT 131.000 21.940 132.170 22.110 ;
        RECT 130.560 20.970 130.890 21.680 ;
        RECT 131.350 21.140 131.680 21.680 ;
        RECT 131.890 21.440 132.170 21.940 ;
        RECT 132.350 21.140 132.520 22.540 ;
        RECT 134.600 22.360 134.770 22.890 ;
        RECT 132.730 22.190 134.770 22.360 ;
        RECT 132.730 21.800 133.060 22.190 ;
      LAYER li1 ;
        RECT 133.380 21.620 133.710 22.010 ;
      LAYER li1 ;
        RECT 131.350 20.970 132.520 21.140 ;
      LAYER li1 ;
        RECT 132.700 21.450 133.710 21.620 ;
        RECT 132.700 20.790 132.870 21.450 ;
      LAYER li1 ;
        RECT 134.540 21.350 134.770 22.190 ;
        RECT 135.270 22.360 135.520 23.360 ;
        RECT 135.700 22.550 136.640 23.860 ;
        RECT 135.270 22.030 136.640 22.360 ;
        RECT 135.270 21.850 135.480 22.030 ;
        RECT 135.150 21.350 135.480 21.850 ;
      LAYER li1 ;
        RECT 130.210 20.620 132.870 20.790 ;
      LAYER li1 ;
        RECT 133.050 20.720 134.000 21.270 ;
        RECT 134.540 20.850 134.870 21.350 ;
        RECT 135.660 20.720 136.610 21.850 ;
      LAYER li1 ;
        RECT 136.820 21.020 137.160 24.090 ;
      LAYER li1 ;
        RECT 137.780 24.080 140.520 24.100 ;
        RECT 137.780 23.910 137.990 24.080 ;
        RECT 138.160 23.910 138.430 24.080 ;
        RECT 138.600 23.910 138.840 24.080 ;
        RECT 139.010 23.910 139.270 24.080 ;
        RECT 139.440 23.910 139.710 24.080 ;
        RECT 139.880 23.910 140.120 24.080 ;
        RECT 140.290 23.910 140.520 24.080 ;
        RECT 137.780 23.030 140.520 23.910 ;
        RECT 138.020 21.710 138.350 22.380 ;
        RECT 138.750 22.050 139.080 23.030 ;
        RECT 139.300 21.710 139.630 22.380 ;
        RECT 140.030 22.050 140.360 23.030 ;
        RECT 137.860 20.710 140.590 21.710 ;
        RECT 5.760 20.260 5.920 20.440 ;
        RECT 6.090 20.260 6.400 20.440 ;
        RECT 6.570 20.260 6.880 20.440 ;
        RECT 7.050 20.260 7.360 20.440 ;
        RECT 7.530 20.260 7.840 20.440 ;
        RECT 8.010 20.260 8.320 20.440 ;
        RECT 8.490 20.260 8.800 20.440 ;
        RECT 8.970 20.260 9.280 20.440 ;
        RECT 9.450 20.260 9.760 20.440 ;
        RECT 9.930 20.260 10.240 20.440 ;
        RECT 10.410 20.260 10.720 20.440 ;
        RECT 10.890 20.260 11.200 20.440 ;
        RECT 11.370 20.260 11.680 20.440 ;
        RECT 11.850 20.260 12.160 20.440 ;
        RECT 12.330 20.260 12.640 20.440 ;
        RECT 12.810 20.260 13.120 20.440 ;
        RECT 13.290 20.260 13.600 20.440 ;
        RECT 13.770 20.260 14.080 20.440 ;
        RECT 14.250 20.260 14.560 20.440 ;
        RECT 14.730 20.260 15.040 20.440 ;
        RECT 15.210 20.260 15.520 20.440 ;
        RECT 15.690 20.260 16.000 20.440 ;
        RECT 16.170 20.260 16.480 20.440 ;
        RECT 16.650 20.260 16.960 20.440 ;
        RECT 17.130 20.260 17.440 20.440 ;
        RECT 17.610 20.260 17.920 20.440 ;
        RECT 18.090 20.260 18.400 20.440 ;
        RECT 18.570 20.260 18.880 20.440 ;
        RECT 19.050 20.260 19.360 20.440 ;
        RECT 19.530 20.260 19.840 20.440 ;
        RECT 20.010 20.260 20.320 20.440 ;
        RECT 20.490 20.260 20.800 20.440 ;
        RECT 20.970 20.260 21.280 20.440 ;
        RECT 21.450 20.260 21.760 20.440 ;
        RECT 21.930 20.260 22.240 20.440 ;
        RECT 22.410 20.260 22.720 20.440 ;
        RECT 22.890 20.260 23.200 20.440 ;
        RECT 23.370 20.260 23.680 20.440 ;
        RECT 23.850 20.260 24.160 20.440 ;
        RECT 24.330 20.260 24.640 20.440 ;
        RECT 24.810 20.260 25.120 20.440 ;
        RECT 25.290 20.260 25.600 20.440 ;
        RECT 25.770 20.260 26.080 20.440 ;
        RECT 26.250 20.260 26.560 20.440 ;
        RECT 26.730 20.260 27.040 20.440 ;
        RECT 27.210 20.260 27.520 20.440 ;
        RECT 27.690 20.260 28.000 20.440 ;
        RECT 28.170 20.260 28.480 20.440 ;
        RECT 28.650 20.260 28.960 20.440 ;
        RECT 29.130 20.260 29.440 20.440 ;
        RECT 29.610 20.260 29.920 20.440 ;
        RECT 30.090 20.260 30.400 20.440 ;
        RECT 30.570 20.260 30.880 20.440 ;
        RECT 31.050 20.260 31.360 20.440 ;
        RECT 31.530 20.260 31.840 20.440 ;
        RECT 32.010 20.260 32.320 20.440 ;
        RECT 32.490 20.260 32.800 20.440 ;
        RECT 32.970 20.260 33.280 20.440 ;
        RECT 33.450 20.260 33.760 20.440 ;
        RECT 33.930 20.260 34.240 20.440 ;
        RECT 34.410 20.260 34.720 20.440 ;
        RECT 34.890 20.260 35.200 20.440 ;
        RECT 35.370 20.260 35.680 20.440 ;
        RECT 35.850 20.260 36.160 20.440 ;
        RECT 36.330 20.260 36.640 20.440 ;
        RECT 36.810 20.260 37.120 20.440 ;
        RECT 37.290 20.260 37.600 20.440 ;
        RECT 37.770 20.260 38.080 20.440 ;
        RECT 38.250 20.260 38.560 20.440 ;
        RECT 38.730 20.260 39.040 20.440 ;
        RECT 39.210 20.260 39.520 20.440 ;
        RECT 39.690 20.260 40.000 20.440 ;
        RECT 40.170 20.260 40.480 20.440 ;
        RECT 40.650 20.260 40.960 20.440 ;
        RECT 41.130 20.260 41.440 20.440 ;
        RECT 41.610 20.260 41.920 20.440 ;
        RECT 42.090 20.260 42.400 20.440 ;
        RECT 42.570 20.260 42.880 20.440 ;
        RECT 43.050 20.260 43.360 20.440 ;
        RECT 43.530 20.260 43.840 20.440 ;
        RECT 44.010 20.260 44.320 20.440 ;
        RECT 44.490 20.260 44.800 20.440 ;
        RECT 44.970 20.260 45.280 20.440 ;
        RECT 45.450 20.260 45.760 20.440 ;
        RECT 45.930 20.260 46.240 20.440 ;
        RECT 46.410 20.260 46.720 20.440 ;
        RECT 46.890 20.260 47.200 20.440 ;
        RECT 47.370 20.260 47.680 20.440 ;
        RECT 47.850 20.260 48.160 20.440 ;
        RECT 48.330 20.260 48.640 20.440 ;
        RECT 48.810 20.260 49.120 20.440 ;
        RECT 49.290 20.260 49.600 20.440 ;
        RECT 49.770 20.260 50.080 20.440 ;
        RECT 50.250 20.260 50.560 20.440 ;
        RECT 50.730 20.260 51.040 20.440 ;
        RECT 51.210 20.260 51.520 20.440 ;
        RECT 51.690 20.260 52.000 20.440 ;
        RECT 52.170 20.260 52.480 20.440 ;
        RECT 52.650 20.260 52.960 20.440 ;
        RECT 53.130 20.260 53.440 20.440 ;
        RECT 53.610 20.260 53.920 20.440 ;
        RECT 54.090 20.260 54.400 20.440 ;
        RECT 54.570 20.260 54.880 20.440 ;
        RECT 55.050 20.260 55.360 20.440 ;
        RECT 55.530 20.260 55.840 20.440 ;
        RECT 56.010 20.260 56.320 20.440 ;
        RECT 56.490 20.260 56.800 20.440 ;
        RECT 56.970 20.260 57.280 20.440 ;
        RECT 57.450 20.260 57.760 20.440 ;
        RECT 57.930 20.260 58.240 20.440 ;
        RECT 58.410 20.260 58.720 20.440 ;
        RECT 58.890 20.260 59.200 20.440 ;
        RECT 59.370 20.260 59.680 20.440 ;
        RECT 59.850 20.260 60.160 20.440 ;
        RECT 60.330 20.260 60.640 20.440 ;
        RECT 60.810 20.260 61.120 20.440 ;
        RECT 61.290 20.260 61.600 20.440 ;
        RECT 61.770 20.260 62.080 20.440 ;
        RECT 62.250 20.260 62.560 20.440 ;
        RECT 62.730 20.260 63.040 20.440 ;
        RECT 63.210 20.260 63.520 20.440 ;
        RECT 63.690 20.260 64.000 20.440 ;
        RECT 64.170 20.260 64.480 20.440 ;
        RECT 64.650 20.260 64.960 20.440 ;
        RECT 65.130 20.260 65.440 20.440 ;
        RECT 65.610 20.260 65.920 20.440 ;
        RECT 66.090 20.260 66.400 20.440 ;
        RECT 66.570 20.260 66.880 20.440 ;
        RECT 67.050 20.260 67.360 20.440 ;
        RECT 67.530 20.260 67.840 20.440 ;
        RECT 68.010 20.260 68.320 20.440 ;
        RECT 68.490 20.260 68.800 20.440 ;
        RECT 68.970 20.260 69.280 20.440 ;
        RECT 69.450 20.260 69.760 20.440 ;
        RECT 69.930 20.260 70.240 20.440 ;
        RECT 70.410 20.260 70.720 20.440 ;
        RECT 70.890 20.260 71.200 20.440 ;
        RECT 71.370 20.260 71.680 20.440 ;
        RECT 71.850 20.260 72.160 20.440 ;
        RECT 72.330 20.260 72.640 20.440 ;
        RECT 72.810 20.260 73.120 20.440 ;
        RECT 73.290 20.260 73.600 20.440 ;
        RECT 73.770 20.260 74.080 20.440 ;
        RECT 74.250 20.260 74.560 20.440 ;
        RECT 74.730 20.260 75.040 20.440 ;
        RECT 75.210 20.260 75.520 20.440 ;
        RECT 75.690 20.260 76.000 20.440 ;
        RECT 76.170 20.260 76.480 20.440 ;
        RECT 76.650 20.260 76.960 20.440 ;
        RECT 77.130 20.260 77.440 20.440 ;
        RECT 77.610 20.260 77.920 20.440 ;
        RECT 78.090 20.260 78.400 20.440 ;
        RECT 78.570 20.260 78.880 20.440 ;
        RECT 79.050 20.260 79.360 20.440 ;
        RECT 79.530 20.260 79.840 20.440 ;
        RECT 80.010 20.260 80.320 20.440 ;
        RECT 80.490 20.260 80.800 20.440 ;
        RECT 80.970 20.260 81.280 20.440 ;
        RECT 81.450 20.260 81.760 20.440 ;
        RECT 81.930 20.260 82.240 20.440 ;
        RECT 82.410 20.260 82.720 20.440 ;
        RECT 82.890 20.260 83.200 20.440 ;
        RECT 83.370 20.260 83.680 20.440 ;
        RECT 83.850 20.260 84.160 20.440 ;
        RECT 84.330 20.260 84.640 20.440 ;
        RECT 84.810 20.260 85.120 20.440 ;
        RECT 85.290 20.260 85.600 20.440 ;
        RECT 85.770 20.260 86.080 20.440 ;
        RECT 86.250 20.260 86.560 20.440 ;
        RECT 86.730 20.260 87.040 20.440 ;
        RECT 87.210 20.260 87.520 20.440 ;
        RECT 87.690 20.260 88.000 20.440 ;
        RECT 88.170 20.260 88.480 20.440 ;
        RECT 88.650 20.260 88.960 20.440 ;
        RECT 89.130 20.260 89.440 20.440 ;
        RECT 89.610 20.260 89.920 20.440 ;
        RECT 90.090 20.260 90.400 20.440 ;
        RECT 90.570 20.260 90.880 20.440 ;
        RECT 91.050 20.260 91.360 20.440 ;
        RECT 91.530 20.260 91.840 20.440 ;
        RECT 92.010 20.260 92.320 20.440 ;
        RECT 92.490 20.260 92.800 20.440 ;
        RECT 92.970 20.260 93.280 20.440 ;
        RECT 93.450 20.260 93.760 20.440 ;
        RECT 93.930 20.260 94.240 20.440 ;
        RECT 94.410 20.260 94.720 20.440 ;
        RECT 94.890 20.260 95.200 20.440 ;
        RECT 95.370 20.260 95.680 20.440 ;
        RECT 95.850 20.260 96.160 20.440 ;
        RECT 96.330 20.260 96.640 20.440 ;
        RECT 96.810 20.260 97.120 20.440 ;
        RECT 97.290 20.260 97.600 20.440 ;
        RECT 97.770 20.260 98.080 20.440 ;
        RECT 98.250 20.260 98.560 20.440 ;
        RECT 98.730 20.260 99.040 20.440 ;
        RECT 99.210 20.260 99.520 20.440 ;
        RECT 99.690 20.260 100.000 20.440 ;
        RECT 100.170 20.260 100.480 20.440 ;
        RECT 100.650 20.260 100.960 20.440 ;
        RECT 101.130 20.260 101.440 20.440 ;
        RECT 101.610 20.260 101.920 20.440 ;
        RECT 102.090 20.260 102.400 20.440 ;
        RECT 102.570 20.260 102.880 20.440 ;
        RECT 103.050 20.260 103.360 20.440 ;
        RECT 103.530 20.260 103.840 20.440 ;
        RECT 104.010 20.260 104.320 20.440 ;
        RECT 104.490 20.260 104.800 20.440 ;
        RECT 104.970 20.260 105.280 20.440 ;
        RECT 105.450 20.260 105.760 20.440 ;
        RECT 105.930 20.260 106.240 20.440 ;
        RECT 106.410 20.260 106.720 20.440 ;
        RECT 106.890 20.260 107.200 20.440 ;
        RECT 107.370 20.260 107.680 20.440 ;
        RECT 107.850 20.260 108.160 20.440 ;
        RECT 108.330 20.260 108.640 20.440 ;
        RECT 108.810 20.260 109.120 20.440 ;
        RECT 109.290 20.260 109.600 20.440 ;
        RECT 109.770 20.260 110.080 20.440 ;
        RECT 110.250 20.260 110.560 20.440 ;
        RECT 110.730 20.260 111.040 20.440 ;
        RECT 111.210 20.260 111.520 20.440 ;
        RECT 111.690 20.260 112.000 20.440 ;
        RECT 112.170 20.260 112.480 20.440 ;
        RECT 112.650 20.260 112.960 20.440 ;
        RECT 113.130 20.260 113.440 20.440 ;
        RECT 113.610 20.260 113.920 20.440 ;
        RECT 114.090 20.260 114.400 20.440 ;
        RECT 114.570 20.260 114.880 20.440 ;
        RECT 115.050 20.260 115.360 20.440 ;
        RECT 115.530 20.260 115.840 20.440 ;
        RECT 116.010 20.260 116.320 20.440 ;
        RECT 116.490 20.260 116.800 20.440 ;
        RECT 116.970 20.260 117.280 20.440 ;
        RECT 117.450 20.260 117.760 20.440 ;
        RECT 117.930 20.260 118.240 20.440 ;
        RECT 118.410 20.260 118.720 20.440 ;
        RECT 118.890 20.260 119.200 20.440 ;
        RECT 119.370 20.260 119.680 20.440 ;
        RECT 119.850 20.260 120.160 20.440 ;
        RECT 120.330 20.260 120.640 20.440 ;
        RECT 120.810 20.260 121.120 20.440 ;
        RECT 121.290 20.260 121.600 20.440 ;
        RECT 121.770 20.260 122.080 20.440 ;
        RECT 122.250 20.260 122.560 20.440 ;
        RECT 122.730 20.260 123.040 20.440 ;
        RECT 123.210 20.260 123.520 20.440 ;
        RECT 123.690 20.260 124.000 20.440 ;
        RECT 124.170 20.260 124.480 20.440 ;
        RECT 124.650 20.260 124.960 20.440 ;
        RECT 125.130 20.260 125.440 20.440 ;
        RECT 125.610 20.260 125.920 20.440 ;
        RECT 126.090 20.260 126.400 20.440 ;
        RECT 126.570 20.260 126.880 20.440 ;
        RECT 127.050 20.260 127.360 20.440 ;
        RECT 127.530 20.260 127.840 20.440 ;
        RECT 128.010 20.260 128.320 20.440 ;
        RECT 128.490 20.260 128.800 20.440 ;
        RECT 128.970 20.260 129.280 20.440 ;
        RECT 129.450 20.260 129.760 20.440 ;
        RECT 129.930 20.260 130.240 20.440 ;
        RECT 130.410 20.260 130.720 20.440 ;
        RECT 130.890 20.260 131.200 20.440 ;
        RECT 131.370 20.260 131.680 20.440 ;
        RECT 131.850 20.260 132.160 20.440 ;
        RECT 132.330 20.260 132.640 20.440 ;
        RECT 132.810 20.260 133.120 20.440 ;
        RECT 133.290 20.260 133.600 20.440 ;
        RECT 133.770 20.260 134.080 20.440 ;
        RECT 134.250 20.260 134.560 20.440 ;
        RECT 134.730 20.260 135.040 20.440 ;
        RECT 135.210 20.260 135.520 20.440 ;
        RECT 135.690 20.260 136.000 20.440 ;
        RECT 136.170 20.260 136.480 20.440 ;
        RECT 136.650 20.260 136.960 20.440 ;
        RECT 137.130 20.260 137.440 20.440 ;
        RECT 137.610 20.260 137.920 20.440 ;
        RECT 138.090 20.260 138.400 20.440 ;
        RECT 138.570 20.260 138.880 20.440 ;
        RECT 139.050 20.260 139.360 20.440 ;
        RECT 139.530 20.260 139.840 20.440 ;
        RECT 140.010 20.260 140.320 20.440 ;
        RECT 140.490 20.260 140.800 20.440 ;
        RECT 140.970 20.260 141.280 20.440 ;
        RECT 141.450 20.260 141.760 20.440 ;
        RECT 141.930 20.260 142.080 20.440 ;
        RECT 6.340 19.960 9.070 19.990 ;
        RECT 6.340 19.790 6.510 19.960 ;
        RECT 6.680 19.790 6.950 19.960 ;
        RECT 7.120 19.790 7.360 19.960 ;
        RECT 7.530 19.790 7.790 19.960 ;
        RECT 7.960 19.790 8.230 19.960 ;
        RECT 8.400 19.790 8.640 19.960 ;
        RECT 8.810 19.790 9.070 19.960 ;
        RECT 6.340 18.990 9.070 19.790 ;
        RECT 9.770 19.950 11.380 19.980 ;
        RECT 9.770 19.780 9.820 19.950 ;
        RECT 9.990 19.780 10.260 19.950 ;
        RECT 10.430 19.780 10.700 19.950 ;
        RECT 10.870 19.780 11.110 19.950 ;
        RECT 11.280 19.780 11.380 19.950 ;
        RECT 13.060 19.950 13.710 20.060 ;
        RECT 9.770 19.500 11.380 19.780 ;
        RECT 10.080 19.100 11.380 19.500 ;
      LAYER li1 ;
        RECT 11.810 19.280 12.390 19.920 ;
      LAYER li1 ;
        RECT 13.060 19.780 13.120 19.950 ;
        RECT 13.290 19.780 13.480 19.950 ;
        RECT 13.650 19.780 13.710 19.950 ;
        RECT 13.060 19.720 13.710 19.780 ;
        RECT 13.300 19.280 13.710 19.720 ;
        RECT 14.090 19.950 15.700 19.980 ;
        RECT 14.090 19.780 14.140 19.950 ;
        RECT 14.310 19.780 14.580 19.950 ;
        RECT 14.750 19.780 15.020 19.950 ;
        RECT 15.190 19.780 15.430 19.950 ;
        RECT 15.600 19.780 15.700 19.950 ;
        RECT 17.380 19.950 18.030 20.060 ;
        RECT 14.090 19.500 15.700 19.780 ;
        RECT 6.500 18.320 6.830 18.990 ;
        RECT 7.230 17.670 7.560 18.650 ;
        RECT 7.780 18.320 8.110 18.990 ;
        RECT 8.510 17.670 8.840 18.650 ;
        RECT 10.080 18.320 10.410 19.100 ;
        RECT 6.260 16.790 9.000 17.670 ;
        RECT 10.620 17.660 10.950 18.650 ;
      LAYER li1 ;
        RECT 12.140 18.410 12.390 19.280 ;
      LAYER li1 ;
        RECT 14.400 19.100 15.700 19.500 ;
      LAYER li1 ;
        RECT 16.130 19.280 16.710 19.920 ;
      LAYER li1 ;
        RECT 17.380 19.780 17.440 19.950 ;
        RECT 17.610 19.780 17.800 19.950 ;
        RECT 17.970 19.780 18.030 19.950 ;
        RECT 17.380 19.720 18.030 19.780 ;
        RECT 17.620 19.280 18.030 19.720 ;
        RECT 18.410 19.950 20.020 19.980 ;
        RECT 18.410 19.780 18.460 19.950 ;
        RECT 18.630 19.780 18.900 19.950 ;
        RECT 19.070 19.780 19.340 19.950 ;
        RECT 19.510 19.780 19.750 19.950 ;
        RECT 19.920 19.780 20.020 19.950 ;
        RECT 21.700 19.950 22.350 20.060 ;
        RECT 18.410 19.500 20.020 19.780 ;
      LAYER li1 ;
        RECT 12.140 18.160 12.850 18.410 ;
      LAYER li1 ;
        RECT 14.400 18.320 14.730 19.100 ;
        RECT 6.260 16.620 6.470 16.790 ;
        RECT 6.640 16.620 6.910 16.790 ;
        RECT 7.080 16.620 7.320 16.790 ;
        RECT 7.490 16.620 7.750 16.790 ;
        RECT 7.920 16.620 8.190 16.790 ;
        RECT 8.360 16.620 8.600 16.790 ;
        RECT 8.770 16.620 9.000 16.790 ;
        RECT 6.260 16.600 9.000 16.620 ;
        RECT 9.850 16.790 11.300 17.660 ;
        RECT 9.850 16.620 10.100 16.790 ;
        RECT 10.270 16.620 10.460 16.790 ;
        RECT 10.630 16.620 10.900 16.790 ;
        RECT 11.070 16.620 11.300 16.790 ;
        RECT 9.850 16.590 11.300 16.620 ;
        RECT 11.740 16.900 12.140 17.170 ;
        RECT 11.740 16.840 12.390 16.900 ;
        RECT 11.740 16.670 11.800 16.840 ;
        RECT 11.970 16.670 12.160 16.840 ;
        RECT 12.330 16.670 12.390 16.840 ;
      LAYER li1 ;
        RECT 12.600 16.820 12.850 18.160 ;
      LAYER li1 ;
        RECT 14.940 17.660 15.270 18.650 ;
      LAYER li1 ;
        RECT 16.460 18.410 16.710 19.280 ;
      LAYER li1 ;
        RECT 18.720 19.100 20.020 19.500 ;
      LAYER li1 ;
        RECT 16.460 18.160 17.170 18.410 ;
      LAYER li1 ;
        RECT 18.720 18.320 19.050 19.100 ;
      LAYER li1 ;
        RECT 21.200 18.850 21.530 19.850 ;
      LAYER li1 ;
        RECT 21.700 19.780 21.760 19.950 ;
        RECT 21.930 19.780 22.120 19.950 ;
        RECT 22.290 19.780 22.350 19.950 ;
        RECT 21.700 19.720 22.350 19.780 ;
        RECT 21.940 19.280 22.350 19.720 ;
        RECT 22.730 19.950 24.340 19.980 ;
        RECT 25.030 19.950 26.280 19.980 ;
        RECT 27.050 19.950 28.660 19.980 ;
        RECT 29.350 19.950 30.600 19.980 ;
        RECT 31.370 19.950 32.980 19.980 ;
        RECT 33.670 19.950 34.920 19.980 ;
        RECT 35.690 19.950 37.300 19.980 ;
        RECT 22.730 19.780 22.780 19.950 ;
        RECT 22.950 19.780 23.220 19.950 ;
        RECT 23.390 19.780 23.660 19.950 ;
        RECT 23.830 19.780 24.070 19.950 ;
        RECT 24.240 19.780 24.340 19.950 ;
        RECT 22.730 19.500 24.340 19.780 ;
        RECT 23.040 19.100 24.340 19.500 ;
        RECT 11.740 16.560 12.390 16.670 ;
        RECT 14.170 16.790 15.620 17.660 ;
        RECT 14.170 16.620 14.420 16.790 ;
        RECT 14.590 16.620 14.780 16.790 ;
        RECT 14.950 16.620 15.220 16.790 ;
        RECT 15.390 16.620 15.620 16.790 ;
        RECT 14.170 16.590 15.620 16.620 ;
        RECT 16.060 16.900 16.460 17.170 ;
        RECT 16.060 16.840 16.710 16.900 ;
        RECT 16.060 16.670 16.120 16.840 ;
        RECT 16.290 16.670 16.480 16.840 ;
        RECT 16.650 16.670 16.710 16.840 ;
      LAYER li1 ;
        RECT 16.920 16.820 17.170 18.160 ;
      LAYER li1 ;
        RECT 19.260 17.660 19.590 18.650 ;
      LAYER li1 ;
        RECT 21.200 18.580 21.960 18.850 ;
      LAYER li1 ;
        RECT 16.060 16.560 16.710 16.670 ;
        RECT 18.490 16.790 19.940 17.660 ;
      LAYER li1 ;
        RECT 21.690 17.170 21.960 18.580 ;
      LAYER li1 ;
        RECT 23.040 18.320 23.370 19.100 ;
        RECT 23.580 17.660 23.910 18.650 ;
      LAYER li1 ;
        RECT 24.600 18.170 24.850 19.850 ;
      LAYER li1 ;
        RECT 25.200 19.780 25.390 19.950 ;
        RECT 25.560 19.780 25.750 19.950 ;
        RECT 25.920 19.780 26.110 19.950 ;
        RECT 25.030 19.410 26.280 19.780 ;
        RECT 26.460 19.230 26.710 19.850 ;
        RECT 27.050 19.780 27.100 19.950 ;
        RECT 27.270 19.780 27.540 19.950 ;
        RECT 27.710 19.780 27.980 19.950 ;
        RECT 28.150 19.780 28.390 19.950 ;
        RECT 28.560 19.780 28.660 19.950 ;
        RECT 27.050 19.500 28.660 19.780 ;
        RECT 25.160 19.060 26.710 19.230 ;
        RECT 25.160 18.600 25.490 19.060 ;
        RECT 18.490 16.620 18.740 16.790 ;
        RECT 18.910 16.620 19.100 16.790 ;
        RECT 19.270 16.620 19.540 16.790 ;
        RECT 19.710 16.620 19.940 16.790 ;
        RECT 18.490 16.590 19.940 16.620 ;
        RECT 20.380 16.900 20.780 17.170 ;
        RECT 20.380 16.840 21.030 16.900 ;
        RECT 20.380 16.670 20.440 16.840 ;
        RECT 20.610 16.670 20.800 16.840 ;
        RECT 20.970 16.670 21.030 16.840 ;
        RECT 20.380 16.560 21.030 16.670 ;
      LAYER li1 ;
        RECT 21.690 16.530 22.270 17.170 ;
      LAYER li1 ;
        RECT 22.810 16.790 24.260 17.660 ;
        RECT 22.810 16.620 23.060 16.790 ;
        RECT 23.230 16.620 23.420 16.790 ;
        RECT 23.590 16.620 23.860 16.790 ;
        RECT 24.030 16.620 24.260 16.790 ;
        RECT 22.810 16.590 24.260 16.620 ;
      LAYER li1 ;
        RECT 24.600 16.590 25.030 18.170 ;
      LAYER li1 ;
        RECT 25.210 16.840 25.770 18.170 ;
      LAYER li1 ;
        RECT 25.950 17.090 26.280 18.880 ;
      LAYER li1 ;
        RECT 26.460 17.340 26.710 19.060 ;
        RECT 27.360 19.100 28.660 19.500 ;
        RECT 27.360 18.320 27.690 19.100 ;
        RECT 27.900 17.660 28.230 18.650 ;
      LAYER li1 ;
        RECT 28.920 18.170 29.170 19.850 ;
      LAYER li1 ;
        RECT 29.520 19.780 29.710 19.950 ;
        RECT 29.880 19.780 30.070 19.950 ;
        RECT 30.240 19.780 30.430 19.950 ;
        RECT 29.350 19.410 30.600 19.780 ;
        RECT 30.780 19.230 31.030 19.850 ;
        RECT 31.370 19.780 31.420 19.950 ;
        RECT 31.590 19.780 31.860 19.950 ;
        RECT 32.030 19.780 32.300 19.950 ;
        RECT 32.470 19.780 32.710 19.950 ;
        RECT 32.880 19.780 32.980 19.950 ;
        RECT 31.370 19.500 32.980 19.780 ;
        RECT 29.480 19.060 31.030 19.230 ;
        RECT 29.480 18.600 29.810 19.060 ;
        RECT 25.210 16.670 25.220 16.840 ;
        RECT 25.390 16.670 25.580 16.840 ;
        RECT 25.750 16.670 25.770 16.840 ;
        RECT 25.210 16.590 25.770 16.670 ;
        RECT 27.130 16.790 28.580 17.660 ;
        RECT 27.130 16.620 27.380 16.790 ;
        RECT 27.550 16.620 27.740 16.790 ;
        RECT 27.910 16.620 28.180 16.790 ;
        RECT 28.350 16.620 28.580 16.790 ;
        RECT 27.130 16.590 28.580 16.620 ;
      LAYER li1 ;
        RECT 28.920 16.590 29.350 18.170 ;
      LAYER li1 ;
        RECT 29.530 16.840 30.090 18.170 ;
      LAYER li1 ;
        RECT 30.270 17.090 30.600 18.880 ;
      LAYER li1 ;
        RECT 30.780 17.340 31.030 19.060 ;
        RECT 31.680 19.100 32.980 19.500 ;
        RECT 31.680 18.320 32.010 19.100 ;
        RECT 32.220 17.660 32.550 18.650 ;
      LAYER li1 ;
        RECT 33.240 18.170 33.490 19.850 ;
      LAYER li1 ;
        RECT 33.840 19.780 34.030 19.950 ;
        RECT 34.200 19.780 34.390 19.950 ;
        RECT 34.560 19.780 34.750 19.950 ;
        RECT 33.670 19.410 34.920 19.780 ;
        RECT 35.100 19.230 35.350 19.850 ;
        RECT 35.690 19.780 35.740 19.950 ;
        RECT 35.910 19.780 36.180 19.950 ;
        RECT 36.350 19.780 36.620 19.950 ;
        RECT 36.790 19.780 37.030 19.950 ;
        RECT 37.200 19.780 37.300 19.950 ;
        RECT 35.690 19.500 37.300 19.780 ;
        RECT 33.800 19.060 35.350 19.230 ;
        RECT 33.800 18.600 34.130 19.060 ;
        RECT 29.530 16.670 29.540 16.840 ;
        RECT 29.710 16.670 29.900 16.840 ;
        RECT 30.070 16.670 30.090 16.840 ;
        RECT 29.530 16.590 30.090 16.670 ;
        RECT 31.450 16.790 32.900 17.660 ;
        RECT 31.450 16.620 31.700 16.790 ;
        RECT 31.870 16.620 32.060 16.790 ;
        RECT 32.230 16.620 32.500 16.790 ;
        RECT 32.670 16.620 32.900 16.790 ;
        RECT 31.450 16.590 32.900 16.620 ;
      LAYER li1 ;
        RECT 33.240 16.590 33.670 18.170 ;
      LAYER li1 ;
        RECT 33.850 16.840 34.410 18.170 ;
      LAYER li1 ;
        RECT 34.590 17.090 34.920 18.880 ;
      LAYER li1 ;
        RECT 35.100 17.340 35.350 19.060 ;
        RECT 36.000 19.100 37.300 19.500 ;
        RECT 38.010 19.950 38.600 19.980 ;
        RECT 38.010 19.780 38.040 19.950 ;
        RECT 38.210 19.780 38.400 19.950 ;
        RECT 38.570 19.780 38.600 19.950 ;
        RECT 39.530 19.950 41.140 19.980 ;
        RECT 41.830 19.950 43.080 19.980 ;
        RECT 43.850 19.950 45.460 19.980 ;
        RECT 36.000 18.320 36.330 19.100 ;
        RECT 38.010 19.020 38.600 19.780 ;
        RECT 36.540 17.660 36.870 18.650 ;
      LAYER li1 ;
        RECT 38.050 18.410 38.760 18.800 ;
        RECT 38.940 18.170 39.270 19.850 ;
      LAYER li1 ;
        RECT 39.530 19.780 39.580 19.950 ;
        RECT 39.750 19.780 40.020 19.950 ;
        RECT 40.190 19.780 40.460 19.950 ;
        RECT 40.630 19.780 40.870 19.950 ;
        RECT 41.040 19.780 41.140 19.950 ;
        RECT 39.530 19.500 41.140 19.780 ;
        RECT 39.840 19.100 41.140 19.500 ;
        RECT 39.840 18.320 40.170 19.100 ;
        RECT 33.850 16.670 33.860 16.840 ;
        RECT 34.030 16.670 34.220 16.840 ;
        RECT 34.390 16.670 34.410 16.840 ;
        RECT 33.850 16.590 34.410 16.670 ;
        RECT 35.770 16.790 37.220 17.660 ;
        RECT 35.770 16.620 36.020 16.790 ;
        RECT 36.190 16.620 36.380 16.790 ;
        RECT 36.550 16.620 36.820 16.790 ;
        RECT 36.990 16.620 37.220 16.790 ;
        RECT 35.770 16.590 37.220 16.620 ;
        RECT 38.010 16.840 38.600 18.170 ;
        RECT 38.010 16.670 38.040 16.840 ;
        RECT 38.210 16.670 38.400 16.840 ;
        RECT 38.570 16.670 38.600 16.840 ;
        RECT 38.010 16.590 38.600 16.670 ;
      LAYER li1 ;
        RECT 38.880 16.590 39.270 18.170 ;
      LAYER li1 ;
        RECT 40.380 17.660 40.710 18.650 ;
      LAYER li1 ;
        RECT 41.400 18.170 41.650 19.850 ;
      LAYER li1 ;
        RECT 42.000 19.780 42.190 19.950 ;
        RECT 42.360 19.780 42.550 19.950 ;
        RECT 42.720 19.780 42.910 19.950 ;
        RECT 41.830 19.410 43.080 19.780 ;
        RECT 43.260 19.230 43.510 19.850 ;
        RECT 43.850 19.780 43.900 19.950 ;
        RECT 44.070 19.780 44.340 19.950 ;
        RECT 44.510 19.780 44.780 19.950 ;
        RECT 44.950 19.780 45.190 19.950 ;
        RECT 45.360 19.780 45.460 19.950 ;
        RECT 43.850 19.500 45.460 19.780 ;
        RECT 41.960 19.060 43.510 19.230 ;
        RECT 41.960 18.600 42.290 19.060 ;
        RECT 39.610 16.790 41.060 17.660 ;
        RECT 39.610 16.620 39.860 16.790 ;
        RECT 40.030 16.620 40.220 16.790 ;
        RECT 40.390 16.620 40.660 16.790 ;
        RECT 40.830 16.620 41.060 16.790 ;
        RECT 39.610 16.590 41.060 16.620 ;
      LAYER li1 ;
        RECT 41.400 16.590 41.830 18.170 ;
      LAYER li1 ;
        RECT 42.010 16.840 42.570 18.170 ;
      LAYER li1 ;
        RECT 42.750 17.090 43.080 18.880 ;
      LAYER li1 ;
        RECT 43.260 17.340 43.510 19.060 ;
        RECT 44.160 19.100 45.460 19.500 ;
        RECT 45.690 19.950 46.280 19.980 ;
        RECT 45.690 19.780 45.720 19.950 ;
        RECT 45.890 19.780 46.080 19.950 ;
        RECT 46.250 19.780 46.280 19.950 ;
        RECT 46.960 19.950 47.910 19.980 ;
        RECT 44.160 18.320 44.490 19.100 ;
        RECT 45.690 19.020 46.280 19.780 ;
      LAYER li1 ;
        RECT 46.530 18.920 46.780 19.850 ;
      LAYER li1 ;
        RECT 46.960 19.780 46.990 19.950 ;
        RECT 47.160 19.780 47.350 19.950 ;
        RECT 47.520 19.780 47.710 19.950 ;
        RECT 47.880 19.780 47.910 19.950 ;
        RECT 49.130 19.950 50.740 19.980 ;
        RECT 46.960 19.100 47.910 19.780 ;
      LAYER li1 ;
        RECT 48.090 18.920 48.360 19.850 ;
      LAYER li1 ;
        RECT 49.130 19.780 49.180 19.950 ;
        RECT 49.350 19.780 49.620 19.950 ;
        RECT 49.790 19.780 50.060 19.950 ;
        RECT 50.230 19.780 50.470 19.950 ;
        RECT 50.640 19.780 50.740 19.950 ;
        RECT 49.130 19.500 50.740 19.780 ;
        RECT 44.700 17.660 45.030 18.650 ;
      LAYER li1 ;
        RECT 45.730 18.230 46.030 18.820 ;
        RECT 46.530 18.750 48.360 18.920 ;
        RECT 46.210 18.230 47.400 18.570 ;
      LAYER li1 ;
        RECT 42.010 16.670 42.020 16.840 ;
        RECT 42.190 16.670 42.380 16.840 ;
        RECT 42.550 16.670 42.570 16.840 ;
        RECT 42.010 16.590 42.570 16.670 ;
        RECT 43.930 16.790 45.380 17.660 ;
        RECT 43.930 16.620 44.180 16.790 ;
        RECT 44.350 16.620 44.540 16.790 ;
        RECT 44.710 16.620 44.980 16.790 ;
        RECT 45.150 16.620 45.380 16.790 ;
        RECT 43.930 16.590 45.380 16.620 ;
        RECT 45.690 16.840 47.360 18.050 ;
      LAYER li1 ;
        RECT 47.580 17.090 47.910 18.570 ;
      LAYER li1 ;
        RECT 45.690 16.670 45.720 16.840 ;
        RECT 45.890 16.670 46.080 16.840 ;
        RECT 46.250 16.670 46.440 16.840 ;
        RECT 46.610 16.670 46.800 16.840 ;
        RECT 46.970 16.670 47.160 16.840 ;
        RECT 47.330 16.670 47.360 16.840 ;
        RECT 45.690 16.590 47.360 16.670 ;
      LAYER li1 ;
        RECT 48.090 16.590 48.360 18.750 ;
      LAYER li1 ;
        RECT 49.440 19.100 50.740 19.500 ;
        RECT 50.970 19.950 51.560 19.980 ;
        RECT 50.970 19.780 51.000 19.950 ;
        RECT 51.170 19.780 51.360 19.950 ;
        RECT 51.530 19.780 51.560 19.950 ;
        RECT 52.240 19.950 53.190 19.980 ;
      LAYER li1 ;
        RECT 48.630 17.120 48.800 18.400 ;
      LAYER li1 ;
        RECT 49.440 18.320 49.770 19.100 ;
        RECT 50.970 19.020 51.560 19.780 ;
      LAYER li1 ;
        RECT 51.810 18.920 52.060 19.850 ;
      LAYER li1 ;
        RECT 52.240 19.780 52.270 19.950 ;
        RECT 52.440 19.780 52.630 19.950 ;
        RECT 52.800 19.780 52.990 19.950 ;
        RECT 53.160 19.780 53.190 19.950 ;
        RECT 54.410 19.950 56.020 19.980 ;
        RECT 52.240 19.100 53.190 19.780 ;
      LAYER li1 ;
        RECT 53.370 18.920 53.640 19.850 ;
      LAYER li1 ;
        RECT 54.410 19.780 54.460 19.950 ;
        RECT 54.630 19.780 54.900 19.950 ;
        RECT 55.070 19.780 55.340 19.950 ;
        RECT 55.510 19.780 55.750 19.950 ;
        RECT 55.920 19.780 56.020 19.950 ;
        RECT 54.410 19.500 56.020 19.780 ;
        RECT 49.980 17.660 50.310 18.650 ;
      LAYER li1 ;
        RECT 51.010 18.230 51.310 18.820 ;
        RECT 51.810 18.750 53.640 18.920 ;
        RECT 51.490 18.230 52.680 18.570 ;
      LAYER li1 ;
        RECT 49.210 16.790 50.660 17.660 ;
        RECT 49.210 16.620 49.460 16.790 ;
        RECT 49.630 16.620 49.820 16.790 ;
        RECT 49.990 16.620 50.260 16.790 ;
        RECT 50.430 16.620 50.660 16.790 ;
        RECT 49.210 16.590 50.660 16.620 ;
        RECT 50.970 16.840 52.640 18.050 ;
      LAYER li1 ;
        RECT 52.860 17.090 53.190 18.570 ;
      LAYER li1 ;
        RECT 50.970 16.670 51.000 16.840 ;
        RECT 51.170 16.670 51.360 16.840 ;
        RECT 51.530 16.670 51.720 16.840 ;
        RECT 51.890 16.670 52.080 16.840 ;
        RECT 52.250 16.670 52.440 16.840 ;
        RECT 52.610 16.670 52.640 16.840 ;
        RECT 50.970 16.590 52.640 16.670 ;
      LAYER li1 ;
        RECT 53.370 16.590 53.640 18.750 ;
      LAYER li1 ;
        RECT 54.720 19.100 56.020 19.500 ;
        RECT 56.250 19.950 56.840 19.980 ;
        RECT 56.250 19.780 56.280 19.950 ;
        RECT 56.450 19.780 56.640 19.950 ;
        RECT 56.810 19.780 56.840 19.950 ;
        RECT 57.770 19.950 59.380 19.980 ;
        RECT 54.720 18.320 55.050 19.100 ;
        RECT 56.250 19.020 56.840 19.780 ;
        RECT 55.260 17.660 55.590 18.650 ;
      LAYER li1 ;
        RECT 56.290 18.410 57.000 18.800 ;
        RECT 57.180 18.170 57.510 19.850 ;
      LAYER li1 ;
        RECT 57.770 19.780 57.820 19.950 ;
        RECT 57.990 19.780 58.260 19.950 ;
        RECT 58.430 19.780 58.700 19.950 ;
        RECT 58.870 19.780 59.110 19.950 ;
        RECT 59.280 19.780 59.380 19.950 ;
        RECT 57.770 19.500 59.380 19.780 ;
        RECT 58.080 19.100 59.380 19.500 ;
        RECT 59.610 19.950 60.560 19.980 ;
        RECT 59.610 19.780 59.640 19.950 ;
        RECT 59.810 19.780 60.000 19.950 ;
        RECT 60.170 19.780 60.360 19.950 ;
        RECT 60.530 19.780 60.560 19.950 ;
        RECT 61.170 19.950 62.120 19.980 ;
        RECT 58.080 18.320 58.410 19.100 ;
        RECT 59.610 19.020 60.560 19.780 ;
      LAYER li1 ;
        RECT 60.740 19.140 60.990 19.850 ;
      LAYER li1 ;
        RECT 61.170 19.780 61.200 19.950 ;
        RECT 61.370 19.780 61.560 19.950 ;
        RECT 61.730 19.780 61.920 19.950 ;
        RECT 62.090 19.780 62.120 19.950 ;
        RECT 62.730 19.950 63.680 19.980 ;
        RECT 61.170 19.320 62.120 19.780 ;
      LAYER li1 ;
        RECT 62.300 19.140 62.550 19.850 ;
        RECT 60.740 18.970 62.550 19.140 ;
      LAYER li1 ;
        RECT 62.730 19.780 62.760 19.950 ;
        RECT 62.930 19.780 63.120 19.950 ;
        RECT 63.290 19.780 63.480 19.950 ;
        RECT 63.650 19.780 63.680 19.950 ;
        RECT 64.490 19.950 66.100 19.980 ;
        RECT 62.730 19.100 63.680 19.780 ;
      LAYER li1 ;
        RECT 60.740 18.800 60.910 18.970 ;
      LAYER li1 ;
        RECT 63.860 18.920 64.190 19.850 ;
        RECT 64.490 19.780 64.540 19.950 ;
        RECT 64.710 19.780 64.980 19.950 ;
        RECT 65.150 19.780 65.420 19.950 ;
        RECT 65.590 19.780 65.830 19.950 ;
        RECT 66.000 19.780 66.100 19.950 ;
        RECT 64.490 19.500 66.100 19.780 ;
        RECT 54.490 16.790 55.940 17.660 ;
        RECT 54.490 16.620 54.740 16.790 ;
        RECT 54.910 16.620 55.100 16.790 ;
        RECT 55.270 16.620 55.540 16.790 ;
        RECT 55.710 16.620 55.940 16.790 ;
        RECT 54.490 16.590 55.940 16.620 ;
        RECT 56.250 16.840 56.840 18.170 ;
        RECT 56.250 16.670 56.280 16.840 ;
        RECT 56.450 16.670 56.640 16.840 ;
        RECT 56.810 16.670 56.840 16.840 ;
        RECT 56.250 16.590 56.840 16.670 ;
      LAYER li1 ;
        RECT 57.120 16.590 57.510 18.170 ;
      LAYER li1 ;
        RECT 58.620 17.660 58.950 18.650 ;
      LAYER li1 ;
        RECT 59.650 18.570 60.910 18.800 ;
      LAYER li1 ;
        RECT 62.950 18.790 64.190 18.920 ;
        RECT 61.090 18.750 64.190 18.790 ;
        RECT 61.090 18.620 63.120 18.750 ;
      LAYER li1 ;
        RECT 60.740 18.440 60.910 18.570 ;
        RECT 60.740 18.270 62.630 18.440 ;
      LAYER li1 ;
        RECT 57.850 16.790 59.300 17.660 ;
        RECT 57.850 16.620 58.100 16.790 ;
        RECT 58.270 16.620 58.460 16.790 ;
        RECT 58.630 16.620 58.900 16.790 ;
        RECT 59.070 16.620 59.300 16.790 ;
        RECT 57.850 16.590 59.300 16.620 ;
        RECT 59.610 16.840 60.560 18.170 ;
        RECT 59.610 16.670 59.640 16.840 ;
        RECT 59.810 16.670 60.000 16.840 ;
        RECT 60.170 16.670 60.360 16.840 ;
        RECT 60.530 16.670 60.560 16.840 ;
        RECT 59.610 16.590 60.560 16.670 ;
      LAYER li1 ;
        RECT 60.740 16.590 60.990 18.270 ;
      LAYER li1 ;
        RECT 61.170 16.840 62.120 18.090 ;
        RECT 61.170 16.670 61.200 16.840 ;
        RECT 61.370 16.670 61.560 16.840 ;
        RECT 61.730 16.670 61.920 16.840 ;
        RECT 62.090 16.670 62.120 16.840 ;
        RECT 61.170 16.590 62.120 16.670 ;
      LAYER li1 ;
        RECT 62.300 16.590 62.630 18.270 ;
        RECT 63.410 18.230 63.740 18.570 ;
      LAYER li1 ;
        RECT 62.810 16.840 63.760 18.050 ;
        RECT 62.810 16.670 62.840 16.840 ;
        RECT 63.010 16.670 63.200 16.840 ;
        RECT 63.370 16.670 63.560 16.840 ;
        RECT 63.730 16.670 63.760 16.840 ;
        RECT 62.810 16.590 63.760 16.670 ;
        RECT 63.940 16.590 64.190 18.750 ;
        RECT 64.800 19.100 66.100 19.500 ;
        RECT 66.400 19.910 68.210 20.080 ;
        RECT 64.800 18.320 65.130 19.100 ;
        RECT 66.400 18.990 66.730 19.910 ;
      LAYER li1 ;
        RECT 66.980 19.510 67.510 19.730 ;
        RECT 66.980 19.340 67.520 19.510 ;
        RECT 66.980 18.990 67.510 19.340 ;
      LAYER li1 ;
        RECT 65.340 17.660 65.670 18.650 ;
      LAYER li1 ;
        RECT 66.370 18.480 66.790 18.810 ;
        RECT 66.980 18.420 67.150 18.990 ;
      LAYER li1 ;
        RECT 68.040 18.890 68.210 19.910 ;
        RECT 68.390 19.950 69.490 19.980 ;
        RECT 68.390 19.780 68.440 19.950 ;
        RECT 68.610 19.780 68.800 19.950 ;
        RECT 68.970 19.780 69.160 19.950 ;
        RECT 69.330 19.780 69.490 19.950 ;
        RECT 70.250 19.950 71.860 19.980 ;
        RECT 72.550 19.950 73.800 19.980 ;
        RECT 74.570 19.950 76.180 19.980 ;
        RECT 76.870 19.950 78.120 19.980 ;
        RECT 79.300 19.960 82.030 19.990 ;
        RECT 68.390 19.070 69.490 19.780 ;
        RECT 69.660 18.890 69.910 19.820 ;
        RECT 70.250 19.780 70.300 19.950 ;
        RECT 70.470 19.780 70.740 19.950 ;
        RECT 70.910 19.780 71.180 19.950 ;
        RECT 71.350 19.780 71.590 19.950 ;
        RECT 71.760 19.780 71.860 19.950 ;
        RECT 70.250 19.500 71.860 19.780 ;
      LAYER li1 ;
        RECT 67.330 18.600 67.840 18.810 ;
      LAYER li1 ;
        RECT 68.040 18.720 69.910 18.890 ;
        RECT 70.560 19.100 71.860 19.500 ;
      LAYER li1 ;
        RECT 66.980 18.250 68.040 18.420 ;
        RECT 67.770 18.170 68.040 18.250 ;
        RECT 68.490 18.230 69.000 18.540 ;
        RECT 69.250 18.230 69.960 18.540 ;
      LAYER li1 ;
        RECT 70.560 18.320 70.890 19.100 ;
        RECT 64.570 16.790 66.020 17.660 ;
        RECT 64.570 16.620 64.820 16.790 ;
        RECT 64.990 16.620 65.180 16.790 ;
        RECT 65.350 16.620 65.620 16.790 ;
        RECT 65.790 16.620 66.020 16.790 ;
        RECT 64.570 16.590 66.020 16.620 ;
        RECT 66.330 16.840 67.590 18.070 ;
      LAYER li1 ;
        RECT 67.770 17.090 68.290 18.170 ;
      LAYER li1 ;
        RECT 66.330 16.670 66.340 16.840 ;
        RECT 66.510 16.670 66.700 16.840 ;
        RECT 66.870 16.670 67.060 16.840 ;
        RECT 67.230 16.670 67.420 16.840 ;
        RECT 66.330 16.590 67.590 16.670 ;
      LAYER li1 ;
        RECT 68.120 16.590 68.290 17.090 ;
      LAYER li1 ;
        RECT 68.550 16.840 69.860 18.050 ;
        RECT 71.100 17.660 71.430 18.650 ;
      LAYER li1 ;
        RECT 72.120 18.170 72.370 19.850 ;
      LAYER li1 ;
        RECT 72.720 19.780 72.910 19.950 ;
        RECT 73.080 19.780 73.270 19.950 ;
        RECT 73.440 19.780 73.630 19.950 ;
        RECT 72.550 19.410 73.800 19.780 ;
        RECT 73.980 19.230 74.230 19.850 ;
        RECT 74.570 19.780 74.620 19.950 ;
        RECT 74.790 19.780 75.060 19.950 ;
        RECT 75.230 19.780 75.500 19.950 ;
        RECT 75.670 19.780 75.910 19.950 ;
        RECT 76.080 19.780 76.180 19.950 ;
        RECT 74.570 19.500 76.180 19.780 ;
        RECT 72.680 19.060 74.230 19.230 ;
        RECT 72.680 18.600 73.010 19.060 ;
        RECT 68.550 16.670 68.580 16.840 ;
        RECT 68.750 16.670 68.940 16.840 ;
        RECT 69.110 16.670 69.300 16.840 ;
        RECT 69.470 16.670 69.660 16.840 ;
        RECT 69.830 16.670 69.860 16.840 ;
        RECT 68.550 16.590 69.860 16.670 ;
        RECT 70.330 16.790 71.780 17.660 ;
        RECT 70.330 16.620 70.580 16.790 ;
        RECT 70.750 16.620 70.940 16.790 ;
        RECT 71.110 16.620 71.380 16.790 ;
        RECT 71.550 16.620 71.780 16.790 ;
        RECT 70.330 16.590 71.780 16.620 ;
      LAYER li1 ;
        RECT 72.120 16.590 72.550 18.170 ;
      LAYER li1 ;
        RECT 72.730 16.840 73.290 18.170 ;
        RECT 73.980 17.340 74.230 19.060 ;
        RECT 74.880 19.100 76.180 19.500 ;
        RECT 74.880 18.320 75.210 19.100 ;
        RECT 75.420 17.660 75.750 18.650 ;
      LAYER li1 ;
        RECT 76.440 18.170 76.690 19.850 ;
      LAYER li1 ;
        RECT 77.040 19.780 77.230 19.950 ;
        RECT 77.400 19.780 77.590 19.950 ;
        RECT 77.760 19.780 77.950 19.950 ;
        RECT 76.870 19.410 78.120 19.780 ;
        RECT 78.300 19.230 78.550 19.850 ;
        RECT 77.000 19.060 78.550 19.230 ;
        RECT 77.000 18.600 77.330 19.060 ;
        RECT 72.730 16.670 72.740 16.840 ;
        RECT 72.910 16.670 73.100 16.840 ;
        RECT 73.270 16.670 73.290 16.840 ;
        RECT 72.730 16.590 73.290 16.670 ;
        RECT 74.650 16.790 76.100 17.660 ;
        RECT 74.650 16.620 74.900 16.790 ;
        RECT 75.070 16.620 75.260 16.790 ;
        RECT 75.430 16.620 75.700 16.790 ;
        RECT 75.870 16.620 76.100 16.790 ;
        RECT 74.650 16.590 76.100 16.620 ;
      LAYER li1 ;
        RECT 76.440 16.590 76.870 18.170 ;
      LAYER li1 ;
        RECT 77.050 16.840 77.610 18.170 ;
      LAYER li1 ;
        RECT 77.790 17.090 78.120 18.880 ;
      LAYER li1 ;
        RECT 78.300 17.340 78.550 19.060 ;
        RECT 79.300 19.790 79.470 19.960 ;
        RECT 79.640 19.790 79.910 19.960 ;
        RECT 80.080 19.790 80.320 19.960 ;
        RECT 80.490 19.790 80.750 19.960 ;
        RECT 80.920 19.790 81.190 19.960 ;
        RECT 81.360 19.790 81.600 19.960 ;
        RECT 81.770 19.790 82.030 19.960 ;
        RECT 83.120 19.950 84.070 19.980 ;
        RECT 79.300 18.990 82.030 19.790 ;
        RECT 79.460 18.320 79.790 18.990 ;
        RECT 80.190 17.670 80.520 18.650 ;
        RECT 80.740 18.320 81.070 18.990 ;
        RECT 81.470 17.670 81.800 18.650 ;
        RECT 82.670 17.990 82.940 19.850 ;
        RECT 83.120 19.780 83.150 19.950 ;
        RECT 83.320 19.780 83.510 19.950 ;
        RECT 83.680 19.780 83.870 19.950 ;
        RECT 84.040 19.780 84.070 19.950 ;
        RECT 84.760 19.950 85.350 19.980 ;
        RECT 83.120 19.350 84.070 19.780 ;
        RECT 84.250 19.350 84.580 19.850 ;
        RECT 83.800 17.990 84.130 18.490 ;
        RECT 82.670 17.820 84.130 17.990 ;
        RECT 77.050 16.670 77.060 16.840 ;
        RECT 77.230 16.670 77.420 16.840 ;
        RECT 77.590 16.670 77.610 16.840 ;
        RECT 77.050 16.590 77.610 16.670 ;
        RECT 79.220 16.790 81.960 17.670 ;
        RECT 82.670 16.890 83.000 17.820 ;
        RECT 79.220 16.620 79.430 16.790 ;
        RECT 79.600 16.620 79.870 16.790 ;
        RECT 80.040 16.620 80.280 16.790 ;
        RECT 80.450 16.620 80.710 16.790 ;
        RECT 80.880 16.620 81.150 16.790 ;
        RECT 81.320 16.620 81.560 16.790 ;
        RECT 81.730 16.620 81.960 16.790 ;
        RECT 83.190 16.840 83.780 17.620 ;
        RECT 83.190 16.670 83.220 16.840 ;
        RECT 83.390 16.670 83.580 16.840 ;
        RECT 83.750 16.670 83.780 16.840 ;
        RECT 83.190 16.640 83.780 16.670 ;
        RECT 83.960 16.710 84.130 17.820 ;
        RECT 84.310 18.430 84.580 19.350 ;
        RECT 84.760 19.780 84.790 19.950 ;
        RECT 84.960 19.780 85.150 19.950 ;
        RECT 85.320 19.780 85.350 19.950 ;
        RECT 89.720 19.950 90.670 19.980 ;
        RECT 84.760 19.100 85.350 19.780 ;
      LAYER li1 ;
        RECT 85.630 19.720 88.570 19.890 ;
        RECT 85.630 18.730 85.800 19.720 ;
      LAYER li1 ;
        RECT 84.310 18.200 84.840 18.430 ;
        RECT 84.310 16.890 84.560 18.200 ;
      LAYER li1 ;
        RECT 85.260 17.860 85.800 18.730 ;
        RECT 85.980 18.240 86.310 19.540 ;
      LAYER li1 ;
        RECT 86.490 19.020 86.760 19.520 ;
        RECT 87.210 19.270 87.540 19.520 ;
        RECT 87.210 19.100 88.220 19.270 ;
        RECT 86.490 18.030 86.660 19.020 ;
        RECT 87.540 18.430 87.870 18.920 ;
        RECT 86.440 17.860 86.660 18.030 ;
        RECT 86.840 18.200 87.870 18.430 ;
        RECT 88.050 18.870 88.220 19.100 ;
      LAYER li1 ;
        RECT 88.400 19.220 88.570 19.720 ;
      LAYER li1 ;
        RECT 89.720 19.780 89.750 19.950 ;
        RECT 89.920 19.780 90.110 19.950 ;
        RECT 90.280 19.780 90.470 19.950 ;
        RECT 90.640 19.780 90.670 19.950 ;
        RECT 89.720 19.400 90.670 19.780 ;
      LAYER li1 ;
        RECT 90.850 19.910 93.510 20.080 ;
        RECT 90.850 19.220 91.020 19.910 ;
        RECT 88.400 19.050 91.020 19.220 ;
      LAYER li1 ;
        RECT 88.050 18.700 90.670 18.870 ;
        RECT 86.440 17.680 86.610 17.860 ;
        RECT 86.840 17.680 87.010 18.200 ;
        RECT 88.050 18.020 88.220 18.700 ;
      LAYER li1 ;
        RECT 90.850 18.520 91.020 19.050 ;
      LAYER li1 ;
        RECT 84.800 17.510 86.610 17.680 ;
        RECT 84.800 16.890 85.050 17.510 ;
        RECT 85.230 17.160 86.260 17.330 ;
        RECT 85.230 16.710 85.400 17.160 ;
        RECT 79.220 16.600 81.960 16.620 ;
        RECT 83.960 16.540 85.400 16.710 ;
        RECT 85.580 16.840 85.910 16.980 ;
        RECT 85.580 16.670 85.610 16.840 ;
        RECT 85.780 16.670 85.910 16.840 ;
        RECT 85.580 16.640 85.910 16.670 ;
        RECT 86.090 16.710 86.260 17.160 ;
        RECT 86.440 16.890 86.610 17.510 ;
        RECT 86.790 17.350 87.010 17.680 ;
        RECT 87.190 17.850 88.220 18.020 ;
        RECT 88.400 18.170 88.730 18.520 ;
      LAYER li1 ;
        RECT 89.170 18.350 91.020 18.520 ;
      LAYER li1 ;
        RECT 91.200 19.020 91.530 19.730 ;
        RECT 91.990 19.560 93.160 19.730 ;
        RECT 91.990 19.020 92.320 19.560 ;
        RECT 91.200 18.170 91.460 19.020 ;
        RECT 92.530 18.760 92.810 19.260 ;
        RECT 88.400 18.000 91.460 18.170 ;
        RECT 87.190 17.150 87.360 17.850 ;
        RECT 88.050 17.820 88.220 17.850 ;
        RECT 87.540 17.470 87.870 17.670 ;
        RECT 88.050 17.650 89.820 17.820 ;
        RECT 87.540 17.350 89.310 17.470 ;
        RECT 87.660 17.300 89.310 17.350 ;
        RECT 87.140 16.890 87.470 17.150 ;
        RECT 87.660 16.710 87.830 17.300 ;
        RECT 86.090 16.540 87.830 16.710 ;
        RECT 88.010 16.840 88.960 17.120 ;
        RECT 88.010 16.670 88.040 16.840 ;
        RECT 88.210 16.670 88.400 16.840 ;
        RECT 88.570 16.670 88.760 16.840 ;
        RECT 88.930 16.670 88.960 16.840 ;
        RECT 88.010 16.640 88.960 16.670 ;
        RECT 89.140 16.710 89.310 17.300 ;
        RECT 89.490 16.890 89.820 17.650 ;
        RECT 91.130 17.420 91.460 18.000 ;
        RECT 91.640 18.590 92.810 18.760 ;
        RECT 91.640 17.240 91.810 18.590 ;
        RECT 92.190 17.910 92.520 18.410 ;
        RECT 92.990 18.160 93.160 19.560 ;
      LAYER li1 ;
        RECT 93.340 19.250 93.510 19.910 ;
      LAYER li1 ;
        RECT 93.690 19.950 94.640 19.980 ;
        RECT 93.690 19.780 93.720 19.950 ;
        RECT 93.890 19.780 94.080 19.950 ;
        RECT 94.250 19.780 94.440 19.950 ;
        RECT 94.610 19.780 94.640 19.950 ;
        RECT 96.300 19.950 97.250 19.980 ;
        RECT 93.690 19.430 94.640 19.780 ;
        RECT 95.180 19.350 95.510 19.850 ;
        RECT 96.300 19.780 96.330 19.950 ;
        RECT 96.500 19.780 96.690 19.950 ;
        RECT 96.860 19.780 97.050 19.950 ;
        RECT 97.220 19.780 97.250 19.950 ;
      LAYER li1 ;
        RECT 93.340 19.140 94.350 19.250 ;
        RECT 93.340 19.080 94.400 19.140 ;
        RECT 94.020 18.970 94.400 19.080 ;
      LAYER li1 ;
        RECT 93.370 18.510 93.700 18.900 ;
      LAYER li1 ;
        RECT 94.020 18.690 94.350 18.970 ;
      LAYER li1 ;
        RECT 95.180 18.510 95.410 19.350 ;
        RECT 95.790 18.850 96.120 19.350 ;
        RECT 96.300 18.850 97.250 19.780 ;
        RECT 98.500 19.960 101.230 19.990 ;
        RECT 98.500 19.790 98.670 19.960 ;
        RECT 98.840 19.790 99.110 19.960 ;
        RECT 99.280 19.790 99.520 19.960 ;
        RECT 99.690 19.790 99.950 19.960 ;
        RECT 100.120 19.790 100.390 19.960 ;
        RECT 100.560 19.790 100.800 19.960 ;
        RECT 100.970 19.790 101.230 19.960 ;
        RECT 103.280 19.950 104.230 19.980 ;
        RECT 93.370 18.340 95.410 18.510 ;
        RECT 92.700 17.990 95.060 18.160 ;
        RECT 92.700 17.670 92.870 17.990 ;
        RECT 95.240 17.810 95.410 18.340 ;
        RECT 90.000 17.070 91.810 17.240 ;
        RECT 91.990 17.500 92.870 17.670 ;
        RECT 90.000 16.710 90.170 17.070 ;
        RECT 89.140 16.540 90.170 16.710 ;
        RECT 90.350 16.840 91.300 16.890 ;
        RECT 90.350 16.670 90.380 16.840 ;
        RECT 90.550 16.670 90.740 16.840 ;
        RECT 90.910 16.670 91.100 16.840 ;
        RECT 91.270 16.670 91.300 16.840 ;
        RECT 90.350 16.590 91.300 16.670 ;
        RECT 91.990 16.590 92.240 17.500 ;
        RECT 93.050 16.840 94.000 17.670 ;
        RECT 94.400 17.640 95.410 17.810 ;
        RECT 95.910 18.670 96.120 18.850 ;
        RECT 95.910 18.340 97.280 18.670 ;
        RECT 94.400 17.170 94.650 17.640 ;
        RECT 94.830 16.840 95.730 17.460 ;
        RECT 95.910 17.340 96.160 18.340 ;
        RECT 93.050 16.670 93.080 16.840 ;
        RECT 93.250 16.670 93.440 16.840 ;
        RECT 93.610 16.670 93.800 16.840 ;
        RECT 93.970 16.670 94.000 16.840 ;
        RECT 95.000 16.670 95.190 16.840 ;
        RECT 95.360 16.670 95.550 16.840 ;
        RECT 95.720 16.670 95.730 16.840 ;
        RECT 93.050 16.640 94.000 16.670 ;
        RECT 94.830 16.640 95.730 16.670 ;
        RECT 96.340 16.840 97.280 18.150 ;
        RECT 96.340 16.670 96.360 16.840 ;
        RECT 96.530 16.670 96.720 16.840 ;
        RECT 96.890 16.670 97.080 16.840 ;
        RECT 97.250 16.670 97.280 16.840 ;
        RECT 96.340 16.610 97.280 16.670 ;
      LAYER li1 ;
        RECT 97.460 16.610 97.800 19.680 ;
      LAYER li1 ;
        RECT 98.500 18.990 101.230 19.790 ;
        RECT 98.660 18.320 98.990 18.990 ;
        RECT 99.390 17.670 99.720 18.650 ;
        RECT 99.940 18.320 100.270 18.990 ;
        RECT 100.670 17.670 101.000 18.650 ;
        RECT 102.830 17.990 103.100 19.850 ;
        RECT 103.280 19.780 103.310 19.950 ;
        RECT 103.480 19.780 103.670 19.950 ;
        RECT 103.840 19.780 104.030 19.950 ;
        RECT 104.200 19.780 104.230 19.950 ;
        RECT 104.920 19.950 105.510 19.980 ;
        RECT 103.280 19.350 104.230 19.780 ;
        RECT 104.410 19.350 104.740 19.850 ;
        RECT 103.960 17.990 104.290 18.490 ;
        RECT 102.830 17.820 104.290 17.990 ;
        RECT 98.420 16.790 101.160 17.670 ;
        RECT 102.830 16.890 103.160 17.820 ;
        RECT 98.420 16.620 98.630 16.790 ;
        RECT 98.800 16.620 99.070 16.790 ;
        RECT 99.240 16.620 99.480 16.790 ;
        RECT 99.650 16.620 99.910 16.790 ;
        RECT 100.080 16.620 100.350 16.790 ;
        RECT 100.520 16.620 100.760 16.790 ;
        RECT 100.930 16.620 101.160 16.790 ;
        RECT 103.350 16.840 103.940 17.620 ;
        RECT 103.350 16.670 103.380 16.840 ;
        RECT 103.550 16.670 103.740 16.840 ;
        RECT 103.910 16.670 103.940 16.840 ;
        RECT 103.350 16.640 103.940 16.670 ;
        RECT 104.120 16.710 104.290 17.820 ;
        RECT 104.470 18.430 104.740 19.350 ;
        RECT 104.920 19.780 104.950 19.950 ;
        RECT 105.120 19.780 105.310 19.950 ;
        RECT 105.480 19.780 105.510 19.950 ;
        RECT 109.880 19.950 110.830 19.980 ;
        RECT 104.920 19.100 105.510 19.780 ;
      LAYER li1 ;
        RECT 105.790 19.720 108.730 19.890 ;
        RECT 105.790 18.730 105.960 19.720 ;
      LAYER li1 ;
        RECT 104.470 18.200 105.000 18.430 ;
        RECT 104.470 16.890 104.720 18.200 ;
      LAYER li1 ;
        RECT 105.420 17.860 105.960 18.730 ;
        RECT 106.140 18.240 106.470 19.540 ;
      LAYER li1 ;
        RECT 106.650 19.020 106.920 19.520 ;
        RECT 107.370 19.270 107.700 19.520 ;
        RECT 107.370 19.100 108.380 19.270 ;
        RECT 106.650 18.030 106.820 19.020 ;
        RECT 107.700 18.430 108.030 18.920 ;
        RECT 106.600 17.860 106.820 18.030 ;
        RECT 107.000 18.200 108.030 18.430 ;
        RECT 108.210 18.870 108.380 19.100 ;
      LAYER li1 ;
        RECT 108.560 19.220 108.730 19.720 ;
      LAYER li1 ;
        RECT 109.880 19.780 109.910 19.950 ;
        RECT 110.080 19.780 110.270 19.950 ;
        RECT 110.440 19.780 110.630 19.950 ;
        RECT 110.800 19.780 110.830 19.950 ;
        RECT 109.880 19.400 110.830 19.780 ;
      LAYER li1 ;
        RECT 111.010 19.910 113.670 20.080 ;
        RECT 111.010 19.220 111.180 19.910 ;
        RECT 108.560 19.050 111.180 19.220 ;
      LAYER li1 ;
        RECT 108.210 18.700 110.830 18.870 ;
        RECT 106.600 17.680 106.770 17.860 ;
        RECT 107.000 17.680 107.170 18.200 ;
        RECT 108.210 18.020 108.380 18.700 ;
      LAYER li1 ;
        RECT 111.010 18.520 111.180 19.050 ;
      LAYER li1 ;
        RECT 104.960 17.510 106.770 17.680 ;
        RECT 104.960 16.890 105.210 17.510 ;
        RECT 105.390 17.160 106.420 17.330 ;
        RECT 105.390 16.710 105.560 17.160 ;
        RECT 98.420 16.600 101.160 16.620 ;
        RECT 104.120 16.540 105.560 16.710 ;
        RECT 105.740 16.840 106.070 16.980 ;
        RECT 105.740 16.670 105.770 16.840 ;
        RECT 105.940 16.670 106.070 16.840 ;
        RECT 105.740 16.640 106.070 16.670 ;
        RECT 106.250 16.710 106.420 17.160 ;
        RECT 106.600 16.890 106.770 17.510 ;
        RECT 106.950 17.350 107.170 17.680 ;
        RECT 107.350 17.850 108.380 18.020 ;
        RECT 108.560 18.170 108.890 18.520 ;
      LAYER li1 ;
        RECT 109.330 18.350 111.180 18.520 ;
      LAYER li1 ;
        RECT 111.360 19.020 111.690 19.730 ;
        RECT 112.150 19.560 113.320 19.730 ;
        RECT 112.150 19.020 112.480 19.560 ;
        RECT 111.360 18.170 111.620 19.020 ;
        RECT 112.690 18.760 112.970 19.260 ;
        RECT 108.560 18.000 111.620 18.170 ;
        RECT 107.350 17.150 107.520 17.850 ;
        RECT 108.210 17.820 108.380 17.850 ;
        RECT 107.700 17.470 108.030 17.670 ;
        RECT 108.210 17.650 109.980 17.820 ;
        RECT 107.700 17.350 109.470 17.470 ;
        RECT 107.820 17.300 109.470 17.350 ;
        RECT 107.300 16.890 107.630 17.150 ;
        RECT 107.820 16.710 107.990 17.300 ;
        RECT 106.250 16.540 107.990 16.710 ;
        RECT 108.170 16.840 109.120 17.120 ;
        RECT 108.170 16.670 108.200 16.840 ;
        RECT 108.370 16.670 108.560 16.840 ;
        RECT 108.730 16.670 108.920 16.840 ;
        RECT 109.090 16.670 109.120 16.840 ;
        RECT 108.170 16.640 109.120 16.670 ;
        RECT 109.300 16.710 109.470 17.300 ;
        RECT 109.650 16.890 109.980 17.650 ;
        RECT 111.290 17.420 111.620 18.000 ;
        RECT 111.800 18.590 112.970 18.760 ;
        RECT 111.800 17.240 111.970 18.590 ;
        RECT 112.350 17.910 112.680 18.410 ;
        RECT 113.150 18.160 113.320 19.560 ;
      LAYER li1 ;
        RECT 113.500 19.250 113.670 19.910 ;
      LAYER li1 ;
        RECT 113.850 19.950 114.800 19.980 ;
        RECT 113.850 19.780 113.880 19.950 ;
        RECT 114.050 19.780 114.240 19.950 ;
        RECT 114.410 19.780 114.600 19.950 ;
        RECT 114.770 19.780 114.800 19.950 ;
        RECT 116.460 19.950 117.410 19.980 ;
        RECT 113.850 19.430 114.800 19.780 ;
        RECT 115.340 19.350 115.670 19.850 ;
        RECT 116.460 19.780 116.490 19.950 ;
        RECT 116.660 19.780 116.850 19.950 ;
        RECT 117.020 19.780 117.210 19.950 ;
        RECT 117.380 19.780 117.410 19.950 ;
      LAYER li1 ;
        RECT 113.500 19.140 114.510 19.250 ;
        RECT 113.500 19.080 114.560 19.140 ;
        RECT 114.180 18.970 114.560 19.080 ;
      LAYER li1 ;
        RECT 113.530 18.510 113.860 18.900 ;
      LAYER li1 ;
        RECT 114.180 18.690 114.510 18.970 ;
      LAYER li1 ;
        RECT 115.340 18.510 115.570 19.350 ;
        RECT 115.950 18.850 116.280 19.350 ;
        RECT 116.460 18.850 117.410 19.780 ;
        RECT 118.250 19.950 119.860 19.980 ;
        RECT 118.250 19.780 118.300 19.950 ;
        RECT 118.470 19.780 118.740 19.950 ;
        RECT 118.910 19.780 119.180 19.950 ;
        RECT 119.350 19.780 119.590 19.950 ;
        RECT 119.760 19.780 119.860 19.950 ;
        RECT 121.540 19.950 122.190 20.060 ;
        RECT 113.530 18.340 115.570 18.510 ;
        RECT 112.860 17.990 115.220 18.160 ;
        RECT 112.860 17.670 113.030 17.990 ;
        RECT 115.400 17.810 115.570 18.340 ;
        RECT 110.160 17.070 111.970 17.240 ;
        RECT 112.150 17.500 113.030 17.670 ;
        RECT 110.160 16.710 110.330 17.070 ;
        RECT 109.300 16.540 110.330 16.710 ;
        RECT 110.510 16.840 111.460 16.890 ;
        RECT 110.510 16.670 110.540 16.840 ;
        RECT 110.710 16.670 110.900 16.840 ;
        RECT 111.070 16.670 111.260 16.840 ;
        RECT 111.430 16.670 111.460 16.840 ;
        RECT 110.510 16.590 111.460 16.670 ;
        RECT 112.150 16.590 112.400 17.500 ;
        RECT 113.210 16.840 114.160 17.670 ;
        RECT 114.560 17.640 115.570 17.810 ;
        RECT 116.070 18.670 116.280 18.850 ;
        RECT 116.070 18.340 117.440 18.670 ;
        RECT 114.560 17.170 114.810 17.640 ;
        RECT 114.990 16.840 115.890 17.460 ;
        RECT 116.070 17.340 116.320 18.340 ;
        RECT 113.210 16.670 113.240 16.840 ;
        RECT 113.410 16.670 113.600 16.840 ;
        RECT 113.770 16.670 113.960 16.840 ;
        RECT 114.130 16.670 114.160 16.840 ;
        RECT 115.160 16.670 115.350 16.840 ;
        RECT 115.520 16.670 115.710 16.840 ;
        RECT 115.880 16.670 115.890 16.840 ;
        RECT 113.210 16.640 114.160 16.670 ;
        RECT 114.990 16.640 115.890 16.670 ;
        RECT 116.500 16.840 117.440 18.150 ;
        RECT 116.500 16.670 116.520 16.840 ;
        RECT 116.690 16.670 116.880 16.840 ;
        RECT 117.050 16.670 117.240 16.840 ;
        RECT 117.410 16.670 117.440 16.840 ;
        RECT 116.500 16.610 117.440 16.670 ;
      LAYER li1 ;
        RECT 117.620 16.610 117.960 19.680 ;
      LAYER li1 ;
        RECT 118.250 19.500 119.860 19.780 ;
        RECT 118.560 19.100 119.860 19.500 ;
      LAYER li1 ;
        RECT 120.290 19.280 120.870 19.920 ;
      LAYER li1 ;
        RECT 121.540 19.780 121.600 19.950 ;
        RECT 121.770 19.780 121.960 19.950 ;
        RECT 122.130 19.780 122.190 19.950 ;
        RECT 121.540 19.720 122.190 19.780 ;
        RECT 121.780 19.280 122.190 19.720 ;
        RECT 122.570 19.950 124.180 19.980 ;
        RECT 122.570 19.780 122.620 19.950 ;
        RECT 122.790 19.780 123.060 19.950 ;
        RECT 123.230 19.780 123.500 19.950 ;
        RECT 123.670 19.780 123.910 19.950 ;
        RECT 124.080 19.780 124.180 19.950 ;
        RECT 125.860 19.950 126.510 20.060 ;
        RECT 122.570 19.500 124.180 19.780 ;
        RECT 118.560 18.320 118.890 19.100 ;
        RECT 119.100 17.660 119.430 18.650 ;
      LAYER li1 ;
        RECT 120.620 18.410 120.870 19.280 ;
      LAYER li1 ;
        RECT 122.880 19.100 124.180 19.500 ;
      LAYER li1 ;
        RECT 124.610 19.280 125.190 19.920 ;
      LAYER li1 ;
        RECT 125.860 19.780 125.920 19.950 ;
        RECT 126.090 19.780 126.280 19.950 ;
        RECT 126.450 19.780 126.510 19.950 ;
        RECT 125.860 19.720 126.510 19.780 ;
        RECT 126.100 19.280 126.510 19.720 ;
        RECT 127.300 19.960 130.030 19.990 ;
        RECT 127.300 19.790 127.470 19.960 ;
        RECT 127.640 19.790 127.910 19.960 ;
        RECT 128.080 19.790 128.320 19.960 ;
        RECT 128.490 19.790 128.750 19.960 ;
        RECT 128.920 19.790 129.190 19.960 ;
        RECT 129.360 19.790 129.600 19.960 ;
        RECT 129.770 19.790 130.030 19.960 ;
      LAYER li1 ;
        RECT 120.620 18.160 121.330 18.410 ;
      LAYER li1 ;
        RECT 122.880 18.320 123.210 19.100 ;
        RECT 118.330 16.790 119.780 17.660 ;
        RECT 118.330 16.620 118.580 16.790 ;
        RECT 118.750 16.620 118.940 16.790 ;
        RECT 119.110 16.620 119.380 16.790 ;
        RECT 119.550 16.620 119.780 16.790 ;
        RECT 118.330 16.590 119.780 16.620 ;
        RECT 120.220 16.900 120.620 17.170 ;
        RECT 120.220 16.840 120.870 16.900 ;
        RECT 120.220 16.670 120.280 16.840 ;
        RECT 120.450 16.670 120.640 16.840 ;
        RECT 120.810 16.670 120.870 16.840 ;
      LAYER li1 ;
        RECT 121.080 16.820 121.330 18.160 ;
      LAYER li1 ;
        RECT 123.420 17.660 123.750 18.650 ;
      LAYER li1 ;
        RECT 124.940 18.410 125.190 19.280 ;
      LAYER li1 ;
        RECT 127.300 18.990 130.030 19.790 ;
        RECT 131.140 19.960 133.870 19.990 ;
        RECT 131.140 19.790 131.310 19.960 ;
        RECT 131.480 19.790 131.750 19.960 ;
        RECT 131.920 19.790 132.160 19.960 ;
        RECT 132.330 19.790 132.590 19.960 ;
        RECT 132.760 19.790 133.030 19.960 ;
        RECT 133.200 19.790 133.440 19.960 ;
        RECT 133.610 19.790 133.870 19.960 ;
        RECT 135.940 19.950 136.590 20.060 ;
        RECT 131.140 18.990 133.870 19.790 ;
      LAYER li1 ;
        RECT 134.690 19.280 135.270 19.920 ;
      LAYER li1 ;
        RECT 135.940 19.780 136.000 19.950 ;
        RECT 136.170 19.780 136.360 19.950 ;
        RECT 136.530 19.780 136.590 19.950 ;
        RECT 135.940 19.720 136.590 19.780 ;
        RECT 136.180 19.280 136.590 19.720 ;
        RECT 137.380 19.960 140.110 19.990 ;
        RECT 137.380 19.790 137.550 19.960 ;
        RECT 137.720 19.790 137.990 19.960 ;
        RECT 138.160 19.790 138.400 19.960 ;
        RECT 138.570 19.790 138.830 19.960 ;
        RECT 139.000 19.790 139.270 19.960 ;
        RECT 139.440 19.790 139.680 19.960 ;
        RECT 139.850 19.790 140.110 19.960 ;
      LAYER li1 ;
        RECT 124.940 18.160 125.650 18.410 ;
      LAYER li1 ;
        RECT 127.460 18.320 127.790 18.990 ;
        RECT 120.220 16.560 120.870 16.670 ;
        RECT 122.650 16.790 124.100 17.660 ;
        RECT 122.650 16.620 122.900 16.790 ;
        RECT 123.070 16.620 123.260 16.790 ;
        RECT 123.430 16.620 123.700 16.790 ;
        RECT 123.870 16.620 124.100 16.790 ;
        RECT 122.650 16.590 124.100 16.620 ;
        RECT 124.540 16.900 124.940 17.170 ;
        RECT 124.540 16.840 125.190 16.900 ;
        RECT 124.540 16.670 124.600 16.840 ;
        RECT 124.770 16.670 124.960 16.840 ;
        RECT 125.130 16.670 125.190 16.840 ;
      LAYER li1 ;
        RECT 125.400 16.820 125.650 18.160 ;
      LAYER li1 ;
        RECT 128.190 17.670 128.520 18.650 ;
        RECT 128.740 18.320 129.070 18.990 ;
        RECT 129.470 17.670 129.800 18.650 ;
        RECT 131.300 18.320 131.630 18.990 ;
        RECT 132.030 17.670 132.360 18.650 ;
        RECT 132.580 18.320 132.910 18.990 ;
        RECT 133.310 17.670 133.640 18.650 ;
      LAYER li1 ;
        RECT 135.020 18.410 135.270 19.280 ;
      LAYER li1 ;
        RECT 137.380 18.990 140.110 19.790 ;
      LAYER li1 ;
        RECT 135.020 18.160 135.730 18.410 ;
      LAYER li1 ;
        RECT 137.540 18.320 137.870 18.990 ;
        RECT 124.540 16.560 125.190 16.670 ;
        RECT 127.220 16.790 129.960 17.670 ;
        RECT 127.220 16.620 127.430 16.790 ;
        RECT 127.600 16.620 127.870 16.790 ;
        RECT 128.040 16.620 128.280 16.790 ;
        RECT 128.450 16.620 128.710 16.790 ;
        RECT 128.880 16.620 129.150 16.790 ;
        RECT 129.320 16.620 129.560 16.790 ;
        RECT 129.730 16.620 129.960 16.790 ;
        RECT 127.220 16.600 129.960 16.620 ;
        RECT 131.060 16.790 133.800 17.670 ;
        RECT 131.060 16.620 131.270 16.790 ;
        RECT 131.440 16.620 131.710 16.790 ;
        RECT 131.880 16.620 132.120 16.790 ;
        RECT 132.290 16.620 132.550 16.790 ;
        RECT 132.720 16.620 132.990 16.790 ;
        RECT 133.160 16.620 133.400 16.790 ;
        RECT 133.570 16.620 133.800 16.790 ;
        RECT 131.060 16.600 133.800 16.620 ;
        RECT 134.620 16.900 135.020 17.170 ;
        RECT 134.620 16.840 135.270 16.900 ;
        RECT 134.620 16.670 134.680 16.840 ;
        RECT 134.850 16.670 135.040 16.840 ;
        RECT 135.210 16.670 135.270 16.840 ;
      LAYER li1 ;
        RECT 135.480 16.820 135.730 18.160 ;
      LAYER li1 ;
        RECT 138.270 17.670 138.600 18.650 ;
        RECT 138.820 18.320 139.150 18.990 ;
        RECT 139.550 17.670 139.880 18.650 ;
        RECT 134.620 16.560 135.270 16.670 ;
        RECT 137.300 16.790 140.040 17.670 ;
        RECT 137.300 16.620 137.510 16.790 ;
        RECT 137.680 16.620 137.950 16.790 ;
        RECT 138.120 16.620 138.360 16.790 ;
        RECT 138.530 16.620 138.790 16.790 ;
        RECT 138.960 16.620 139.230 16.790 ;
        RECT 139.400 16.620 139.640 16.790 ;
        RECT 139.810 16.620 140.040 16.790 ;
        RECT 137.300 16.600 140.040 16.620 ;
        RECT 5.760 16.190 5.920 16.360 ;
        RECT 6.090 16.190 6.400 16.360 ;
        RECT 6.570 16.190 6.880 16.360 ;
        RECT 7.050 16.190 7.360 16.360 ;
        RECT 7.530 16.190 7.840 16.360 ;
        RECT 8.010 16.190 8.320 16.360 ;
        RECT 8.490 16.190 8.800 16.360 ;
        RECT 8.970 16.190 9.280 16.360 ;
        RECT 9.450 16.190 9.760 16.360 ;
        RECT 9.930 16.190 10.240 16.360 ;
        RECT 10.410 16.190 10.720 16.360 ;
        RECT 10.890 16.190 11.200 16.360 ;
        RECT 11.370 16.190 11.680 16.360 ;
        RECT 11.850 16.190 12.160 16.360 ;
        RECT 12.330 16.190 12.640 16.360 ;
        RECT 12.810 16.190 13.120 16.360 ;
        RECT 13.290 16.190 13.600 16.360 ;
        RECT 13.770 16.190 14.080 16.360 ;
        RECT 14.250 16.190 14.560 16.360 ;
        RECT 14.730 16.190 15.040 16.360 ;
        RECT 15.210 16.190 15.520 16.360 ;
        RECT 15.690 16.190 16.000 16.360 ;
        RECT 16.170 16.190 16.480 16.360 ;
        RECT 16.650 16.190 16.960 16.360 ;
        RECT 17.130 16.190 17.440 16.360 ;
        RECT 17.610 16.190 17.920 16.360 ;
        RECT 18.090 16.190 18.400 16.360 ;
        RECT 18.570 16.190 18.880 16.360 ;
        RECT 19.050 16.190 19.360 16.360 ;
        RECT 19.530 16.190 19.840 16.360 ;
        RECT 20.010 16.190 20.320 16.360 ;
        RECT 20.490 16.190 20.800 16.360 ;
        RECT 20.970 16.190 21.280 16.360 ;
        RECT 21.450 16.190 21.760 16.360 ;
        RECT 21.930 16.190 22.240 16.360 ;
        RECT 22.410 16.190 22.720 16.360 ;
        RECT 22.890 16.190 23.200 16.360 ;
        RECT 23.370 16.190 23.680 16.360 ;
        RECT 23.850 16.190 24.160 16.360 ;
        RECT 24.330 16.190 24.640 16.360 ;
        RECT 24.810 16.190 25.120 16.360 ;
        RECT 25.290 16.190 25.600 16.360 ;
        RECT 25.770 16.190 26.080 16.360 ;
        RECT 26.250 16.190 26.560 16.360 ;
        RECT 26.730 16.190 27.040 16.360 ;
        RECT 27.210 16.190 27.520 16.360 ;
        RECT 27.690 16.190 28.000 16.360 ;
        RECT 28.170 16.190 28.480 16.360 ;
        RECT 28.650 16.190 28.960 16.360 ;
        RECT 29.130 16.190 29.440 16.360 ;
        RECT 29.610 16.190 29.920 16.360 ;
        RECT 30.090 16.190 30.400 16.360 ;
        RECT 30.570 16.190 30.880 16.360 ;
        RECT 31.050 16.190 31.360 16.360 ;
        RECT 31.530 16.190 31.840 16.360 ;
        RECT 32.010 16.190 32.320 16.360 ;
        RECT 32.490 16.190 32.800 16.360 ;
        RECT 32.970 16.190 33.280 16.360 ;
        RECT 33.450 16.190 33.760 16.360 ;
        RECT 33.930 16.190 34.240 16.360 ;
        RECT 34.410 16.190 34.720 16.360 ;
        RECT 34.890 16.190 35.200 16.360 ;
        RECT 35.370 16.190 35.680 16.360 ;
        RECT 35.850 16.190 36.160 16.360 ;
        RECT 36.330 16.190 36.640 16.360 ;
        RECT 36.810 16.190 37.120 16.360 ;
        RECT 37.290 16.190 37.440 16.360 ;
        RECT 37.920 16.190 38.080 16.360 ;
        RECT 38.250 16.190 38.560 16.360 ;
        RECT 38.730 16.190 39.040 16.360 ;
        RECT 39.210 16.190 39.520 16.360 ;
        RECT 39.690 16.190 40.000 16.360 ;
        RECT 40.170 16.190 40.480 16.360 ;
        RECT 40.650 16.190 40.960 16.360 ;
        RECT 41.130 16.190 41.440 16.360 ;
        RECT 41.610 16.190 41.920 16.360 ;
        RECT 42.090 16.190 42.400 16.360 ;
        RECT 42.570 16.190 42.880 16.360 ;
        RECT 43.050 16.190 43.360 16.360 ;
        RECT 43.530 16.190 43.840 16.360 ;
        RECT 44.010 16.190 44.320 16.360 ;
        RECT 44.490 16.190 44.800 16.360 ;
        RECT 44.970 16.190 45.280 16.360 ;
        RECT 45.450 16.190 45.760 16.360 ;
        RECT 45.930 16.190 46.240 16.360 ;
        RECT 46.410 16.190 46.720 16.360 ;
        RECT 46.890 16.190 47.200 16.360 ;
        RECT 47.370 16.190 47.680 16.360 ;
        RECT 47.850 16.190 48.160 16.360 ;
        RECT 48.330 16.190 48.640 16.360 ;
        RECT 48.810 16.190 49.120 16.360 ;
        RECT 49.290 16.190 49.600 16.360 ;
        RECT 49.770 16.190 50.080 16.360 ;
        RECT 50.250 16.190 50.560 16.360 ;
        RECT 50.730 16.190 51.040 16.360 ;
        RECT 51.210 16.190 51.520 16.360 ;
        RECT 51.690 16.190 52.000 16.360 ;
        RECT 52.170 16.190 52.480 16.360 ;
        RECT 52.650 16.190 52.960 16.360 ;
        RECT 53.130 16.190 53.440 16.360 ;
        RECT 53.610 16.190 53.920 16.360 ;
        RECT 54.090 16.190 54.400 16.360 ;
        RECT 54.570 16.190 54.880 16.360 ;
        RECT 55.050 16.190 55.360 16.360 ;
        RECT 55.530 16.190 55.840 16.360 ;
        RECT 56.010 16.190 56.320 16.360 ;
        RECT 56.490 16.190 56.800 16.360 ;
        RECT 56.970 16.190 57.280 16.360 ;
        RECT 57.450 16.190 57.760 16.360 ;
        RECT 57.930 16.190 58.240 16.360 ;
        RECT 58.410 16.190 58.720 16.360 ;
        RECT 58.890 16.190 59.200 16.360 ;
        RECT 59.370 16.190 59.680 16.360 ;
        RECT 59.850 16.190 60.160 16.360 ;
        RECT 60.330 16.190 60.640 16.360 ;
        RECT 60.810 16.190 61.120 16.360 ;
        RECT 61.290 16.190 61.600 16.360 ;
        RECT 61.770 16.190 62.080 16.360 ;
        RECT 62.250 16.190 62.560 16.360 ;
        RECT 62.730 16.190 63.040 16.360 ;
        RECT 63.210 16.190 63.520 16.360 ;
        RECT 63.690 16.190 64.000 16.360 ;
        RECT 64.170 16.190 64.480 16.360 ;
        RECT 64.650 16.190 64.960 16.360 ;
        RECT 65.130 16.190 65.440 16.360 ;
        RECT 65.610 16.190 65.920 16.360 ;
        RECT 66.090 16.190 66.400 16.360 ;
        RECT 66.570 16.190 66.880 16.360 ;
        RECT 67.050 16.190 67.360 16.360 ;
        RECT 67.530 16.190 67.840 16.360 ;
        RECT 68.010 16.190 68.320 16.360 ;
        RECT 68.490 16.190 68.800 16.360 ;
        RECT 68.970 16.190 69.280 16.360 ;
        RECT 69.450 16.190 69.760 16.360 ;
        RECT 69.930 16.190 70.240 16.360 ;
        RECT 70.410 16.190 70.720 16.360 ;
        RECT 70.890 16.190 71.200 16.360 ;
        RECT 71.370 16.190 71.680 16.360 ;
        RECT 71.850 16.190 72.160 16.360 ;
        RECT 72.330 16.190 72.640 16.360 ;
        RECT 72.810 16.190 73.120 16.360 ;
        RECT 73.290 16.190 73.600 16.360 ;
        RECT 73.770 16.190 74.080 16.360 ;
        RECT 74.250 16.190 74.560 16.360 ;
        RECT 74.730 16.190 75.040 16.360 ;
        RECT 75.210 16.190 75.520 16.360 ;
        RECT 75.690 16.190 76.000 16.360 ;
        RECT 76.170 16.190 76.480 16.360 ;
        RECT 76.650 16.190 76.960 16.360 ;
        RECT 77.130 16.190 77.440 16.360 ;
        RECT 77.610 16.190 77.920 16.360 ;
        RECT 78.090 16.190 78.400 16.360 ;
        RECT 78.570 16.190 78.880 16.360 ;
        RECT 79.050 16.190 79.360 16.360 ;
        RECT 79.530 16.190 79.840 16.360 ;
        RECT 80.010 16.190 80.320 16.360 ;
        RECT 80.490 16.190 80.800 16.360 ;
        RECT 80.970 16.190 81.280 16.360 ;
        RECT 81.450 16.190 81.760 16.360 ;
        RECT 81.930 16.190 82.240 16.360 ;
        RECT 82.410 16.190 82.720 16.360 ;
        RECT 82.890 16.190 83.200 16.360 ;
        RECT 83.370 16.190 83.680 16.360 ;
        RECT 83.850 16.190 84.160 16.360 ;
        RECT 84.330 16.190 84.640 16.360 ;
        RECT 84.810 16.190 85.120 16.360 ;
        RECT 85.290 16.190 85.600 16.360 ;
        RECT 85.770 16.190 86.080 16.360 ;
        RECT 86.250 16.190 86.560 16.360 ;
        RECT 86.730 16.190 87.040 16.360 ;
        RECT 87.210 16.190 87.520 16.360 ;
        RECT 87.690 16.190 88.000 16.360 ;
        RECT 88.170 16.190 88.480 16.360 ;
        RECT 88.650 16.190 88.960 16.360 ;
        RECT 89.130 16.190 89.440 16.360 ;
        RECT 89.610 16.190 89.920 16.360 ;
        RECT 90.090 16.190 90.400 16.360 ;
        RECT 90.570 16.190 90.880 16.360 ;
        RECT 91.050 16.190 91.360 16.360 ;
        RECT 91.530 16.190 91.840 16.360 ;
        RECT 92.010 16.190 92.320 16.360 ;
        RECT 92.490 16.190 92.800 16.360 ;
        RECT 92.970 16.190 93.280 16.360 ;
        RECT 93.450 16.190 93.760 16.360 ;
        RECT 93.930 16.190 94.240 16.360 ;
        RECT 94.410 16.190 94.720 16.360 ;
        RECT 94.890 16.190 95.200 16.360 ;
        RECT 95.370 16.190 95.680 16.360 ;
        RECT 95.850 16.190 96.160 16.360 ;
        RECT 96.330 16.190 96.640 16.360 ;
        RECT 96.810 16.190 97.120 16.360 ;
        RECT 97.290 16.190 97.600 16.360 ;
        RECT 97.770 16.190 98.080 16.360 ;
        RECT 98.250 16.190 98.560 16.360 ;
        RECT 98.730 16.190 99.040 16.360 ;
        RECT 99.210 16.190 99.520 16.360 ;
        RECT 99.690 16.190 100.000 16.360 ;
        RECT 100.170 16.190 100.480 16.360 ;
        RECT 100.650 16.190 100.960 16.360 ;
        RECT 101.130 16.190 101.440 16.360 ;
        RECT 101.610 16.190 101.920 16.360 ;
        RECT 102.090 16.190 102.400 16.360 ;
        RECT 102.570 16.190 102.880 16.360 ;
        RECT 103.050 16.190 103.360 16.360 ;
        RECT 103.530 16.190 103.840 16.360 ;
        RECT 104.010 16.190 104.320 16.360 ;
        RECT 104.490 16.190 104.800 16.360 ;
        RECT 104.970 16.190 105.280 16.360 ;
        RECT 105.450 16.190 105.760 16.360 ;
        RECT 105.930 16.190 106.240 16.360 ;
        RECT 106.410 16.190 106.720 16.360 ;
        RECT 106.890 16.190 107.200 16.360 ;
        RECT 107.370 16.190 107.680 16.360 ;
        RECT 107.850 16.190 108.160 16.360 ;
        RECT 108.330 16.190 108.640 16.360 ;
        RECT 108.810 16.190 109.120 16.360 ;
        RECT 109.290 16.190 109.600 16.360 ;
        RECT 109.770 16.190 110.080 16.360 ;
        RECT 110.250 16.190 110.560 16.360 ;
        RECT 110.730 16.190 111.040 16.360 ;
        RECT 111.210 16.190 111.520 16.360 ;
        RECT 111.690 16.190 112.000 16.360 ;
        RECT 112.170 16.190 112.480 16.360 ;
        RECT 112.650 16.190 112.960 16.360 ;
        RECT 113.130 16.190 113.440 16.360 ;
        RECT 113.610 16.190 113.920 16.360 ;
        RECT 114.090 16.190 114.400 16.360 ;
        RECT 114.570 16.190 114.880 16.360 ;
        RECT 115.050 16.190 115.360 16.360 ;
        RECT 115.530 16.190 115.840 16.360 ;
        RECT 116.010 16.190 116.320 16.360 ;
        RECT 116.490 16.190 116.800 16.360 ;
        RECT 116.970 16.190 117.280 16.360 ;
        RECT 117.450 16.190 117.760 16.360 ;
        RECT 117.930 16.190 118.240 16.360 ;
        RECT 118.410 16.190 118.720 16.360 ;
        RECT 118.890 16.190 119.200 16.360 ;
        RECT 119.370 16.190 119.680 16.360 ;
        RECT 119.850 16.190 120.160 16.360 ;
        RECT 120.330 16.190 120.640 16.360 ;
        RECT 120.810 16.190 121.120 16.360 ;
        RECT 121.290 16.190 121.600 16.360 ;
        RECT 121.770 16.190 122.080 16.360 ;
        RECT 122.250 16.190 122.560 16.360 ;
        RECT 122.730 16.190 123.040 16.360 ;
        RECT 123.210 16.190 123.520 16.360 ;
        RECT 123.690 16.190 124.000 16.360 ;
        RECT 124.170 16.190 124.480 16.360 ;
        RECT 124.650 16.190 124.960 16.360 ;
        RECT 125.130 16.190 125.440 16.360 ;
        RECT 125.610 16.190 125.920 16.360 ;
        RECT 126.090 16.190 126.400 16.360 ;
        RECT 126.570 16.190 126.880 16.360 ;
        RECT 127.050 16.190 127.360 16.360 ;
        RECT 127.530 16.190 127.840 16.360 ;
        RECT 128.010 16.190 128.320 16.360 ;
        RECT 128.490 16.190 128.800 16.360 ;
        RECT 128.970 16.190 129.280 16.360 ;
        RECT 129.450 16.190 129.760 16.360 ;
        RECT 129.930 16.190 130.240 16.360 ;
        RECT 130.410 16.190 130.720 16.360 ;
        RECT 130.890 16.190 131.200 16.360 ;
        RECT 131.370 16.190 131.680 16.360 ;
        RECT 131.850 16.190 132.160 16.360 ;
        RECT 132.330 16.190 132.640 16.360 ;
        RECT 132.810 16.190 133.120 16.360 ;
        RECT 133.290 16.190 133.600 16.360 ;
        RECT 133.770 16.190 134.080 16.360 ;
        RECT 134.250 16.190 134.560 16.360 ;
        RECT 134.730 16.190 135.040 16.360 ;
        RECT 135.210 16.190 135.520 16.360 ;
        RECT 135.690 16.190 136.000 16.360 ;
        RECT 136.170 16.190 136.480 16.360 ;
        RECT 136.650 16.190 136.960 16.360 ;
        RECT 137.130 16.190 137.440 16.360 ;
        RECT 137.610 16.190 137.920 16.360 ;
        RECT 138.090 16.190 138.400 16.360 ;
        RECT 138.570 16.190 138.880 16.360 ;
        RECT 139.050 16.190 139.360 16.360 ;
        RECT 139.530 16.190 139.840 16.360 ;
        RECT 140.010 16.190 140.320 16.360 ;
        RECT 140.490 16.190 140.800 16.360 ;
        RECT 140.970 16.190 141.280 16.360 ;
        RECT 141.450 16.190 141.600 16.360 ;
      LAYER mcon ;
        RECT 6.510 142.840 6.680 143.010 ;
        RECT 6.950 142.840 7.120 143.010 ;
        RECT 7.360 142.840 7.530 143.010 ;
        RECT 7.790 142.840 7.960 143.010 ;
        RECT 8.230 142.840 8.400 143.010 ;
        RECT 8.640 142.840 8.810 143.010 ;
        RECT 12.160 142.850 12.330 143.020 ;
        RECT 12.520 142.850 12.690 143.020 ;
        RECT 13.710 142.840 13.880 143.010 ;
        RECT 14.150 142.840 14.320 143.010 ;
        RECT 14.560 142.840 14.730 143.010 ;
        RECT 14.990 142.840 15.160 143.010 ;
        RECT 15.430 142.840 15.600 143.010 ;
        RECT 15.840 142.840 16.010 143.010 ;
        RECT 18.840 142.850 19.010 143.020 ;
        RECT 19.200 142.850 19.370 143.020 ;
      LAYER L1M1_PR_C ;
        RECT 20.790 144.030 20.960 144.200 ;
      LAYER mcon ;
        RECT 20.710 142.850 20.880 143.020 ;
        RECT 21.070 142.850 21.240 143.020 ;
        RECT 23.130 142.850 23.300 143.020 ;
        RECT 23.490 142.850 23.660 143.020 ;
        RECT 23.850 142.850 24.020 143.020 ;
      LAYER L1M1_PR_C ;
        RECT 28.950 143.290 29.120 143.460 ;
      LAYER mcon ;
        RECT 25.070 142.850 25.240 143.020 ;
        RECT 25.430 142.850 25.600 143.020 ;
        RECT 25.790 142.850 25.960 143.020 ;
        RECT 29.610 142.850 29.780 143.020 ;
        RECT 29.970 142.850 30.140 143.020 ;
        RECT 31.530 142.850 31.700 143.020 ;
        RECT 31.890 142.850 32.060 143.020 ;
        RECT 32.250 142.850 32.420 143.020 ;
        RECT 33.340 142.850 33.510 143.020 ;
        RECT 33.780 142.850 33.950 143.020 ;
        RECT 34.220 142.850 34.390 143.020 ;
        RECT 34.630 142.850 34.800 143.020 ;
      LAYER L1M1_PR_C ;
        RECT 38.070 144.030 38.240 144.200 ;
        RECT 36.630 143.290 36.800 143.460 ;
      LAYER mcon ;
        RECT 37.030 142.850 37.200 143.020 ;
        RECT 37.390 142.850 37.560 143.020 ;
        RECT 37.750 142.850 37.920 143.020 ;
        RECT 38.110 142.850 38.280 143.020 ;
        RECT 39.630 142.840 39.800 143.010 ;
        RECT 40.070 142.840 40.240 143.010 ;
        RECT 40.480 142.840 40.650 143.010 ;
        RECT 40.910 142.840 41.080 143.010 ;
        RECT 41.350 142.840 41.520 143.010 ;
        RECT 41.760 142.840 41.930 143.010 ;
        RECT 45.760 142.850 45.930 143.020 ;
        RECT 46.120 142.850 46.290 143.020 ;
        RECT 47.310 142.840 47.480 143.010 ;
        RECT 47.750 142.840 47.920 143.010 ;
        RECT 48.160 142.840 48.330 143.010 ;
        RECT 48.590 142.840 48.760 143.010 ;
        RECT 49.030 142.840 49.200 143.010 ;
        RECT 49.440 142.840 49.610 143.010 ;
      LAYER L1M1_PR_C ;
        RECT 51.990 144.030 52.160 144.200 ;
        RECT 50.550 143.290 50.720 143.460 ;
      LAYER mcon ;
        RECT 50.950 142.850 51.120 143.020 ;
        RECT 51.310 142.850 51.480 143.020 ;
        RECT 51.670 142.850 51.840 143.020 ;
        RECT 52.030 142.850 52.200 143.020 ;
        RECT 53.550 142.840 53.720 143.010 ;
        RECT 53.990 142.840 54.160 143.010 ;
        RECT 54.400 142.840 54.570 143.010 ;
        RECT 54.830 142.840 55.000 143.010 ;
        RECT 55.270 142.840 55.440 143.010 ;
        RECT 55.680 142.840 55.850 143.010 ;
        RECT 57.390 142.840 57.560 143.010 ;
        RECT 57.830 142.840 58.000 143.010 ;
        RECT 58.240 142.840 58.410 143.010 ;
        RECT 58.670 142.840 58.840 143.010 ;
        RECT 59.110 142.840 59.280 143.010 ;
        RECT 59.520 142.840 59.690 143.010 ;
      LAYER L1M1_PR_C ;
        RECT 61.110 144.030 61.280 144.200 ;
      LAYER mcon ;
        RECT 61.070 142.850 61.240 143.020 ;
        RECT 61.430 142.850 61.600 143.020 ;
        RECT 61.790 142.850 61.960 143.020 ;
        RECT 62.710 142.850 62.880 143.020 ;
        RECT 63.070 142.850 63.240 143.020 ;
      LAYER L1M1_PR_C ;
        RECT 63.990 143.290 64.160 143.460 ;
      LAYER mcon ;
        RECT 67.670 142.850 67.840 143.020 ;
        RECT 68.030 142.850 68.200 143.020 ;
        RECT 68.390 142.850 68.560 143.020 ;
      LAYER L1M1_PR_C ;
        RECT 72.150 143.660 72.320 143.830 ;
      LAYER mcon ;
        RECT 71.640 142.850 71.810 143.020 ;
        RECT 72.000 142.850 72.170 143.020 ;
        RECT 72.360 142.850 72.530 143.020 ;
      LAYER L1M1_PR_C ;
        RECT 77.910 144.030 78.080 144.200 ;
      LAYER mcon ;
        RECT 74.250 142.850 74.420 143.020 ;
        RECT 74.610 142.850 74.780 143.020 ;
        RECT 74.970 142.850 75.140 143.020 ;
        RECT 76.060 142.850 76.230 143.020 ;
        RECT 76.500 142.850 76.670 143.020 ;
        RECT 76.940 142.850 77.110 143.020 ;
        RECT 77.350 142.850 77.520 143.020 ;
        RECT 77.880 142.850 78.050 143.020 ;
        RECT 78.240 142.850 78.410 143.020 ;
        RECT 78.600 142.850 78.770 143.020 ;
        RECT 79.440 142.850 79.610 143.020 ;
        RECT 79.800 142.850 79.970 143.020 ;
        RECT 80.160 142.850 80.330 143.020 ;
        RECT 81.000 142.850 81.170 143.020 ;
        RECT 81.360 142.850 81.530 143.020 ;
        RECT 81.720 142.850 81.890 143.020 ;
        RECT 82.780 142.850 82.950 143.020 ;
        RECT 83.220 142.850 83.390 143.020 ;
        RECT 83.660 142.850 83.830 143.020 ;
        RECT 84.070 142.850 84.240 143.020 ;
      LAYER L1M1_PR_C ;
        RECT 87.510 144.030 87.680 144.200 ;
        RECT 86.070 143.290 86.240 143.460 ;
      LAYER mcon ;
        RECT 86.470 142.850 86.640 143.020 ;
        RECT 86.830 142.850 87.000 143.020 ;
        RECT 87.190 142.850 87.360 143.020 ;
        RECT 87.550 142.850 87.720 143.020 ;
        RECT 89.070 142.840 89.240 143.010 ;
        RECT 89.510 142.840 89.680 143.010 ;
        RECT 89.920 142.840 90.090 143.010 ;
        RECT 90.350 142.840 90.520 143.010 ;
        RECT 90.790 142.840 90.960 143.010 ;
        RECT 91.200 142.840 91.370 143.010 ;
        RECT 92.910 142.840 93.080 143.010 ;
        RECT 93.350 142.840 93.520 143.010 ;
        RECT 93.760 142.840 93.930 143.010 ;
        RECT 94.190 142.840 94.360 143.010 ;
        RECT 94.630 142.840 94.800 143.010 ;
        RECT 95.040 142.840 95.210 143.010 ;
        RECT 96.220 142.850 96.390 143.020 ;
        RECT 96.660 142.850 96.830 143.020 ;
        RECT 97.100 142.850 97.270 143.020 ;
        RECT 97.510 142.850 97.680 143.020 ;
      LAYER L1M1_PR_C ;
        RECT 99.510 144.030 99.680 144.200 ;
        RECT 98.070 143.290 98.240 143.460 ;
      LAYER mcon ;
        RECT 98.470 142.850 98.640 143.020 ;
        RECT 98.830 142.850 99.000 143.020 ;
        RECT 99.190 142.850 99.360 143.020 ;
        RECT 99.550 142.850 99.720 143.020 ;
        RECT 100.540 142.850 100.710 143.020 ;
        RECT 100.980 142.850 101.150 143.020 ;
        RECT 101.420 142.850 101.590 143.020 ;
        RECT 101.830 142.850 102.000 143.020 ;
        RECT 102.790 142.850 102.960 143.020 ;
        RECT 103.150 142.850 103.320 143.020 ;
        RECT 103.510 142.850 103.680 143.020 ;
        RECT 103.870 142.850 104.040 143.020 ;
      LAYER L1M1_PR_C ;
        RECT 108.150 144.770 108.320 144.940 ;
      LAYER mcon ;
        RECT 104.860 142.850 105.030 143.020 ;
        RECT 105.300 142.850 105.470 143.020 ;
        RECT 105.740 142.850 105.910 143.020 ;
        RECT 106.150 142.850 106.320 143.020 ;
      LAYER L1M1_PR_C ;
        RECT 106.710 143.290 106.880 143.460 ;
      LAYER mcon ;
        RECT 107.110 142.850 107.280 143.020 ;
        RECT 107.470 142.850 107.640 143.020 ;
        RECT 107.830 142.850 108.000 143.020 ;
        RECT 108.190 142.850 108.360 143.020 ;
        RECT 109.710 142.840 109.880 143.010 ;
        RECT 110.150 142.840 110.320 143.010 ;
        RECT 110.560 142.840 110.730 143.010 ;
        RECT 110.990 142.840 111.160 143.010 ;
        RECT 111.430 142.840 111.600 143.010 ;
        RECT 111.840 142.840 112.010 143.010 ;
        RECT 113.550 142.840 113.720 143.010 ;
        RECT 113.990 142.840 114.160 143.010 ;
        RECT 114.400 142.840 114.570 143.010 ;
        RECT 114.830 142.840 115.000 143.010 ;
        RECT 115.270 142.840 115.440 143.010 ;
        RECT 115.680 142.840 115.850 143.010 ;
        RECT 117.390 142.840 117.560 143.010 ;
        RECT 117.830 142.840 118.000 143.010 ;
        RECT 118.240 142.840 118.410 143.010 ;
        RECT 118.670 142.840 118.840 143.010 ;
        RECT 119.110 142.840 119.280 143.010 ;
        RECT 119.520 142.840 119.690 143.010 ;
        RECT 121.230 142.840 121.400 143.010 ;
        RECT 121.670 142.840 121.840 143.010 ;
        RECT 122.080 142.840 122.250 143.010 ;
        RECT 122.510 142.840 122.680 143.010 ;
        RECT 122.950 142.840 123.120 143.010 ;
        RECT 123.360 142.840 123.530 143.010 ;
        RECT 124.540 142.850 124.710 143.020 ;
        RECT 124.980 142.850 125.150 143.020 ;
        RECT 125.420 142.850 125.590 143.020 ;
        RECT 125.830 142.850 126.000 143.020 ;
        RECT 128.800 142.850 128.970 143.020 ;
        RECT 129.160 142.850 129.330 143.020 ;
        RECT 130.350 142.840 130.520 143.010 ;
        RECT 130.790 142.840 130.960 143.010 ;
        RECT 131.200 142.840 131.370 143.010 ;
        RECT 131.630 142.840 131.800 143.010 ;
        RECT 132.070 142.840 132.240 143.010 ;
        RECT 132.480 142.840 132.650 143.010 ;
        RECT 133.990 142.850 134.160 143.020 ;
        RECT 134.350 142.850 134.520 143.020 ;
        RECT 134.710 142.850 134.880 143.020 ;
        RECT 135.070 142.850 135.240 143.020 ;
        RECT 136.590 142.840 136.760 143.010 ;
        RECT 137.030 142.840 137.200 143.010 ;
        RECT 137.440 142.840 137.610 143.010 ;
        RECT 137.870 142.840 138.040 143.010 ;
        RECT 138.310 142.840 138.480 143.010 ;
        RECT 138.720 142.840 138.890 143.010 ;
        RECT 139.900 142.850 140.070 143.020 ;
        RECT 140.340 142.850 140.510 143.020 ;
        RECT 140.780 142.850 140.950 143.020 ;
        RECT 141.190 142.850 141.360 143.020 ;
      LAYER L1M1_PR_C ;
        RECT 33.750 140.700 33.920 140.870 ;
        RECT 51.030 140.700 51.200 140.870 ;
        RECT 64.950 141.440 65.120 141.610 ;
        RECT 71.670 140.700 71.840 140.870 ;
        RECT 66.390 139.220 66.560 139.390 ;
        RECT 74.550 140.330 74.720 140.500 ;
        RECT 72.150 139.590 72.320 139.760 ;
        RECT 79.350 140.330 79.520 140.500 ;
        RECT 75.990 139.220 76.160 139.390 ;
        RECT 82.230 140.700 82.400 140.870 ;
        RECT 98.550 141.070 98.720 141.240 ;
        RECT 93.750 139.220 93.920 139.390 ;
        RECT 101.430 140.700 101.600 140.870 ;
        RECT 109.590 141.070 109.760 141.240 ;
        RECT 112.950 139.220 113.120 139.390 ;
        RECT 30.870 136.630 31.040 136.800 ;
      LAYER mcon ;
        RECT 6.510 134.700 6.680 134.870 ;
        RECT 6.950 134.700 7.120 134.870 ;
        RECT 7.360 134.700 7.530 134.870 ;
        RECT 7.790 134.700 7.960 134.870 ;
        RECT 8.230 134.700 8.400 134.870 ;
        RECT 8.640 134.700 8.810 134.870 ;
        RECT 9.820 134.710 9.990 134.880 ;
        RECT 10.260 134.710 10.430 134.880 ;
        RECT 10.700 134.710 10.870 134.880 ;
        RECT 11.110 134.710 11.280 134.880 ;
        RECT 13.030 134.710 13.200 134.880 ;
        RECT 13.390 134.710 13.560 134.880 ;
        RECT 13.750 134.710 13.920 134.880 ;
        RECT 14.110 134.710 14.280 134.880 ;
        RECT 15.630 134.700 15.800 134.870 ;
        RECT 16.070 134.700 16.240 134.870 ;
        RECT 16.480 134.700 16.650 134.870 ;
        RECT 16.910 134.700 17.080 134.870 ;
        RECT 17.350 134.700 17.520 134.870 ;
        RECT 17.760 134.700 17.930 134.870 ;
        RECT 19.470 134.700 19.640 134.870 ;
        RECT 19.910 134.700 20.080 134.870 ;
        RECT 20.320 134.700 20.490 134.870 ;
        RECT 20.750 134.700 20.920 134.870 ;
        RECT 21.190 134.700 21.360 134.870 ;
        RECT 21.600 134.700 21.770 134.870 ;
        RECT 23.310 134.700 23.480 134.870 ;
        RECT 23.750 134.700 23.920 134.870 ;
        RECT 24.160 134.700 24.330 134.870 ;
        RECT 24.590 134.700 24.760 134.870 ;
        RECT 25.030 134.700 25.200 134.870 ;
        RECT 25.440 134.700 25.610 134.870 ;
        RECT 27.150 134.700 27.320 134.870 ;
        RECT 27.590 134.700 27.760 134.870 ;
        RECT 28.000 134.700 28.170 134.870 ;
        RECT 28.430 134.700 28.600 134.870 ;
        RECT 28.870 134.700 29.040 134.870 ;
        RECT 29.280 134.700 29.450 134.870 ;
      LAYER L1M1_PR_C ;
        RECT 32.310 136.260 32.480 136.430 ;
      LAYER mcon ;
        RECT 31.270 134.710 31.440 134.880 ;
        RECT 31.630 134.710 31.800 134.880 ;
        RECT 31.990 134.710 32.160 134.880 ;
        RECT 32.350 134.710 32.520 134.880 ;
        RECT 33.340 134.710 33.510 134.880 ;
        RECT 33.780 134.710 33.950 134.880 ;
        RECT 34.220 134.710 34.390 134.880 ;
        RECT 34.630 134.710 34.800 134.880 ;
        RECT 35.160 134.710 35.330 134.880 ;
        RECT 35.520 134.710 35.690 134.880 ;
      LAYER L1M1_PR_C ;
        RECT 36.150 135.150 36.320 135.320 ;
      LAYER mcon ;
        RECT 37.230 134.700 37.400 134.870 ;
        RECT 37.670 134.700 37.840 134.870 ;
        RECT 38.080 134.700 38.250 134.870 ;
        RECT 38.510 134.700 38.680 134.870 ;
        RECT 38.950 134.700 39.120 134.870 ;
        RECT 39.360 134.700 39.530 134.870 ;
        RECT 41.070 134.700 41.240 134.870 ;
        RECT 41.510 134.700 41.680 134.870 ;
        RECT 41.920 134.700 42.090 134.870 ;
        RECT 42.350 134.700 42.520 134.870 ;
        RECT 42.790 134.700 42.960 134.870 ;
        RECT 43.200 134.700 43.370 134.870 ;
        RECT 44.910 134.700 45.080 134.870 ;
        RECT 45.350 134.700 45.520 134.870 ;
        RECT 45.760 134.700 45.930 134.870 ;
        RECT 46.190 134.700 46.360 134.870 ;
        RECT 46.630 134.700 46.800 134.870 ;
        RECT 47.040 134.700 47.210 134.870 ;
        RECT 48.750 134.700 48.920 134.870 ;
        RECT 49.190 134.700 49.360 134.870 ;
        RECT 49.600 134.700 49.770 134.870 ;
        RECT 50.030 134.700 50.200 134.870 ;
        RECT 50.470 134.700 50.640 134.870 ;
        RECT 50.880 134.700 51.050 134.870 ;
        RECT 52.590 134.700 52.760 134.870 ;
        RECT 53.030 134.700 53.200 134.870 ;
        RECT 53.440 134.700 53.610 134.870 ;
        RECT 53.870 134.700 54.040 134.870 ;
        RECT 54.310 134.700 54.480 134.870 ;
        RECT 54.720 134.700 54.890 134.870 ;
      LAYER L1M1_PR_C ;
        RECT 63.990 137.370 64.160 137.540 ;
      LAYER mcon ;
        RECT 56.430 134.700 56.600 134.870 ;
        RECT 56.870 134.700 57.040 134.870 ;
        RECT 57.280 134.700 57.450 134.870 ;
        RECT 57.710 134.700 57.880 134.870 ;
        RECT 58.150 134.700 58.320 134.870 ;
        RECT 58.560 134.700 58.730 134.870 ;
        RECT 59.740 134.710 59.910 134.880 ;
        RECT 60.180 134.710 60.350 134.880 ;
        RECT 60.620 134.710 60.790 134.880 ;
        RECT 61.030 134.710 61.200 134.880 ;
        RECT 63.000 134.710 63.170 134.880 ;
        RECT 63.360 134.710 63.530 134.880 ;
        RECT 65.070 134.700 65.240 134.870 ;
        RECT 65.510 134.700 65.680 134.870 ;
        RECT 65.920 134.700 66.090 134.870 ;
        RECT 66.350 134.700 66.520 134.870 ;
        RECT 66.790 134.700 66.960 134.870 ;
        RECT 67.200 134.700 67.370 134.870 ;
      LAYER L1M1_PR_C ;
        RECT 76.950 136.630 77.120 136.800 ;
        RECT 77.910 136.260 78.080 136.430 ;
        RECT 75.510 135.890 75.680 136.060 ;
        RECT 78.390 136.260 78.560 136.430 ;
        RECT 76.470 135.890 76.640 136.060 ;
      LAYER mcon ;
        RECT 68.910 134.700 69.080 134.870 ;
        RECT 69.350 134.700 69.520 134.870 ;
        RECT 69.760 134.700 69.930 134.870 ;
        RECT 70.190 134.700 70.360 134.870 ;
        RECT 70.630 134.700 70.800 134.870 ;
        RECT 71.040 134.700 71.210 134.870 ;
        RECT 72.220 134.710 72.390 134.880 ;
        RECT 72.660 134.710 72.830 134.880 ;
        RECT 73.100 134.710 73.270 134.880 ;
        RECT 73.510 134.710 73.680 134.880 ;
        RECT 77.560 134.710 77.730 134.880 ;
        RECT 77.920 134.710 78.090 134.880 ;
        RECT 78.280 134.710 78.450 134.880 ;
      LAYER L1M1_PR_C ;
        RECT 87.030 136.630 87.200 136.800 ;
      LAYER mcon ;
        RECT 79.950 134.700 80.120 134.870 ;
        RECT 80.390 134.700 80.560 134.870 ;
        RECT 80.800 134.700 80.970 134.870 ;
        RECT 81.230 134.700 81.400 134.870 ;
        RECT 81.670 134.700 81.840 134.870 ;
        RECT 82.080 134.700 82.250 134.870 ;
        RECT 83.790 134.700 83.960 134.870 ;
        RECT 84.230 134.700 84.400 134.870 ;
        RECT 84.640 134.700 84.810 134.870 ;
        RECT 85.070 134.700 85.240 134.870 ;
        RECT 85.510 134.700 85.680 134.870 ;
        RECT 85.920 134.700 86.090 134.870 ;
      LAYER L1M1_PR_C ;
        RECT 89.430 136.260 89.600 136.430 ;
        RECT 89.910 135.890 90.080 136.060 ;
        RECT 90.870 135.890 91.040 136.060 ;
        RECT 90.390 135.520 90.560 135.690 ;
      LAYER mcon ;
        RECT 87.440 134.710 87.610 134.880 ;
        RECT 87.800 134.710 87.970 134.880 ;
        RECT 88.160 134.710 88.330 134.880 ;
        RECT 90.800 134.710 90.970 134.880 ;
        RECT 91.160 134.710 91.330 134.880 ;
        RECT 91.520 134.710 91.690 134.880 ;
        RECT 91.880 134.710 92.050 134.880 ;
      LAYER L1M1_PR_C ;
        RECT 98.550 136.630 98.720 136.800 ;
      LAYER mcon ;
        RECT 92.910 134.700 93.080 134.870 ;
        RECT 93.350 134.700 93.520 134.870 ;
        RECT 93.760 134.700 93.930 134.870 ;
        RECT 94.190 134.700 94.360 134.870 ;
        RECT 94.630 134.700 94.800 134.870 ;
        RECT 95.040 134.700 95.210 134.870 ;
        RECT 96.220 134.710 96.390 134.880 ;
        RECT 96.660 134.710 96.830 134.880 ;
        RECT 97.100 134.710 97.270 134.880 ;
        RECT 97.510 134.710 97.680 134.880 ;
      LAYER L1M1_PR_C ;
        RECT 100.950 136.260 101.120 136.430 ;
        RECT 101.430 135.890 101.600 136.060 ;
        RECT 101.910 135.890 102.080 136.060 ;
      LAYER mcon ;
        RECT 98.960 134.710 99.130 134.880 ;
        RECT 99.320 134.710 99.490 134.880 ;
        RECT 99.680 134.710 99.850 134.880 ;
        RECT 102.320 134.710 102.490 134.880 ;
        RECT 102.680 134.710 102.850 134.880 ;
        RECT 103.040 134.710 103.210 134.880 ;
        RECT 103.400 134.710 103.570 134.880 ;
      LAYER L1M1_PR_C ;
        RECT 110.070 136.630 110.240 136.800 ;
      LAYER mcon ;
        RECT 104.430 134.700 104.600 134.870 ;
        RECT 104.870 134.700 105.040 134.870 ;
        RECT 105.280 134.700 105.450 134.870 ;
        RECT 105.710 134.700 105.880 134.870 ;
        RECT 106.150 134.700 106.320 134.870 ;
        RECT 106.560 134.700 106.730 134.870 ;
        RECT 107.740 134.710 107.910 134.880 ;
        RECT 108.180 134.710 108.350 134.880 ;
        RECT 108.620 134.710 108.790 134.880 ;
        RECT 109.030 134.710 109.200 134.880 ;
      LAYER L1M1_PR_C ;
        RECT 111.510 135.890 111.680 136.060 ;
      LAYER mcon ;
        RECT 110.470 134.710 110.640 134.880 ;
        RECT 110.830 134.710 111.000 134.880 ;
        RECT 111.190 134.710 111.360 134.880 ;
        RECT 111.550 134.710 111.720 134.880 ;
        RECT 113.070 134.700 113.240 134.870 ;
        RECT 113.510 134.700 113.680 134.870 ;
        RECT 113.920 134.700 114.090 134.870 ;
        RECT 114.350 134.700 114.520 134.870 ;
        RECT 114.790 134.700 114.960 134.870 ;
        RECT 115.200 134.700 115.370 134.870 ;
        RECT 116.380 134.710 116.550 134.880 ;
        RECT 116.820 134.710 116.990 134.880 ;
        RECT 117.260 134.710 117.430 134.880 ;
        RECT 117.670 134.710 117.840 134.880 ;
      LAYER L1M1_PR_C ;
        RECT 119.670 135.890 119.840 136.060 ;
        RECT 118.230 135.150 118.400 135.320 ;
      LAYER mcon ;
        RECT 118.630 134.710 118.800 134.880 ;
        RECT 118.990 134.710 119.160 134.880 ;
        RECT 119.350 134.710 119.520 134.880 ;
        RECT 119.710 134.710 119.880 134.880 ;
        RECT 121.230 134.700 121.400 134.870 ;
        RECT 121.670 134.700 121.840 134.870 ;
        RECT 122.080 134.700 122.250 134.870 ;
        RECT 122.510 134.700 122.680 134.870 ;
        RECT 122.950 134.700 123.120 134.870 ;
        RECT 123.360 134.700 123.530 134.870 ;
        RECT 125.070 134.700 125.240 134.870 ;
        RECT 125.510 134.700 125.680 134.870 ;
        RECT 125.920 134.700 126.090 134.870 ;
        RECT 126.350 134.700 126.520 134.870 ;
        RECT 126.790 134.700 126.960 134.870 ;
        RECT 127.200 134.700 127.370 134.870 ;
        RECT 128.910 134.700 129.080 134.870 ;
        RECT 129.350 134.700 129.520 134.870 ;
        RECT 129.760 134.700 129.930 134.870 ;
        RECT 130.190 134.700 130.360 134.870 ;
        RECT 130.630 134.700 130.800 134.870 ;
        RECT 131.040 134.700 131.210 134.870 ;
        RECT 132.750 134.700 132.920 134.870 ;
        RECT 133.190 134.700 133.360 134.870 ;
        RECT 133.600 134.700 133.770 134.870 ;
        RECT 134.030 134.700 134.200 134.870 ;
        RECT 134.470 134.700 134.640 134.870 ;
        RECT 134.880 134.700 135.050 134.870 ;
        RECT 136.590 134.700 136.760 134.870 ;
        RECT 137.030 134.700 137.200 134.870 ;
        RECT 137.440 134.700 137.610 134.870 ;
        RECT 137.870 134.700 138.040 134.870 ;
        RECT 138.310 134.700 138.480 134.870 ;
        RECT 138.720 134.700 138.890 134.870 ;
        RECT 139.900 134.710 140.070 134.880 ;
        RECT 140.340 134.710 140.510 134.880 ;
        RECT 140.780 134.710 140.950 134.880 ;
        RECT 141.190 134.710 141.360 134.880 ;
      LAYER L1M1_PR_C ;
        RECT 32.790 133.300 32.960 133.470 ;
        RECT 31.830 132.560 32.000 132.730 ;
        RECT 32.790 132.560 32.960 132.730 ;
        RECT 34.230 132.190 34.400 132.360 ;
        RECT 35.190 132.190 35.360 132.360 ;
        RECT 74.550 132.930 74.720 133.100 ;
        RECT 78.870 132.190 79.040 132.360 ;
        RECT 79.350 132.190 79.520 132.360 ;
        RECT 76.470 131.080 76.640 131.250 ;
        RECT 80.790 131.450 80.960 131.620 ;
        RECT 85.110 133.300 85.280 133.470 ;
        RECT 81.270 131.080 81.440 131.250 ;
        RECT 87.510 132.190 87.680 132.360 ;
        RECT 88.950 132.560 89.120 132.730 ;
        RECT 87.990 132.190 88.160 132.360 ;
        RECT 98.070 131.820 98.240 131.990 ;
        RECT 100.470 132.190 100.640 132.360 ;
        RECT 101.430 132.560 101.600 132.730 ;
        RECT 100.950 132.190 101.120 132.360 ;
        RECT 107.670 133.300 107.840 133.470 ;
        RECT 105.750 132.560 105.920 132.730 ;
        RECT 106.230 132.560 106.400 132.730 ;
        RECT 107.670 132.190 107.840 132.360 ;
        RECT 111.510 132.190 111.680 132.360 ;
        RECT 114.390 132.560 114.560 132.730 ;
        RECT 125.910 132.930 126.080 133.100 ;
      LAYER mcon ;
        RECT 6.510 126.560 6.680 126.730 ;
        RECT 6.950 126.560 7.120 126.730 ;
        RECT 7.360 126.560 7.530 126.730 ;
        RECT 7.790 126.560 7.960 126.730 ;
        RECT 8.230 126.560 8.400 126.730 ;
        RECT 8.640 126.560 8.810 126.730 ;
        RECT 10.350 126.560 10.520 126.730 ;
        RECT 10.790 126.560 10.960 126.730 ;
        RECT 11.200 126.560 11.370 126.730 ;
        RECT 11.630 126.560 11.800 126.730 ;
        RECT 12.070 126.560 12.240 126.730 ;
        RECT 12.480 126.560 12.650 126.730 ;
        RECT 13.660 126.570 13.830 126.740 ;
        RECT 14.100 126.570 14.270 126.740 ;
        RECT 14.540 126.570 14.710 126.740 ;
        RECT 14.950 126.570 15.120 126.740 ;
      LAYER L1M1_PR_C ;
        RECT 16.950 127.750 17.120 127.920 ;
        RECT 34.710 129.230 34.880 129.400 ;
        RECT 15.510 127.010 15.680 127.180 ;
      LAYER mcon ;
        RECT 15.910 126.570 16.080 126.740 ;
        RECT 16.270 126.570 16.440 126.740 ;
        RECT 16.630 126.570 16.800 126.740 ;
        RECT 16.990 126.570 17.160 126.740 ;
        RECT 18.510 126.560 18.680 126.730 ;
        RECT 18.950 126.560 19.120 126.730 ;
        RECT 19.360 126.560 19.530 126.730 ;
        RECT 19.790 126.560 19.960 126.730 ;
        RECT 20.230 126.560 20.400 126.730 ;
        RECT 20.640 126.560 20.810 126.730 ;
        RECT 22.350 126.560 22.520 126.730 ;
        RECT 22.790 126.560 22.960 126.730 ;
        RECT 23.200 126.560 23.370 126.730 ;
        RECT 23.630 126.560 23.800 126.730 ;
        RECT 24.070 126.560 24.240 126.730 ;
        RECT 24.480 126.560 24.650 126.730 ;
        RECT 26.190 126.560 26.360 126.730 ;
        RECT 26.630 126.560 26.800 126.730 ;
        RECT 27.040 126.560 27.210 126.730 ;
        RECT 27.470 126.560 27.640 126.730 ;
        RECT 27.910 126.560 28.080 126.730 ;
        RECT 28.320 126.560 28.490 126.730 ;
        RECT 30.030 126.560 30.200 126.730 ;
        RECT 30.470 126.560 30.640 126.730 ;
        RECT 30.880 126.560 31.050 126.730 ;
        RECT 31.310 126.560 31.480 126.730 ;
        RECT 31.750 126.560 31.920 126.730 ;
        RECT 32.160 126.560 32.330 126.730 ;
      LAYER L1M1_PR_C ;
        RECT 36.630 129.230 36.800 129.400 ;
      LAYER mcon ;
        RECT 35.160 126.570 35.330 126.740 ;
        RECT 35.520 126.570 35.690 126.740 ;
        RECT 35.880 126.570 36.050 126.740 ;
        RECT 36.240 126.570 36.410 126.740 ;
        RECT 36.600 126.570 36.770 126.740 ;
      LAYER L1M1_PR_C ;
        RECT 39.510 127.750 39.680 127.920 ;
        RECT 45.750 128.120 45.920 128.290 ;
        RECT 46.710 128.120 46.880 128.290 ;
        RECT 44.310 127.750 44.480 127.920 ;
        RECT 47.670 128.120 47.840 128.290 ;
        RECT 45.270 127.750 45.440 127.920 ;
      LAYER mcon ;
        RECT 38.410 126.570 38.580 126.740 ;
        RECT 38.770 126.570 38.940 126.740 ;
        RECT 39.130 126.570 39.300 126.740 ;
        RECT 39.490 126.570 39.660 126.740 ;
        RECT 40.590 126.560 40.760 126.730 ;
        RECT 41.030 126.560 41.200 126.730 ;
        RECT 41.440 126.560 41.610 126.730 ;
        RECT 41.870 126.560 42.040 126.730 ;
        RECT 42.310 126.560 42.480 126.730 ;
        RECT 42.720 126.560 42.890 126.730 ;
        RECT 46.360 126.570 46.530 126.740 ;
        RECT 46.720 126.570 46.890 126.740 ;
        RECT 47.080 126.570 47.250 126.740 ;
        RECT 48.220 126.570 48.390 126.740 ;
        RECT 48.660 126.570 48.830 126.740 ;
        RECT 49.100 126.570 49.270 126.740 ;
        RECT 49.510 126.570 49.680 126.740 ;
        RECT 50.520 126.570 50.690 126.740 ;
        RECT 50.880 126.570 51.050 126.740 ;
      LAYER L1M1_PR_C ;
        RECT 52.470 127.750 52.640 127.920 ;
      LAYER mcon ;
        RECT 52.390 126.570 52.560 126.740 ;
        RECT 52.750 126.570 52.920 126.740 ;
        RECT 54.810 126.570 54.980 126.740 ;
        RECT 55.170 126.570 55.340 126.740 ;
        RECT 55.530 126.570 55.700 126.740 ;
      LAYER L1M1_PR_C ;
        RECT 58.230 127.010 58.400 127.180 ;
      LAYER mcon ;
        RECT 56.750 126.570 56.920 126.740 ;
        RECT 57.110 126.570 57.280 126.740 ;
        RECT 57.470 126.570 57.640 126.740 ;
        RECT 61.290 126.570 61.460 126.740 ;
        RECT 61.650 126.570 61.820 126.740 ;
        RECT 63.210 126.570 63.380 126.740 ;
        RECT 63.570 126.570 63.740 126.740 ;
        RECT 63.930 126.570 64.100 126.740 ;
        RECT 65.020 126.570 65.190 126.740 ;
        RECT 65.460 126.570 65.630 126.740 ;
        RECT 65.900 126.570 66.070 126.740 ;
        RECT 66.310 126.570 66.480 126.740 ;
        RECT 67.800 126.570 67.970 126.740 ;
        RECT 68.160 126.570 68.330 126.740 ;
      LAYER L1M1_PR_C ;
        RECT 68.790 127.380 68.960 127.550 ;
      LAYER mcon ;
        RECT 69.870 126.560 70.040 126.730 ;
        RECT 70.310 126.560 70.480 126.730 ;
        RECT 70.720 126.560 70.890 126.730 ;
        RECT 71.150 126.560 71.320 126.730 ;
        RECT 71.590 126.560 71.760 126.730 ;
        RECT 72.000 126.560 72.170 126.730 ;
      LAYER L1M1_PR_C ;
        RECT 75.510 127.750 75.680 127.920 ;
        RECT 78.390 127.750 78.560 127.920 ;
        RECT 74.550 127.010 74.720 127.180 ;
      LAYER mcon ;
        RECT 75.040 126.570 75.210 126.740 ;
        RECT 75.400 126.570 75.570 126.740 ;
        RECT 75.760 126.570 75.930 126.740 ;
        RECT 76.120 126.570 76.290 126.740 ;
        RECT 76.480 126.570 76.650 126.740 ;
      LAYER L1M1_PR_C ;
        RECT 82.230 128.120 82.400 128.290 ;
        RECT 82.710 128.120 82.880 128.290 ;
        RECT 83.190 129.230 83.360 129.400 ;
        RECT 80.790 127.750 80.960 127.920 ;
        RECT 97.590 129.230 97.760 129.400 ;
      LAYER mcon ;
        RECT 77.290 126.570 77.460 126.740 ;
        RECT 77.650 126.570 77.820 126.740 ;
        RECT 78.010 126.570 78.180 126.740 ;
        RECT 78.370 126.570 78.540 126.740 ;
        RECT 78.940 126.570 79.110 126.740 ;
        RECT 79.380 126.570 79.550 126.740 ;
        RECT 79.820 126.570 79.990 126.740 ;
        RECT 80.230 126.570 80.400 126.740 ;
        RECT 80.760 126.570 80.930 126.740 ;
        RECT 81.120 126.570 81.290 126.740 ;
        RECT 82.030 126.570 82.200 126.740 ;
        RECT 82.390 126.570 82.560 126.740 ;
        RECT 82.750 126.570 82.920 126.740 ;
        RECT 84.750 126.560 84.920 126.730 ;
        RECT 85.190 126.560 85.360 126.730 ;
        RECT 85.600 126.560 85.770 126.730 ;
        RECT 86.030 126.560 86.200 126.730 ;
        RECT 86.470 126.560 86.640 126.730 ;
        RECT 86.880 126.560 87.050 126.730 ;
        RECT 88.590 126.560 88.760 126.730 ;
        RECT 89.030 126.560 89.200 126.730 ;
        RECT 89.440 126.560 89.610 126.730 ;
        RECT 89.870 126.560 90.040 126.730 ;
        RECT 90.310 126.560 90.480 126.730 ;
        RECT 90.720 126.560 90.890 126.730 ;
        RECT 92.430 126.560 92.600 126.730 ;
        RECT 92.870 126.560 93.040 126.730 ;
        RECT 93.280 126.560 93.450 126.730 ;
        RECT 93.710 126.560 93.880 126.730 ;
        RECT 94.150 126.560 94.320 126.730 ;
        RECT 94.560 126.560 94.730 126.730 ;
        RECT 95.740 126.570 95.910 126.740 ;
        RECT 96.180 126.570 96.350 126.740 ;
        RECT 96.620 126.570 96.790 126.740 ;
        RECT 97.030 126.570 97.200 126.740 ;
      LAYER L1M1_PR_C ;
        RECT 99.030 128.120 99.200 128.290 ;
        RECT 99.990 128.120 100.160 128.290 ;
        RECT 100.470 128.120 100.640 128.290 ;
        RECT 100.950 127.750 101.120 127.920 ;
        RECT 112.470 129.230 112.640 129.400 ;
      LAYER mcon ;
        RECT 98.000 126.570 98.170 126.740 ;
        RECT 98.360 126.570 98.530 126.740 ;
        RECT 98.720 126.570 98.890 126.740 ;
        RECT 101.360 126.570 101.530 126.740 ;
        RECT 101.720 126.570 101.890 126.740 ;
        RECT 102.080 126.570 102.250 126.740 ;
        RECT 102.440 126.570 102.610 126.740 ;
        RECT 103.470 126.560 103.640 126.730 ;
        RECT 103.910 126.560 104.080 126.730 ;
        RECT 104.320 126.560 104.490 126.730 ;
        RECT 104.750 126.560 104.920 126.730 ;
        RECT 105.190 126.560 105.360 126.730 ;
        RECT 105.600 126.560 105.770 126.730 ;
        RECT 107.310 126.560 107.480 126.730 ;
        RECT 107.750 126.560 107.920 126.730 ;
        RECT 108.160 126.560 108.330 126.730 ;
        RECT 108.590 126.560 108.760 126.730 ;
        RECT 109.030 126.560 109.200 126.730 ;
        RECT 109.440 126.560 109.610 126.730 ;
      LAYER L1M1_PR_C ;
        RECT 111.030 127.010 111.200 127.180 ;
      LAYER mcon ;
        RECT 111.430 126.570 111.600 126.740 ;
        RECT 111.790 126.570 111.960 126.740 ;
        RECT 112.150 126.570 112.320 126.740 ;
        RECT 112.510 126.570 112.680 126.740 ;
        RECT 114.030 126.560 114.200 126.730 ;
        RECT 114.470 126.560 114.640 126.730 ;
        RECT 114.880 126.560 115.050 126.730 ;
        RECT 115.310 126.560 115.480 126.730 ;
        RECT 115.750 126.560 115.920 126.730 ;
        RECT 116.160 126.560 116.330 126.730 ;
      LAYER L1M1_PR_C ;
        RECT 120.150 127.750 120.320 127.920 ;
        RECT 118.710 127.010 118.880 127.180 ;
      LAYER mcon ;
        RECT 119.110 126.570 119.280 126.740 ;
        RECT 119.470 126.570 119.640 126.740 ;
        RECT 119.830 126.570 120.000 126.740 ;
        RECT 120.190 126.570 120.360 126.740 ;
        RECT 121.710 126.560 121.880 126.730 ;
        RECT 122.150 126.560 122.320 126.730 ;
        RECT 122.560 126.560 122.730 126.730 ;
        RECT 122.990 126.560 123.160 126.730 ;
        RECT 123.430 126.560 123.600 126.730 ;
        RECT 123.840 126.560 124.010 126.730 ;
        RECT 125.550 126.560 125.720 126.730 ;
        RECT 125.990 126.560 126.160 126.730 ;
        RECT 126.400 126.560 126.570 126.730 ;
        RECT 126.830 126.560 127.000 126.730 ;
        RECT 127.270 126.560 127.440 126.730 ;
        RECT 127.680 126.560 127.850 126.730 ;
        RECT 129.390 126.560 129.560 126.730 ;
        RECT 129.830 126.560 130.000 126.730 ;
        RECT 130.240 126.560 130.410 126.730 ;
        RECT 130.670 126.560 130.840 126.730 ;
        RECT 131.110 126.560 131.280 126.730 ;
        RECT 131.520 126.560 131.690 126.730 ;
        RECT 133.230 126.560 133.400 126.730 ;
        RECT 133.670 126.560 133.840 126.730 ;
        RECT 134.080 126.560 134.250 126.730 ;
        RECT 134.510 126.560 134.680 126.730 ;
        RECT 134.950 126.560 135.120 126.730 ;
        RECT 135.360 126.560 135.530 126.730 ;
        RECT 137.070 126.560 137.240 126.730 ;
        RECT 137.510 126.560 137.680 126.730 ;
        RECT 137.920 126.560 138.090 126.730 ;
        RECT 138.350 126.560 138.520 126.730 ;
        RECT 138.790 126.560 138.960 126.730 ;
        RECT 139.200 126.560 139.370 126.730 ;
        RECT 140.380 126.570 140.550 126.740 ;
        RECT 140.820 126.570 140.990 126.740 ;
        RECT 141.260 126.570 141.430 126.740 ;
        RECT 141.670 126.570 141.840 126.740 ;
      LAYER L1M1_PR_C ;
        RECT 11.670 124.420 11.840 124.590 ;
        RECT 23.190 122.940 23.360 123.110 ;
        RECT 29.910 124.420 30.080 124.590 ;
        RECT 38.070 124.790 38.240 124.960 ;
        RECT 44.310 125.160 44.480 125.330 ;
        RECT 41.430 122.940 41.600 123.110 ;
        RECT 58.230 125.160 58.400 125.330 ;
        RECT 46.230 124.050 46.400 124.220 ;
        RECT 47.670 124.420 47.840 124.590 ;
        RECT 77.430 125.160 77.600 125.330 ;
        RECT 59.670 122.940 59.840 123.110 ;
        RECT 75.030 124.050 75.200 124.220 ;
        RECT 75.990 124.050 76.160 124.220 ;
        RECT 76.950 124.050 77.120 124.220 ;
        RECT 90.870 124.420 91.040 124.590 ;
        RECT 94.230 125.160 94.400 125.330 ;
        RECT 91.830 123.680 92.000 123.850 ;
        RECT 96.630 124.050 96.800 124.220 ;
        RECT 98.070 124.420 98.240 124.590 ;
        RECT 97.110 124.050 97.280 124.220 ;
        RECT 101.430 124.420 101.600 124.590 ;
        RECT 102.390 124.420 102.560 124.590 ;
        RECT 103.830 124.050 104.000 124.220 ;
        RECT 104.790 124.050 104.960 124.220 ;
        RECT 102.870 123.310 103.040 123.480 ;
        RECT 107.190 124.420 107.360 124.590 ;
        RECT 111.990 124.790 112.160 124.960 ;
        RECT 108.150 122.940 108.320 123.110 ;
        RECT 114.870 124.420 115.040 124.590 ;
        RECT 126.390 124.790 126.560 124.960 ;
        RECT 20.310 121.090 20.480 121.260 ;
        RECT 12.150 120.350 12.320 120.520 ;
      LAYER mcon ;
        RECT 6.510 118.420 6.680 118.590 ;
        RECT 6.950 118.420 7.120 118.590 ;
        RECT 7.360 118.420 7.530 118.590 ;
        RECT 7.790 118.420 7.960 118.590 ;
        RECT 8.230 118.420 8.400 118.590 ;
        RECT 8.640 118.420 8.810 118.590 ;
        RECT 11.160 118.430 11.330 118.600 ;
        RECT 11.520 118.430 11.690 118.600 ;
        RECT 13.230 118.420 13.400 118.590 ;
        RECT 13.670 118.420 13.840 118.590 ;
        RECT 14.080 118.420 14.250 118.590 ;
        RECT 14.510 118.420 14.680 118.590 ;
        RECT 14.950 118.420 15.120 118.590 ;
        RECT 15.360 118.420 15.530 118.590 ;
        RECT 17.070 118.420 17.240 118.590 ;
        RECT 17.510 118.420 17.680 118.590 ;
        RECT 17.920 118.420 18.090 118.590 ;
        RECT 18.350 118.420 18.520 118.590 ;
        RECT 18.790 118.420 18.960 118.590 ;
        RECT 19.200 118.420 19.370 118.590 ;
      LAYER L1M1_PR_C ;
        RECT 22.230 119.980 22.400 120.150 ;
        RECT 28.950 121.090 29.120 121.260 ;
      LAYER mcon ;
        RECT 20.760 118.430 20.930 118.600 ;
        RECT 21.120 118.430 21.290 118.600 ;
        RECT 21.480 118.430 21.650 118.600 ;
        RECT 21.840 118.430 22.010 118.600 ;
        RECT 22.200 118.430 22.370 118.600 ;
      LAYER L1M1_PR_C ;
        RECT 24.630 119.610 24.800 119.780 ;
        RECT 25.110 119.610 25.280 119.780 ;
      LAYER mcon ;
        RECT 24.010 118.430 24.180 118.600 ;
        RECT 24.370 118.430 24.540 118.600 ;
        RECT 24.730 118.430 24.900 118.600 ;
        RECT 25.090 118.430 25.260 118.600 ;
        RECT 25.660 118.430 25.830 118.600 ;
        RECT 26.100 118.430 26.270 118.600 ;
        RECT 26.540 118.430 26.710 118.600 ;
        RECT 26.950 118.430 27.120 118.600 ;
      LAYER L1M1_PR_C ;
        RECT 30.870 119.980 31.040 120.150 ;
        RECT 36.150 121.090 36.320 121.260 ;
      LAYER mcon ;
        RECT 29.400 118.430 29.570 118.600 ;
        RECT 29.760 118.430 29.930 118.600 ;
        RECT 30.120 118.430 30.290 118.600 ;
        RECT 30.480 118.430 30.650 118.600 ;
        RECT 30.840 118.430 31.010 118.600 ;
      LAYER L1M1_PR_C ;
        RECT 33.270 119.610 33.440 119.780 ;
        RECT 33.750 119.610 33.920 119.780 ;
        RECT 37.590 120.350 37.760 120.520 ;
      LAYER mcon ;
        RECT 32.650 118.430 32.820 118.600 ;
        RECT 33.010 118.430 33.180 118.600 ;
        RECT 33.370 118.430 33.540 118.600 ;
        RECT 33.730 118.430 33.900 118.600 ;
        RECT 34.300 118.430 34.470 118.600 ;
        RECT 34.740 118.430 34.910 118.600 ;
        RECT 35.180 118.430 35.350 118.600 ;
        RECT 35.590 118.430 35.760 118.600 ;
      LAYER L1M1_PR_C ;
        RECT 43.830 121.090 44.000 121.260 ;
        RECT 45.270 120.720 45.440 120.890 ;
      LAYER mcon ;
        RECT 36.550 118.430 36.720 118.600 ;
        RECT 36.910 118.430 37.080 118.600 ;
        RECT 37.270 118.430 37.440 118.600 ;
        RECT 37.630 118.430 37.800 118.600 ;
        RECT 39.150 118.420 39.320 118.590 ;
        RECT 39.590 118.420 39.760 118.590 ;
        RECT 40.000 118.420 40.170 118.590 ;
        RECT 40.430 118.420 40.600 118.590 ;
        RECT 40.870 118.420 41.040 118.590 ;
        RECT 41.280 118.420 41.450 118.590 ;
        RECT 44.230 118.430 44.400 118.600 ;
        RECT 44.590 118.430 44.760 118.600 ;
        RECT 44.950 118.430 45.120 118.600 ;
        RECT 45.310 118.430 45.480 118.600 ;
        RECT 46.830 118.420 47.000 118.590 ;
        RECT 47.270 118.420 47.440 118.590 ;
        RECT 47.680 118.420 47.850 118.590 ;
        RECT 48.110 118.420 48.280 118.590 ;
        RECT 48.550 118.420 48.720 118.590 ;
        RECT 48.960 118.420 49.130 118.590 ;
        RECT 51.000 118.430 51.170 118.600 ;
        RECT 51.360 118.430 51.530 118.600 ;
      LAYER L1M1_PR_C ;
        RECT 52.950 119.610 53.120 119.780 ;
      LAYER mcon ;
        RECT 52.870 118.430 53.040 118.600 ;
        RECT 53.230 118.430 53.400 118.600 ;
        RECT 55.290 118.430 55.460 118.600 ;
        RECT 55.650 118.430 55.820 118.600 ;
        RECT 56.010 118.430 56.180 118.600 ;
      LAYER L1M1_PR_C ;
        RECT 60.630 118.870 60.800 119.040 ;
      LAYER mcon ;
        RECT 57.230 118.430 57.400 118.600 ;
        RECT 57.590 118.430 57.760 118.600 ;
        RECT 57.950 118.430 58.120 118.600 ;
        RECT 61.770 118.430 61.940 118.600 ;
        RECT 62.130 118.430 62.300 118.600 ;
      LAYER L1M1_PR_C ;
        RECT 68.790 120.350 68.960 120.520 ;
      LAYER mcon ;
        RECT 63.690 118.430 63.860 118.600 ;
        RECT 64.050 118.430 64.220 118.600 ;
        RECT 64.410 118.430 64.580 118.600 ;
        RECT 65.500 118.430 65.670 118.600 ;
        RECT 65.940 118.430 66.110 118.600 ;
        RECT 66.380 118.430 66.550 118.600 ;
        RECT 66.790 118.430 66.960 118.600 ;
        RECT 67.800 118.430 67.970 118.600 ;
        RECT 68.160 118.430 68.330 118.600 ;
      LAYER L1M1_PR_C ;
        RECT 75.510 120.720 75.680 120.890 ;
      LAYER mcon ;
        RECT 69.870 118.420 70.040 118.590 ;
        RECT 70.310 118.420 70.480 118.590 ;
        RECT 70.720 118.420 70.890 118.590 ;
        RECT 71.150 118.420 71.320 118.590 ;
        RECT 71.590 118.420 71.760 118.590 ;
        RECT 72.000 118.420 72.170 118.590 ;
      LAYER L1M1_PR_C ;
        RECT 74.070 118.870 74.240 119.040 ;
      LAYER mcon ;
        RECT 74.470 118.430 74.640 118.600 ;
        RECT 74.830 118.430 75.000 118.600 ;
        RECT 75.190 118.430 75.360 118.600 ;
        RECT 75.550 118.430 75.720 118.600 ;
      LAYER L1M1_PR_C ;
        RECT 78.390 119.980 78.560 120.150 ;
        RECT 79.830 119.980 80.000 120.150 ;
        RECT 80.310 119.610 80.480 119.780 ;
      LAYER mcon ;
        RECT 76.540 118.430 76.710 118.600 ;
        RECT 76.980 118.430 77.150 118.600 ;
        RECT 77.420 118.430 77.590 118.600 ;
        RECT 77.830 118.430 78.000 118.600 ;
        RECT 78.350 118.430 78.520 118.600 ;
        RECT 78.710 118.430 78.880 118.600 ;
        RECT 79.070 118.430 79.240 118.600 ;
      LAYER L1M1_PR_C ;
        RECT 83.190 119.610 83.360 119.780 ;
      LAYER mcon ;
        RECT 79.990 118.430 80.160 118.600 ;
        RECT 80.350 118.430 80.520 118.600 ;
        RECT 80.860 118.430 81.030 118.600 ;
        RECT 81.300 118.430 81.470 118.600 ;
        RECT 81.740 118.430 81.910 118.600 ;
        RECT 82.150 118.430 82.320 118.600 ;
        RECT 82.680 118.430 82.850 118.600 ;
        RECT 83.040 118.430 83.210 118.600 ;
      LAYER L1M1_PR_C ;
        RECT 83.670 118.870 83.840 119.040 ;
        RECT 86.550 119.610 86.720 119.780 ;
      LAYER mcon ;
        RECT 84.220 118.430 84.390 118.600 ;
        RECT 84.660 118.430 84.830 118.600 ;
        RECT 85.100 118.430 85.270 118.600 ;
        RECT 85.510 118.430 85.680 118.600 ;
        RECT 86.040 118.430 86.210 118.600 ;
        RECT 86.400 118.430 86.570 118.600 ;
        RECT 86.760 118.430 86.930 118.600 ;
        RECT 87.120 118.430 87.290 118.600 ;
      LAYER L1M1_PR_C ;
        RECT 90.390 119.980 90.560 120.150 ;
        RECT 91.830 119.980 92.000 120.150 ;
        RECT 92.310 119.610 92.480 119.780 ;
        RECT 87.990 118.870 88.160 119.040 ;
      LAYER mcon ;
        RECT 88.540 118.430 88.710 118.600 ;
        RECT 88.980 118.430 89.150 118.600 ;
        RECT 89.420 118.430 89.590 118.600 ;
        RECT 89.830 118.430 90.000 118.600 ;
        RECT 90.350 118.430 90.520 118.600 ;
        RECT 90.710 118.430 90.880 118.600 ;
        RECT 91.070 118.430 91.240 118.600 ;
      LAYER L1M1_PR_C ;
        RECT 95.670 121.090 95.840 121.260 ;
        RECT 95.190 119.610 95.360 119.780 ;
      LAYER mcon ;
        RECT 91.990 118.430 92.160 118.600 ;
        RECT 92.350 118.430 92.520 118.600 ;
        RECT 92.860 118.430 93.030 118.600 ;
        RECT 93.300 118.430 93.470 118.600 ;
        RECT 93.740 118.430 93.910 118.600 ;
        RECT 94.150 118.430 94.320 118.600 ;
      LAYER L1M1_PR_C ;
        RECT 96.150 119.610 96.320 119.780 ;
        RECT 96.630 119.610 96.800 119.780 ;
        RECT 97.590 119.610 97.760 119.780 ;
      LAYER mcon ;
        RECT 94.680 118.430 94.850 118.600 ;
        RECT 95.040 118.430 95.210 118.600 ;
      LAYER L1M1_PR_C ;
        RECT 101.910 120.720 102.080 120.890 ;
        RECT 101.430 119.610 101.600 119.780 ;
      LAYER mcon ;
        RECT 96.700 118.430 96.870 118.600 ;
        RECT 97.060 118.430 97.230 118.600 ;
        RECT 97.420 118.430 97.590 118.600 ;
        RECT 97.780 118.430 97.950 118.600 ;
        RECT 98.140 118.430 98.310 118.600 ;
        RECT 98.620 118.430 98.790 118.600 ;
        RECT 99.060 118.430 99.230 118.600 ;
        RECT 99.500 118.430 99.670 118.600 ;
        RECT 99.910 118.430 100.080 118.600 ;
        RECT 100.920 118.430 101.090 118.600 ;
        RECT 101.280 118.430 101.450 118.600 ;
      LAYER L1M1_PR_C ;
        RECT 105.750 121.090 105.920 121.260 ;
        RECT 106.710 119.980 106.880 120.150 ;
        RECT 104.310 119.610 104.480 119.780 ;
        RECT 107.190 119.980 107.360 120.150 ;
        RECT 105.270 119.610 105.440 119.780 ;
      LAYER mcon ;
        RECT 102.460 118.430 102.630 118.600 ;
        RECT 102.900 118.430 103.070 118.600 ;
        RECT 103.340 118.430 103.510 118.600 ;
        RECT 103.750 118.430 103.920 118.600 ;
        RECT 106.360 118.430 106.530 118.600 ;
        RECT 106.720 118.430 106.890 118.600 ;
        RECT 107.080 118.430 107.250 118.600 ;
        RECT 108.750 118.420 108.920 118.590 ;
        RECT 109.190 118.420 109.360 118.590 ;
        RECT 109.600 118.420 109.770 118.590 ;
        RECT 110.030 118.420 110.200 118.590 ;
        RECT 110.470 118.420 110.640 118.590 ;
        RECT 110.880 118.420 111.050 118.590 ;
        RECT 112.590 118.420 112.760 118.590 ;
        RECT 113.030 118.420 113.200 118.590 ;
        RECT 113.440 118.420 113.610 118.590 ;
        RECT 113.870 118.420 114.040 118.590 ;
        RECT 114.310 118.420 114.480 118.590 ;
        RECT 114.720 118.420 114.890 118.590 ;
        RECT 116.430 118.420 116.600 118.590 ;
        RECT 116.870 118.420 117.040 118.590 ;
        RECT 117.280 118.420 117.450 118.590 ;
        RECT 117.710 118.420 117.880 118.590 ;
        RECT 118.150 118.420 118.320 118.590 ;
        RECT 118.560 118.420 118.730 118.590 ;
        RECT 120.270 118.420 120.440 118.590 ;
        RECT 120.710 118.420 120.880 118.590 ;
        RECT 121.120 118.420 121.290 118.590 ;
        RECT 121.550 118.420 121.720 118.590 ;
        RECT 121.990 118.420 122.160 118.590 ;
        RECT 122.400 118.420 122.570 118.590 ;
        RECT 124.110 118.420 124.280 118.590 ;
        RECT 124.550 118.420 124.720 118.590 ;
        RECT 124.960 118.420 125.130 118.590 ;
        RECT 125.390 118.420 125.560 118.590 ;
        RECT 125.830 118.420 126.000 118.590 ;
        RECT 126.240 118.420 126.410 118.590 ;
        RECT 127.950 118.420 128.120 118.590 ;
        RECT 128.390 118.420 128.560 118.590 ;
        RECT 128.800 118.420 128.970 118.590 ;
        RECT 129.230 118.420 129.400 118.590 ;
        RECT 129.670 118.420 129.840 118.590 ;
        RECT 130.080 118.420 130.250 118.590 ;
        RECT 131.790 118.420 131.960 118.590 ;
        RECT 132.230 118.420 132.400 118.590 ;
        RECT 132.640 118.420 132.810 118.590 ;
        RECT 133.070 118.420 133.240 118.590 ;
        RECT 133.510 118.420 133.680 118.590 ;
        RECT 133.920 118.420 134.090 118.590 ;
        RECT 135.630 118.420 135.800 118.590 ;
        RECT 136.070 118.420 136.240 118.590 ;
        RECT 136.480 118.420 136.650 118.590 ;
        RECT 136.910 118.420 137.080 118.590 ;
        RECT 137.350 118.420 137.520 118.590 ;
        RECT 137.760 118.420 137.930 118.590 ;
        RECT 138.940 118.430 139.110 118.600 ;
        RECT 139.380 118.430 139.550 118.600 ;
        RECT 139.820 118.430 139.990 118.600 ;
        RECT 140.230 118.430 140.400 118.600 ;
      LAYER L1M1_PR_C ;
        RECT 15.510 116.280 15.680 116.450 ;
        RECT 14.070 114.800 14.240 114.970 ;
        RECT 25.110 116.280 25.280 116.450 ;
        RECT 26.070 116.280 26.240 116.450 ;
        RECT 42.870 116.280 43.040 116.450 ;
        RECT 43.830 116.280 44.000 116.450 ;
        RECT 45.270 115.910 45.440 116.080 ;
        RECT 46.230 115.910 46.400 116.080 ;
        RECT 50.070 116.650 50.240 116.820 ;
        RECT 44.310 115.170 44.480 115.340 ;
        RECT 52.470 115.910 52.640 116.080 ;
        RECT 57.750 115.910 57.920 116.080 ;
        RECT 56.310 115.540 56.480 115.710 ;
        RECT 60.630 117.020 60.800 117.190 ;
        RECT 62.070 115.910 62.240 116.080 ;
        RECT 66.870 115.170 67.040 115.340 ;
        RECT 68.310 115.170 68.480 115.340 ;
        RECT 71.670 116.650 71.840 116.820 ;
        RECT 74.550 116.280 74.720 116.450 ;
        RECT 74.070 115.540 74.240 115.710 ;
        RECT 86.070 117.020 86.240 117.190 ;
        RECT 90.390 116.280 90.560 116.450 ;
        RECT 88.950 114.800 89.120 114.970 ;
        RECT 93.270 117.020 93.440 117.190 ;
        RECT 95.670 115.910 95.840 116.080 ;
        RECT 96.630 116.280 96.800 116.450 ;
        RECT 96.150 115.910 96.320 116.080 ;
        RECT 101.910 116.280 102.080 116.450 ;
        RECT 100.470 115.910 100.640 116.080 ;
        RECT 104.790 116.280 104.960 116.450 ;
        RECT 108.630 115.910 108.800 116.080 ;
        RECT 112.950 116.280 113.120 116.450 ;
        RECT 111.510 114.800 111.680 114.970 ;
        RECT 117.270 114.800 117.440 114.970 ;
        RECT 122.070 116.280 122.240 116.450 ;
        RECT 118.710 114.800 118.880 114.970 ;
        RECT 122.550 114.800 122.720 114.970 ;
        RECT 8.790 112.210 8.960 112.380 ;
      LAYER mcon ;
        RECT 6.350 110.290 6.520 110.460 ;
        RECT 6.710 110.290 6.880 110.460 ;
        RECT 7.070 110.290 7.240 110.460 ;
        RECT 7.990 110.290 8.160 110.460 ;
        RECT 8.350 110.290 8.520 110.460 ;
      LAYER L1M1_PR_C ;
        RECT 9.270 111.100 9.440 111.270 ;
      LAYER mcon ;
        RECT 12.950 110.290 13.120 110.460 ;
        RECT 13.310 110.290 13.480 110.460 ;
        RECT 13.670 110.290 13.840 110.460 ;
      LAYER L1M1_PR_C ;
        RECT 20.790 112.950 20.960 113.120 ;
      LAYER mcon ;
        RECT 16.920 110.290 17.090 110.460 ;
        RECT 17.280 110.290 17.450 110.460 ;
        RECT 17.640 110.290 17.810 110.460 ;
      LAYER L1M1_PR_C ;
        RECT 27.030 111.840 27.200 112.010 ;
        RECT 24.630 111.470 24.800 111.640 ;
        RECT 27.990 111.840 28.160 112.010 ;
        RECT 25.590 111.470 25.760 111.640 ;
      LAYER mcon ;
        RECT 19.530 110.290 19.700 110.460 ;
        RECT 19.890 110.290 20.060 110.460 ;
        RECT 20.250 110.290 20.420 110.460 ;
        RECT 21.340 110.290 21.510 110.460 ;
        RECT 21.780 110.290 21.950 110.460 ;
        RECT 22.220 110.290 22.390 110.460 ;
        RECT 22.630 110.290 22.800 110.460 ;
      LAYER L1M1_PR_C ;
        RECT 25.590 110.730 25.760 110.900 ;
      LAYER mcon ;
        RECT 26.680 110.290 26.850 110.460 ;
        RECT 27.040 110.290 27.210 110.460 ;
        RECT 27.400 110.290 27.570 110.460 ;
        RECT 29.070 110.280 29.240 110.450 ;
        RECT 29.510 110.280 29.680 110.450 ;
        RECT 29.920 110.280 30.090 110.450 ;
        RECT 30.350 110.280 30.520 110.450 ;
        RECT 30.790 110.280 30.960 110.450 ;
        RECT 31.200 110.280 31.370 110.450 ;
        RECT 32.910 110.280 33.080 110.450 ;
        RECT 33.350 110.280 33.520 110.450 ;
        RECT 33.760 110.280 33.930 110.450 ;
        RECT 34.190 110.280 34.360 110.450 ;
        RECT 34.630 110.280 34.800 110.450 ;
        RECT 35.040 110.280 35.210 110.450 ;
      LAYER L1M1_PR_C ;
        RECT 39.030 111.470 39.200 111.640 ;
        RECT 37.590 110.730 37.760 110.900 ;
      LAYER mcon ;
        RECT 37.990 110.290 38.160 110.460 ;
        RECT 38.350 110.290 38.520 110.460 ;
        RECT 38.710 110.290 38.880 110.460 ;
        RECT 39.070 110.290 39.240 110.460 ;
      LAYER L1M1_PR_C ;
        RECT 45.750 111.840 45.920 112.010 ;
      LAYER mcon ;
        RECT 40.060 110.290 40.230 110.460 ;
        RECT 40.500 110.290 40.670 110.460 ;
        RECT 40.940 110.290 41.110 110.460 ;
        RECT 41.350 110.290 41.520 110.460 ;
        RECT 41.880 110.290 42.050 110.460 ;
        RECT 42.240 110.290 42.410 110.460 ;
        RECT 42.600 110.290 42.770 110.460 ;
      LAYER L1M1_PR_C ;
        RECT 44.310 111.100 44.480 111.270 ;
      LAYER mcon ;
        RECT 43.440 110.290 43.610 110.460 ;
        RECT 43.800 110.290 43.970 110.460 ;
        RECT 44.160 110.290 44.330 110.460 ;
        RECT 45.000 110.290 45.170 110.460 ;
        RECT 45.360 110.290 45.530 110.460 ;
        RECT 45.720 110.290 45.890 110.460 ;
      LAYER L1M1_PR_C ;
        RECT 52.470 111.840 52.640 112.010 ;
      LAYER mcon ;
        RECT 46.780 110.290 46.950 110.460 ;
        RECT 47.220 110.290 47.390 110.460 ;
        RECT 47.660 110.290 47.830 110.460 ;
        RECT 48.070 110.290 48.240 110.460 ;
        RECT 48.600 110.290 48.770 110.460 ;
        RECT 48.960 110.290 49.130 110.460 ;
        RECT 49.320 110.290 49.490 110.460 ;
      LAYER L1M1_PR_C ;
        RECT 51.030 111.100 51.200 111.270 ;
      LAYER mcon ;
        RECT 50.160 110.290 50.330 110.460 ;
        RECT 50.520 110.290 50.690 110.460 ;
        RECT 50.880 110.290 51.050 110.460 ;
        RECT 51.720 110.290 51.890 110.460 ;
        RECT 52.080 110.290 52.250 110.460 ;
        RECT 52.440 110.290 52.610 110.460 ;
      LAYER L1M1_PR_C ;
        RECT 59.190 111.840 59.360 112.010 ;
        RECT 55.350 111.470 55.520 111.640 ;
      LAYER mcon ;
        RECT 53.500 110.290 53.670 110.460 ;
        RECT 53.940 110.290 54.110 110.460 ;
        RECT 54.380 110.290 54.550 110.460 ;
        RECT 54.790 110.290 54.960 110.460 ;
        RECT 55.320 110.290 55.490 110.460 ;
        RECT 55.680 110.290 55.850 110.460 ;
        RECT 56.040 110.290 56.210 110.460 ;
        RECT 56.880 110.290 57.050 110.460 ;
        RECT 57.240 110.290 57.410 110.460 ;
        RECT 57.600 110.290 57.770 110.460 ;
        RECT 58.440 110.290 58.610 110.460 ;
        RECT 58.800 110.290 58.970 110.460 ;
        RECT 59.160 110.290 59.330 110.460 ;
      LAYER L1M1_PR_C ;
        RECT 66.870 111.840 67.040 112.010 ;
        RECT 72.150 112.950 72.320 113.120 ;
      LAYER mcon ;
        RECT 60.220 110.290 60.390 110.460 ;
        RECT 60.660 110.290 60.830 110.460 ;
        RECT 61.100 110.290 61.270 110.460 ;
        RECT 61.510 110.290 61.680 110.460 ;
        RECT 63.000 110.290 63.170 110.460 ;
        RECT 63.360 110.290 63.530 110.460 ;
        RECT 63.720 110.290 63.890 110.460 ;
      LAYER L1M1_PR_C ;
        RECT 65.430 111.100 65.600 111.270 ;
      LAYER mcon ;
        RECT 64.560 110.290 64.730 110.460 ;
        RECT 64.920 110.290 65.090 110.460 ;
        RECT 65.280 110.290 65.450 110.460 ;
        RECT 66.120 110.290 66.290 110.460 ;
        RECT 66.480 110.290 66.650 110.460 ;
        RECT 66.840 110.290 67.010 110.460 ;
        RECT 68.430 110.280 68.600 110.450 ;
        RECT 68.870 110.280 69.040 110.450 ;
        RECT 69.280 110.280 69.450 110.450 ;
        RECT 69.710 110.280 69.880 110.450 ;
        RECT 70.150 110.280 70.320 110.450 ;
        RECT 70.560 110.280 70.730 110.450 ;
      LAYER L1M1_PR_C ;
        RECT 73.590 111.470 73.760 111.640 ;
      LAYER mcon ;
        RECT 72.550 110.290 72.720 110.460 ;
        RECT 72.910 110.290 73.080 110.460 ;
        RECT 73.270 110.290 73.440 110.460 ;
        RECT 73.630 110.290 73.800 110.460 ;
      LAYER L1M1_PR_C ;
        RECT 82.710 112.950 82.880 113.120 ;
        RECT 78.870 111.470 79.040 111.640 ;
        RECT 79.830 111.840 80.000 112.010 ;
      LAYER mcon ;
        RECT 74.620 110.290 74.790 110.460 ;
        RECT 75.060 110.290 75.230 110.460 ;
        RECT 75.500 110.290 75.670 110.460 ;
        RECT 75.910 110.290 76.080 110.460 ;
        RECT 77.920 110.290 78.090 110.460 ;
        RECT 78.280 110.290 78.450 110.460 ;
        RECT 78.640 110.290 78.810 110.460 ;
      LAYER L1M1_PR_C ;
        RECT 79.830 110.730 80.000 110.900 ;
      LAYER mcon ;
        RECT 80.860 110.290 81.030 110.460 ;
        RECT 81.300 110.290 81.470 110.460 ;
        RECT 81.740 110.290 81.910 110.460 ;
        RECT 82.150 110.290 82.320 110.460 ;
      LAYER L1M1_PR_C ;
        RECT 89.910 112.950 90.080 113.120 ;
        RECT 85.110 111.840 85.280 112.010 ;
        RECT 85.590 111.470 85.760 111.640 ;
        RECT 86.550 111.470 86.720 111.640 ;
        RECT 91.830 111.470 92.000 111.640 ;
        RECT 93.750 111.470 93.920 111.640 ;
      LAYER mcon ;
        RECT 83.120 110.290 83.290 110.460 ;
        RECT 83.480 110.290 83.650 110.460 ;
        RECT 83.840 110.290 84.010 110.460 ;
        RECT 86.480 110.290 86.650 110.460 ;
        RECT 86.840 110.290 87.010 110.460 ;
        RECT 87.200 110.290 87.370 110.460 ;
        RECT 87.560 110.290 87.730 110.460 ;
        RECT 88.060 110.290 88.230 110.460 ;
        RECT 88.500 110.290 88.670 110.460 ;
        RECT 88.940 110.290 89.110 110.460 ;
        RECT 89.350 110.290 89.520 110.460 ;
        RECT 90.400 110.290 90.570 110.460 ;
        RECT 90.760 110.290 90.930 110.460 ;
        RECT 91.120 110.290 91.290 110.460 ;
        RECT 91.480 110.290 91.650 110.460 ;
        RECT 91.840 110.290 92.010 110.460 ;
      LAYER L1M1_PR_C ;
        RECT 99.990 111.840 100.160 112.010 ;
        RECT 96.150 111.470 96.320 111.640 ;
      LAYER mcon ;
        RECT 92.650 110.290 92.820 110.460 ;
        RECT 93.010 110.290 93.180 110.460 ;
        RECT 93.370 110.290 93.540 110.460 ;
        RECT 93.730 110.290 93.900 110.460 ;
        RECT 94.300 110.290 94.470 110.460 ;
        RECT 94.740 110.290 94.910 110.460 ;
        RECT 95.180 110.290 95.350 110.460 ;
        RECT 95.590 110.290 95.760 110.460 ;
        RECT 96.120 110.290 96.290 110.460 ;
        RECT 96.480 110.290 96.650 110.460 ;
        RECT 96.840 110.290 97.010 110.460 ;
        RECT 97.680 110.290 97.850 110.460 ;
        RECT 98.040 110.290 98.210 110.460 ;
        RECT 98.400 110.290 98.570 110.460 ;
        RECT 99.240 110.290 99.410 110.460 ;
        RECT 99.600 110.290 99.770 110.460 ;
        RECT 99.960 110.290 100.130 110.460 ;
      LAYER L1M1_PR_C ;
        RECT 106.710 111.840 106.880 112.010 ;
        RECT 102.870 111.470 103.040 111.640 ;
      LAYER mcon ;
        RECT 101.020 110.290 101.190 110.460 ;
        RECT 101.460 110.290 101.630 110.460 ;
        RECT 101.900 110.290 102.070 110.460 ;
        RECT 102.310 110.290 102.480 110.460 ;
        RECT 102.840 110.290 103.010 110.460 ;
        RECT 103.200 110.290 103.370 110.460 ;
        RECT 103.560 110.290 103.730 110.460 ;
        RECT 104.400 110.290 104.570 110.460 ;
        RECT 104.760 110.290 104.930 110.460 ;
        RECT 105.120 110.290 105.290 110.460 ;
        RECT 105.960 110.290 106.130 110.460 ;
        RECT 106.320 110.290 106.490 110.460 ;
        RECT 106.680 110.290 106.850 110.460 ;
        RECT 107.740 110.290 107.910 110.460 ;
        RECT 108.180 110.290 108.350 110.460 ;
        RECT 108.620 110.290 108.790 110.460 ;
        RECT 109.030 110.290 109.200 110.460 ;
      LAYER L1M1_PR_C ;
        RECT 110.070 111.840 110.240 112.010 ;
      LAYER mcon ;
        RECT 110.030 110.290 110.200 110.460 ;
        RECT 110.390 110.290 110.560 110.460 ;
        RECT 110.750 110.290 110.920 110.460 ;
        RECT 111.670 110.290 111.840 110.460 ;
        RECT 112.030 110.290 112.200 110.460 ;
      LAYER L1M1_PR_C ;
        RECT 112.950 111.470 113.120 111.640 ;
      LAYER mcon ;
        RECT 116.630 110.290 116.800 110.460 ;
        RECT 116.990 110.290 117.160 110.460 ;
        RECT 117.350 110.290 117.520 110.460 ;
      LAYER L1M1_PR_C ;
        RECT 121.110 111.100 121.280 111.270 ;
        RECT 124.470 112.950 124.640 113.120 ;
      LAYER mcon ;
        RECT 120.600 110.290 120.770 110.460 ;
        RECT 120.960 110.290 121.130 110.460 ;
        RECT 121.320 110.290 121.490 110.460 ;
        RECT 123.210 110.290 123.380 110.460 ;
        RECT 123.570 110.290 123.740 110.460 ;
        RECT 123.930 110.290 124.100 110.460 ;
        RECT 125.550 110.280 125.720 110.450 ;
        RECT 125.990 110.280 126.160 110.450 ;
        RECT 126.400 110.280 126.570 110.450 ;
        RECT 126.830 110.280 127.000 110.450 ;
        RECT 127.270 110.280 127.440 110.450 ;
        RECT 127.680 110.280 127.850 110.450 ;
        RECT 129.390 110.280 129.560 110.450 ;
        RECT 129.830 110.280 130.000 110.450 ;
        RECT 130.240 110.280 130.410 110.450 ;
        RECT 130.670 110.280 130.840 110.450 ;
        RECT 131.110 110.280 131.280 110.450 ;
        RECT 131.520 110.280 131.690 110.450 ;
        RECT 133.230 110.280 133.400 110.450 ;
        RECT 133.670 110.280 133.840 110.450 ;
        RECT 134.080 110.280 134.250 110.450 ;
        RECT 134.510 110.280 134.680 110.450 ;
        RECT 134.950 110.280 135.120 110.450 ;
        RECT 135.360 110.280 135.530 110.450 ;
        RECT 137.070 110.280 137.240 110.450 ;
        RECT 137.510 110.280 137.680 110.450 ;
        RECT 137.920 110.280 138.090 110.450 ;
        RECT 138.350 110.280 138.520 110.450 ;
        RECT 138.790 110.280 138.960 110.450 ;
        RECT 139.200 110.280 139.370 110.450 ;
        RECT 140.380 110.290 140.550 110.460 ;
        RECT 140.820 110.290 140.990 110.460 ;
        RECT 141.260 110.290 141.430 110.460 ;
        RECT 141.670 110.290 141.840 110.460 ;
      LAYER L1M1_PR_C ;
        RECT 23.190 108.140 23.360 108.310 ;
        RECT 24.150 108.140 24.320 108.310 ;
        RECT 25.590 107.770 25.760 107.940 ;
        RECT 26.550 107.770 26.720 107.940 ;
        RECT 24.630 106.660 24.800 106.830 ;
        RECT 31.830 108.140 32.000 108.310 ;
        RECT 32.310 108.140 32.480 108.310 ;
        RECT 47.190 106.660 47.360 106.830 ;
        RECT 52.950 108.880 53.120 109.050 ;
        RECT 61.110 108.510 61.280 108.680 ;
        RECT 69.270 108.510 69.440 108.680 ;
        RECT 70.710 107.770 70.880 107.940 ;
        RECT 75.990 108.140 76.160 108.310 ;
        RECT 74.070 107.770 74.240 107.940 ;
        RECT 75.510 107.770 75.680 107.940 ;
        RECT 78.390 108.140 78.560 108.310 ;
        RECT 79.350 108.140 79.520 108.310 ;
        RECT 80.790 107.770 80.960 107.940 ;
        RECT 81.750 107.770 81.920 107.940 ;
        RECT 79.830 106.660 80.000 106.830 ;
        RECT 87.030 108.140 87.200 108.310 ;
        RECT 86.550 107.770 86.720 107.940 ;
        RECT 87.990 108.140 88.160 108.310 ;
        RECT 84.150 107.030 84.320 107.200 ;
        RECT 92.310 108.140 92.480 108.310 ;
        RECT 96.150 107.770 96.320 107.940 ;
        RECT 99.030 108.140 99.200 108.310 ;
        RECT 102.870 107.770 103.040 107.940 ;
        RECT 107.670 108.510 107.840 108.680 ;
        RECT 109.590 107.770 109.760 107.940 ;
        RECT 112.470 108.880 112.640 109.050 ;
        RECT 113.910 108.140 114.080 108.310 ;
        RECT 117.270 108.880 117.440 109.050 ;
        RECT 123.990 108.510 124.160 108.680 ;
        RECT 118.710 106.660 118.880 106.830 ;
        RECT 125.430 107.770 125.600 107.940 ;
      LAYER mcon ;
        RECT 6.510 102.140 6.680 102.310 ;
        RECT 6.950 102.140 7.120 102.310 ;
        RECT 7.360 102.140 7.530 102.310 ;
        RECT 7.790 102.140 7.960 102.310 ;
        RECT 8.230 102.140 8.400 102.310 ;
        RECT 8.640 102.140 8.810 102.310 ;
        RECT 10.190 102.150 10.360 102.320 ;
        RECT 10.550 102.150 10.720 102.320 ;
        RECT 10.910 102.150 11.080 102.320 ;
        RECT 11.830 102.150 12.000 102.320 ;
        RECT 12.190 102.150 12.360 102.320 ;
      LAYER L1M1_PR_C ;
        RECT 13.110 103.330 13.280 103.500 ;
      LAYER mcon ;
        RECT 16.790 102.150 16.960 102.320 ;
        RECT 17.150 102.150 17.320 102.320 ;
        RECT 17.510 102.150 17.680 102.320 ;
      LAYER L1M1_PR_C ;
        RECT 21.270 102.960 21.440 103.130 ;
        RECT 24.630 103.330 24.800 103.500 ;
      LAYER mcon ;
        RECT 20.760 102.150 20.930 102.320 ;
        RECT 21.120 102.150 21.290 102.320 ;
        RECT 21.480 102.150 21.650 102.320 ;
      LAYER L1M1_PR_C ;
        RECT 27.990 104.810 28.160 104.980 ;
        RECT 31.350 104.810 31.520 104.980 ;
        RECT 27.510 103.330 27.680 103.500 ;
      LAYER mcon ;
        RECT 23.370 102.150 23.540 102.320 ;
        RECT 23.730 102.150 23.900 102.320 ;
        RECT 24.090 102.150 24.260 102.320 ;
        RECT 25.180 102.150 25.350 102.320 ;
        RECT 25.620 102.150 25.790 102.320 ;
        RECT 26.060 102.150 26.230 102.320 ;
        RECT 26.470 102.150 26.640 102.320 ;
        RECT 27.000 102.150 27.170 102.320 ;
        RECT 27.360 102.150 27.530 102.320 ;
        RECT 28.540 102.150 28.710 102.320 ;
        RECT 28.980 102.150 29.150 102.320 ;
        RECT 29.420 102.150 29.590 102.320 ;
        RECT 29.830 102.150 30.000 102.320 ;
      LAYER L1M1_PR_C ;
        RECT 33.270 104.810 33.440 104.980 ;
      LAYER mcon ;
        RECT 31.800 102.150 31.970 102.320 ;
        RECT 32.160 102.150 32.330 102.320 ;
        RECT 32.520 102.150 32.690 102.320 ;
        RECT 32.880 102.150 33.050 102.320 ;
        RECT 33.240 102.150 33.410 102.320 ;
      LAYER L1M1_PR_C ;
        RECT 36.150 103.330 36.320 103.500 ;
        RECT 44.790 103.700 44.960 103.870 ;
        RECT 40.950 103.330 41.120 103.500 ;
      LAYER mcon ;
        RECT 35.050 102.150 35.220 102.320 ;
        RECT 35.410 102.150 35.580 102.320 ;
        RECT 35.770 102.150 35.940 102.320 ;
        RECT 36.130 102.150 36.300 102.320 ;
        RECT 37.230 102.140 37.400 102.310 ;
        RECT 37.670 102.140 37.840 102.310 ;
        RECT 38.080 102.140 38.250 102.310 ;
        RECT 38.510 102.140 38.680 102.310 ;
        RECT 38.950 102.140 39.120 102.310 ;
        RECT 39.360 102.140 39.530 102.310 ;
        RECT 40.920 102.150 41.090 102.320 ;
        RECT 41.280 102.150 41.450 102.320 ;
        RECT 41.640 102.150 41.810 102.320 ;
        RECT 42.480 102.150 42.650 102.320 ;
        RECT 42.840 102.150 43.010 102.320 ;
        RECT 43.200 102.150 43.370 102.320 ;
        RECT 44.040 102.150 44.210 102.320 ;
        RECT 44.400 102.150 44.570 102.320 ;
        RECT 44.760 102.150 44.930 102.320 ;
      LAYER L1M1_PR_C ;
        RECT 51.510 103.700 51.680 103.870 ;
      LAYER mcon ;
        RECT 45.820 102.150 45.990 102.320 ;
        RECT 46.260 102.150 46.430 102.320 ;
        RECT 46.700 102.150 46.870 102.320 ;
        RECT 47.110 102.150 47.280 102.320 ;
        RECT 47.640 102.150 47.810 102.320 ;
        RECT 48.000 102.150 48.170 102.320 ;
        RECT 48.360 102.150 48.530 102.320 ;
      LAYER L1M1_PR_C ;
        RECT 50.070 102.960 50.240 103.130 ;
      LAYER mcon ;
        RECT 49.200 102.150 49.370 102.320 ;
        RECT 49.560 102.150 49.730 102.320 ;
        RECT 49.920 102.150 50.090 102.320 ;
        RECT 50.760 102.150 50.930 102.320 ;
        RECT 51.120 102.150 51.290 102.320 ;
        RECT 51.480 102.150 51.650 102.320 ;
      LAYER L1M1_PR_C ;
        RECT 58.230 103.700 58.400 103.870 ;
        RECT 54.390 103.330 54.560 103.500 ;
      LAYER mcon ;
        RECT 52.540 102.150 52.710 102.320 ;
        RECT 52.980 102.150 53.150 102.320 ;
        RECT 53.420 102.150 53.590 102.320 ;
        RECT 53.830 102.150 54.000 102.320 ;
        RECT 54.360 102.150 54.530 102.320 ;
        RECT 54.720 102.150 54.890 102.320 ;
        RECT 55.080 102.150 55.250 102.320 ;
        RECT 55.920 102.150 56.090 102.320 ;
        RECT 56.280 102.150 56.450 102.320 ;
        RECT 56.640 102.150 56.810 102.320 ;
        RECT 57.480 102.150 57.650 102.320 ;
        RECT 57.840 102.150 58.010 102.320 ;
        RECT 58.200 102.150 58.370 102.320 ;
      LAYER L1M1_PR_C ;
        RECT 62.550 104.810 62.720 104.980 ;
      LAYER mcon ;
        RECT 59.260 102.150 59.430 102.320 ;
        RECT 59.700 102.150 59.870 102.320 ;
        RECT 60.140 102.150 60.310 102.320 ;
        RECT 60.550 102.150 60.720 102.320 ;
        RECT 61.560 102.150 61.730 102.320 ;
        RECT 61.920 102.150 62.090 102.320 ;
        RECT 63.100 102.150 63.270 102.320 ;
        RECT 63.540 102.150 63.710 102.320 ;
        RECT 63.980 102.150 64.150 102.320 ;
        RECT 64.390 102.150 64.560 102.320 ;
      LAYER L1M1_PR_C ;
        RECT 65.430 102.960 65.600 103.130 ;
      LAYER mcon ;
        RECT 65.390 102.150 65.560 102.320 ;
        RECT 65.750 102.150 65.920 102.320 ;
        RECT 66.110 102.150 66.280 102.320 ;
        RECT 67.030 102.150 67.200 102.320 ;
        RECT 67.390 102.150 67.560 102.320 ;
      LAYER L1M1_PR_C ;
        RECT 68.310 103.330 68.480 103.500 ;
      LAYER mcon ;
        RECT 71.990 102.150 72.160 102.320 ;
        RECT 72.350 102.150 72.520 102.320 ;
        RECT 72.710 102.150 72.880 102.320 ;
      LAYER L1M1_PR_C ;
        RECT 76.470 102.960 76.640 103.130 ;
        RECT 79.830 104.810 80.000 104.980 ;
      LAYER mcon ;
        RECT 75.960 102.150 76.130 102.320 ;
        RECT 76.320 102.150 76.490 102.320 ;
        RECT 76.680 102.150 76.850 102.320 ;
      LAYER L1M1_PR_C ;
        RECT 86.070 103.700 86.240 103.870 ;
        RECT 82.230 103.330 82.400 103.500 ;
      LAYER mcon ;
        RECT 78.570 102.150 78.740 102.320 ;
        RECT 78.930 102.150 79.100 102.320 ;
        RECT 79.290 102.150 79.460 102.320 ;
        RECT 80.380 102.150 80.550 102.320 ;
        RECT 80.820 102.150 80.990 102.320 ;
        RECT 81.260 102.150 81.430 102.320 ;
        RECT 81.670 102.150 81.840 102.320 ;
        RECT 82.200 102.150 82.370 102.320 ;
        RECT 82.560 102.150 82.730 102.320 ;
        RECT 82.920 102.150 83.090 102.320 ;
        RECT 83.760 102.150 83.930 102.320 ;
        RECT 84.120 102.150 84.290 102.320 ;
        RECT 84.480 102.150 84.650 102.320 ;
        RECT 85.320 102.150 85.490 102.320 ;
        RECT 85.680 102.150 85.850 102.320 ;
        RECT 86.040 102.150 86.210 102.320 ;
      LAYER L1M1_PR_C ;
        RECT 92.790 103.700 92.960 103.870 ;
        RECT 88.950 103.330 89.120 103.500 ;
        RECT 98.550 104.810 98.720 104.980 ;
      LAYER mcon ;
        RECT 87.100 102.150 87.270 102.320 ;
        RECT 87.540 102.150 87.710 102.320 ;
        RECT 87.980 102.150 88.150 102.320 ;
        RECT 88.390 102.150 88.560 102.320 ;
        RECT 88.920 102.150 89.090 102.320 ;
        RECT 89.280 102.150 89.450 102.320 ;
        RECT 89.640 102.150 89.810 102.320 ;
        RECT 90.480 102.150 90.650 102.320 ;
        RECT 90.840 102.150 91.010 102.320 ;
        RECT 91.200 102.150 91.370 102.320 ;
        RECT 92.040 102.150 92.210 102.320 ;
        RECT 92.400 102.150 92.570 102.320 ;
        RECT 92.760 102.150 92.930 102.320 ;
        RECT 94.350 102.140 94.520 102.310 ;
        RECT 94.790 102.140 94.960 102.310 ;
        RECT 95.200 102.140 95.370 102.310 ;
        RECT 95.630 102.140 95.800 102.310 ;
        RECT 96.070 102.140 96.240 102.310 ;
        RECT 96.480 102.140 96.650 102.310 ;
      LAYER L1M1_PR_C ;
        RECT 99.990 103.700 100.160 103.870 ;
        RECT 101.430 103.330 101.600 103.500 ;
        RECT 102.390 103.330 102.560 103.500 ;
        RECT 109.590 103.700 109.760 103.870 ;
        RECT 105.750 103.330 105.920 103.500 ;
      LAYER mcon ;
        RECT 98.960 102.150 99.130 102.320 ;
        RECT 99.320 102.150 99.490 102.320 ;
        RECT 99.680 102.150 99.850 102.320 ;
        RECT 102.320 102.150 102.490 102.320 ;
        RECT 102.680 102.150 102.850 102.320 ;
        RECT 103.040 102.150 103.210 102.320 ;
        RECT 103.400 102.150 103.570 102.320 ;
        RECT 103.900 102.150 104.070 102.320 ;
        RECT 104.340 102.150 104.510 102.320 ;
        RECT 104.780 102.150 104.950 102.320 ;
        RECT 105.190 102.150 105.360 102.320 ;
        RECT 105.720 102.150 105.890 102.320 ;
        RECT 106.080 102.150 106.250 102.320 ;
        RECT 106.440 102.150 106.610 102.320 ;
        RECT 107.280 102.150 107.450 102.320 ;
        RECT 107.640 102.150 107.810 102.320 ;
        RECT 108.000 102.150 108.170 102.320 ;
        RECT 108.840 102.150 109.010 102.320 ;
        RECT 109.200 102.150 109.370 102.320 ;
        RECT 109.560 102.150 109.730 102.320 ;
      LAYER L1M1_PR_C ;
        RECT 116.310 103.700 116.480 103.870 ;
        RECT 112.470 103.330 112.640 103.500 ;
      LAYER mcon ;
        RECT 110.620 102.150 110.790 102.320 ;
        RECT 111.060 102.150 111.230 102.320 ;
        RECT 111.500 102.150 111.670 102.320 ;
        RECT 111.910 102.150 112.080 102.320 ;
        RECT 112.440 102.150 112.610 102.320 ;
        RECT 112.800 102.150 112.970 102.320 ;
        RECT 113.160 102.150 113.330 102.320 ;
        RECT 114.000 102.150 114.170 102.320 ;
        RECT 114.360 102.150 114.530 102.320 ;
        RECT 114.720 102.150 114.890 102.320 ;
        RECT 115.560 102.150 115.730 102.320 ;
        RECT 115.920 102.150 116.090 102.320 ;
        RECT 116.280 102.150 116.450 102.320 ;
      LAYER L1M1_PR_C ;
        RECT 125.430 103.700 125.600 103.870 ;
      LAYER mcon ;
        RECT 117.870 102.140 118.040 102.310 ;
        RECT 118.310 102.140 118.480 102.310 ;
        RECT 118.720 102.140 118.890 102.310 ;
        RECT 119.150 102.140 119.320 102.310 ;
        RECT 119.590 102.140 119.760 102.310 ;
        RECT 120.000 102.140 120.170 102.310 ;
        RECT 121.560 102.150 121.730 102.320 ;
        RECT 121.920 102.150 122.090 102.320 ;
        RECT 122.280 102.150 122.450 102.320 ;
      LAYER L1M1_PR_C ;
        RECT 123.990 102.960 124.160 103.130 ;
      LAYER mcon ;
        RECT 123.120 102.150 123.290 102.320 ;
        RECT 123.480 102.150 123.650 102.320 ;
        RECT 123.840 102.150 124.010 102.320 ;
        RECT 124.680 102.150 124.850 102.320 ;
        RECT 125.040 102.150 125.210 102.320 ;
        RECT 125.400 102.150 125.570 102.320 ;
      LAYER L1M1_PR_C ;
        RECT 135.990 104.070 136.160 104.240 ;
      LAYER mcon ;
        RECT 126.990 102.140 127.160 102.310 ;
        RECT 127.430 102.140 127.600 102.310 ;
        RECT 127.840 102.140 128.010 102.310 ;
        RECT 128.270 102.140 128.440 102.310 ;
        RECT 128.710 102.140 128.880 102.310 ;
        RECT 129.120 102.140 129.290 102.310 ;
        RECT 130.830 102.140 131.000 102.310 ;
        RECT 131.270 102.140 131.440 102.310 ;
        RECT 131.680 102.140 131.850 102.310 ;
        RECT 132.110 102.140 132.280 102.310 ;
        RECT 132.550 102.140 132.720 102.310 ;
        RECT 132.960 102.140 133.130 102.310 ;
        RECT 135.000 102.150 135.170 102.320 ;
        RECT 135.360 102.150 135.530 102.320 ;
        RECT 137.070 102.140 137.240 102.310 ;
        RECT 137.510 102.140 137.680 102.310 ;
        RECT 137.920 102.140 138.090 102.310 ;
        RECT 138.350 102.140 138.520 102.310 ;
        RECT 138.790 102.140 138.960 102.310 ;
        RECT 139.200 102.140 139.370 102.310 ;
        RECT 140.380 102.150 140.550 102.320 ;
        RECT 140.820 102.150 140.990 102.320 ;
        RECT 141.260 102.150 141.430 102.320 ;
        RECT 141.670 102.150 141.840 102.320 ;
      LAYER L1M1_PR_C ;
        RECT 16.470 100.740 16.640 100.910 ;
        RECT 22.230 100.000 22.400 100.170 ;
        RECT 17.910 98.520 18.080 98.690 ;
        RECT 29.430 100.000 29.600 100.170 ;
        RECT 32.310 100.370 32.480 100.540 ;
        RECT 23.190 98.520 23.360 98.690 ;
        RECT 33.750 100.000 33.920 100.170 ;
        RECT 29.910 98.520 30.080 98.690 ;
        RECT 36.630 98.520 36.800 98.690 ;
        RECT 38.070 98.890 38.240 99.060 ;
        RECT 43.350 100.370 43.520 100.540 ;
        RECT 44.790 99.630 44.960 99.800 ;
        RECT 50.070 100.370 50.240 100.540 ;
        RECT 51.510 99.630 51.680 99.800 ;
        RECT 54.390 100.000 54.560 100.170 ;
        RECT 58.230 99.630 58.400 99.800 ;
        RECT 61.110 100.000 61.280 100.170 ;
        RECT 62.070 100.000 62.240 100.170 ;
        RECT 66.870 100.740 67.040 100.910 ;
        RECT 62.550 99.630 62.720 99.800 ;
        RECT 63.510 99.630 63.680 99.800 ;
        RECT 64.470 99.630 64.640 99.800 ;
        RECT 75.030 100.370 75.200 100.540 ;
        RECT 72.630 99.630 72.800 99.800 ;
        RECT 74.070 99.630 74.240 99.800 ;
        RECT 74.550 99.630 74.720 99.800 ;
        RECT 68.310 98.520 68.480 98.690 ;
        RECT 78.870 100.000 79.040 100.170 ;
        RECT 81.750 99.630 81.920 99.800 ;
        RECT 84.630 100.000 84.800 100.170 ;
        RECT 88.470 99.630 88.640 99.800 ;
        RECT 93.270 100.000 93.440 100.170 ;
        RECT 97.110 99.630 97.280 99.800 ;
        RECT 99.990 100.370 100.160 100.540 ;
        RECT 102.870 100.000 103.040 100.170 ;
        RECT 103.350 100.000 103.520 100.170 ;
        RECT 108.630 100.000 108.800 100.170 ;
        RECT 107.190 98.890 107.360 99.060 ;
        RECT 111.990 99.260 112.160 99.430 ;
        RECT 113.910 100.000 114.080 100.170 ;
        RECT 118.710 100.000 118.880 100.170 ;
        RECT 128.310 100.000 128.480 100.170 ;
        RECT 132.150 99.630 132.320 99.800 ;
      LAYER mcon ;
        RECT 6.350 94.010 6.520 94.180 ;
        RECT 6.710 94.010 6.880 94.180 ;
        RECT 7.070 94.010 7.240 94.180 ;
        RECT 7.990 94.010 8.160 94.180 ;
        RECT 8.350 94.010 8.520 94.180 ;
      LAYER L1M1_PR_C ;
        RECT 9.270 94.450 9.440 94.620 ;
      LAYER mcon ;
        RECT 12.950 94.010 13.120 94.180 ;
        RECT 13.310 94.010 13.480 94.180 ;
        RECT 13.670 94.010 13.840 94.180 ;
      LAYER L1M1_PR_C ;
        RECT 20.790 96.670 20.960 96.840 ;
      LAYER mcon ;
        RECT 16.920 94.010 17.090 94.180 ;
        RECT 17.280 94.010 17.450 94.180 ;
        RECT 17.640 94.010 17.810 94.180 ;
      LAYER L1M1_PR_C ;
        RECT 27.510 95.560 27.680 95.730 ;
        RECT 25.110 95.190 25.280 95.360 ;
        RECT 27.990 95.560 28.160 95.730 ;
        RECT 26.070 95.190 26.240 95.360 ;
      LAYER mcon ;
        RECT 19.530 94.010 19.700 94.180 ;
        RECT 19.890 94.010 20.060 94.180 ;
        RECT 20.250 94.010 20.420 94.180 ;
        RECT 21.870 94.000 22.040 94.170 ;
        RECT 22.310 94.000 22.480 94.170 ;
        RECT 22.720 94.000 22.890 94.170 ;
        RECT 23.150 94.000 23.320 94.170 ;
        RECT 23.590 94.000 23.760 94.170 ;
        RECT 24.000 94.000 24.170 94.170 ;
      LAYER L1M1_PR_C ;
        RECT 26.070 94.450 26.240 94.620 ;
      LAYER mcon ;
        RECT 27.160 94.010 27.330 94.180 ;
        RECT 27.520 94.010 27.690 94.180 ;
        RECT 27.880 94.010 28.050 94.180 ;
      LAYER L1M1_PR_C ;
        RECT 34.710 96.670 34.880 96.840 ;
      LAYER mcon ;
        RECT 29.550 94.000 29.720 94.170 ;
        RECT 29.990 94.000 30.160 94.170 ;
        RECT 30.400 94.000 30.570 94.170 ;
        RECT 30.830 94.000 31.000 94.170 ;
        RECT 31.270 94.000 31.440 94.170 ;
        RECT 31.680 94.000 31.850 94.170 ;
      LAYER L1M1_PR_C ;
        RECT 37.590 96.670 37.760 96.840 ;
        RECT 33.270 94.450 33.440 94.620 ;
      LAYER mcon ;
        RECT 33.670 94.010 33.840 94.180 ;
        RECT 34.030 94.010 34.200 94.180 ;
        RECT 34.390 94.010 34.560 94.180 ;
        RECT 34.750 94.010 34.920 94.180 ;
      LAYER L1M1_PR_C ;
        RECT 39.030 96.300 39.200 96.470 ;
      LAYER mcon ;
        RECT 35.740 94.010 35.910 94.180 ;
        RECT 36.180 94.010 36.350 94.180 ;
        RECT 36.620 94.010 36.790 94.180 ;
        RECT 37.030 94.010 37.200 94.180 ;
        RECT 37.990 94.010 38.160 94.180 ;
        RECT 38.350 94.010 38.520 94.180 ;
        RECT 38.710 94.010 38.880 94.180 ;
        RECT 39.070 94.010 39.240 94.180 ;
      LAYER L1M1_PR_C ;
        RECT 45.750 95.560 45.920 95.730 ;
        RECT 41.910 95.190 42.080 95.360 ;
      LAYER mcon ;
        RECT 40.060 94.010 40.230 94.180 ;
        RECT 40.500 94.010 40.670 94.180 ;
        RECT 40.940 94.010 41.110 94.180 ;
        RECT 41.350 94.010 41.520 94.180 ;
        RECT 41.880 94.010 42.050 94.180 ;
        RECT 42.240 94.010 42.410 94.180 ;
        RECT 42.600 94.010 42.770 94.180 ;
        RECT 43.440 94.010 43.610 94.180 ;
        RECT 43.800 94.010 43.970 94.180 ;
        RECT 44.160 94.010 44.330 94.180 ;
        RECT 45.000 94.010 45.170 94.180 ;
        RECT 45.360 94.010 45.530 94.180 ;
        RECT 45.720 94.010 45.890 94.180 ;
      LAYER L1M1_PR_C ;
        RECT 52.470 95.560 52.640 95.730 ;
      LAYER mcon ;
        RECT 46.780 94.010 46.950 94.180 ;
        RECT 47.220 94.010 47.390 94.180 ;
        RECT 47.660 94.010 47.830 94.180 ;
        RECT 48.070 94.010 48.240 94.180 ;
        RECT 48.600 94.010 48.770 94.180 ;
        RECT 48.960 94.010 49.130 94.180 ;
        RECT 49.320 94.010 49.490 94.180 ;
      LAYER L1M1_PR_C ;
        RECT 51.030 94.820 51.200 94.990 ;
      LAYER mcon ;
        RECT 50.160 94.010 50.330 94.180 ;
        RECT 50.520 94.010 50.690 94.180 ;
        RECT 50.880 94.010 51.050 94.180 ;
        RECT 51.720 94.010 51.890 94.180 ;
        RECT 52.080 94.010 52.250 94.180 ;
        RECT 52.440 94.010 52.610 94.180 ;
      LAYER L1M1_PR_C ;
        RECT 59.190 95.560 59.360 95.730 ;
        RECT 55.350 95.190 55.520 95.360 ;
      LAYER mcon ;
        RECT 53.500 94.010 53.670 94.180 ;
        RECT 53.940 94.010 54.110 94.180 ;
        RECT 54.380 94.010 54.550 94.180 ;
        RECT 54.790 94.010 54.960 94.180 ;
        RECT 55.320 94.010 55.490 94.180 ;
        RECT 55.680 94.010 55.850 94.180 ;
        RECT 56.040 94.010 56.210 94.180 ;
        RECT 56.880 94.010 57.050 94.180 ;
        RECT 57.240 94.010 57.410 94.180 ;
        RECT 57.600 94.010 57.770 94.180 ;
        RECT 58.440 94.010 58.610 94.180 ;
        RECT 58.800 94.010 58.970 94.180 ;
        RECT 59.160 94.010 59.330 94.180 ;
      LAYER L1M1_PR_C ;
        RECT 63.510 96.670 63.680 96.840 ;
      LAYER mcon ;
        RECT 60.220 94.010 60.390 94.180 ;
        RECT 60.660 94.010 60.830 94.180 ;
        RECT 61.100 94.010 61.270 94.180 ;
        RECT 61.510 94.010 61.680 94.180 ;
      LAYER L1M1_PR_C ;
        RECT 62.070 94.450 62.240 94.620 ;
      LAYER mcon ;
        RECT 62.470 94.010 62.640 94.180 ;
        RECT 62.830 94.010 63.000 94.180 ;
        RECT 63.190 94.010 63.360 94.180 ;
        RECT 63.550 94.010 63.720 94.180 ;
      LAYER L1M1_PR_C ;
        RECT 67.350 96.670 67.520 96.840 ;
        RECT 69.750 96.670 69.920 96.840 ;
        RECT 66.870 95.190 67.040 95.360 ;
      LAYER mcon ;
        RECT 64.540 94.010 64.710 94.180 ;
        RECT 64.980 94.010 65.150 94.180 ;
        RECT 65.420 94.010 65.590 94.180 ;
        RECT 65.830 94.010 66.000 94.180 ;
        RECT 66.360 94.010 66.530 94.180 ;
        RECT 66.720 94.010 66.890 94.180 ;
      LAYER L1M1_PR_C ;
        RECT 71.190 96.300 71.360 96.470 ;
      LAYER mcon ;
        RECT 67.900 94.010 68.070 94.180 ;
        RECT 68.340 94.010 68.510 94.180 ;
        RECT 68.780 94.010 68.950 94.180 ;
        RECT 69.190 94.010 69.360 94.180 ;
        RECT 70.150 94.010 70.320 94.180 ;
        RECT 70.510 94.010 70.680 94.180 ;
        RECT 70.870 94.010 71.040 94.180 ;
        RECT 71.230 94.010 71.400 94.180 ;
      LAYER L1M1_PR_C ;
        RECT 74.070 95.930 74.240 96.100 ;
        RECT 75.990 96.300 76.160 96.470 ;
        RECT 75.030 95.190 75.200 95.360 ;
        RECT 75.990 95.190 76.160 95.360 ;
        RECT 77.430 95.560 77.600 95.730 ;
      LAYER mcon ;
        RECT 72.220 94.010 72.390 94.180 ;
        RECT 72.660 94.010 72.830 94.180 ;
        RECT 73.100 94.010 73.270 94.180 ;
        RECT 73.510 94.010 73.680 94.180 ;
        RECT 75.040 94.010 75.210 94.180 ;
        RECT 75.400 94.010 75.570 94.180 ;
        RECT 75.760 94.010 75.930 94.180 ;
      LAYER L1M1_PR_C ;
        RECT 83.670 95.560 83.840 95.730 ;
      LAYER mcon ;
        RECT 77.980 94.010 78.150 94.180 ;
        RECT 78.420 94.010 78.590 94.180 ;
        RECT 78.860 94.010 79.030 94.180 ;
        RECT 79.270 94.010 79.440 94.180 ;
        RECT 79.800 94.010 79.970 94.180 ;
        RECT 80.160 94.010 80.330 94.180 ;
        RECT 80.520 94.010 80.690 94.180 ;
      LAYER L1M1_PR_C ;
        RECT 81.270 94.820 81.440 94.990 ;
      LAYER mcon ;
        RECT 81.360 94.010 81.530 94.180 ;
        RECT 81.720 94.010 81.890 94.180 ;
        RECT 82.080 94.010 82.250 94.180 ;
        RECT 82.920 94.010 83.090 94.180 ;
        RECT 83.280 94.010 83.450 94.180 ;
        RECT 83.640 94.010 83.810 94.180 ;
      LAYER L1M1_PR_C ;
        RECT 90.390 95.560 90.560 95.730 ;
      LAYER mcon ;
        RECT 84.700 94.010 84.870 94.180 ;
        RECT 85.140 94.010 85.310 94.180 ;
        RECT 85.580 94.010 85.750 94.180 ;
        RECT 85.990 94.010 86.160 94.180 ;
        RECT 86.520 94.010 86.690 94.180 ;
        RECT 86.880 94.010 87.050 94.180 ;
        RECT 87.240 94.010 87.410 94.180 ;
      LAYER L1M1_PR_C ;
        RECT 87.990 94.820 88.160 94.990 ;
      LAYER mcon ;
        RECT 88.080 94.010 88.250 94.180 ;
        RECT 88.440 94.010 88.610 94.180 ;
        RECT 88.800 94.010 88.970 94.180 ;
        RECT 89.640 94.010 89.810 94.180 ;
        RECT 90.000 94.010 90.170 94.180 ;
        RECT 90.360 94.010 90.530 94.180 ;
      LAYER L1M1_PR_C ;
        RECT 93.270 95.560 93.440 95.730 ;
        RECT 93.750 95.560 93.920 95.730 ;
        RECT 95.190 95.560 95.360 95.730 ;
        RECT 95.670 96.670 95.840 96.840 ;
      LAYER mcon ;
        RECT 91.420 94.010 91.590 94.180 ;
        RECT 91.860 94.010 92.030 94.180 ;
        RECT 92.300 94.010 92.470 94.180 ;
        RECT 92.710 94.010 92.880 94.180 ;
        RECT 93.240 94.010 93.410 94.180 ;
        RECT 93.600 94.010 93.770 94.180 ;
        RECT 94.510 94.010 94.680 94.180 ;
        RECT 94.870 94.010 95.040 94.180 ;
        RECT 95.230 94.010 95.400 94.180 ;
      LAYER L1M1_PR_C ;
        RECT 102.870 95.560 103.040 95.730 ;
      LAYER mcon ;
        RECT 96.700 94.010 96.870 94.180 ;
        RECT 97.140 94.010 97.310 94.180 ;
        RECT 97.580 94.010 97.750 94.180 ;
        RECT 97.990 94.010 98.160 94.180 ;
        RECT 99.000 94.010 99.170 94.180 ;
        RECT 99.360 94.010 99.530 94.180 ;
        RECT 99.720 94.010 99.890 94.180 ;
      LAYER L1M1_PR_C ;
        RECT 100.950 94.820 101.120 94.990 ;
      LAYER mcon ;
        RECT 100.560 94.010 100.730 94.180 ;
        RECT 100.920 94.010 101.090 94.180 ;
        RECT 101.280 94.010 101.450 94.180 ;
        RECT 102.120 94.010 102.290 94.180 ;
        RECT 102.480 94.010 102.650 94.180 ;
        RECT 102.840 94.010 103.010 94.180 ;
      LAYER L1M1_PR_C ;
        RECT 109.590 95.560 109.760 95.730 ;
      LAYER mcon ;
        RECT 103.900 94.010 104.070 94.180 ;
        RECT 104.340 94.010 104.510 94.180 ;
        RECT 104.780 94.010 104.950 94.180 ;
        RECT 105.190 94.010 105.360 94.180 ;
        RECT 105.720 94.010 105.890 94.180 ;
        RECT 106.080 94.010 106.250 94.180 ;
        RECT 106.440 94.010 106.610 94.180 ;
      LAYER L1M1_PR_C ;
        RECT 108.150 94.820 108.320 94.990 ;
      LAYER mcon ;
        RECT 107.280 94.010 107.450 94.180 ;
        RECT 107.640 94.010 107.810 94.180 ;
        RECT 108.000 94.010 108.170 94.180 ;
        RECT 108.840 94.010 109.010 94.180 ;
        RECT 109.200 94.010 109.370 94.180 ;
        RECT 109.560 94.010 109.730 94.180 ;
      LAYER L1M1_PR_C ;
        RECT 114.390 96.670 114.560 96.840 ;
        RECT 112.470 95.560 112.640 95.730 ;
        RECT 113.910 95.560 114.080 95.730 ;
        RECT 116.790 96.670 116.960 96.840 ;
      LAYER mcon ;
        RECT 110.620 94.010 110.790 94.180 ;
        RECT 111.060 94.010 111.230 94.180 ;
        RECT 111.500 94.010 111.670 94.180 ;
        RECT 111.910 94.010 112.080 94.180 ;
        RECT 112.430 94.010 112.600 94.180 ;
        RECT 112.790 94.010 112.960 94.180 ;
        RECT 113.150 94.010 113.320 94.180 ;
      LAYER L1M1_PR_C ;
        RECT 118.230 96.670 118.400 96.840 ;
      LAYER mcon ;
        RECT 114.070 94.010 114.240 94.180 ;
        RECT 114.430 94.010 114.600 94.180 ;
        RECT 114.940 94.010 115.110 94.180 ;
        RECT 115.380 94.010 115.550 94.180 ;
        RECT 115.820 94.010 115.990 94.180 ;
        RECT 116.230 94.010 116.400 94.180 ;
        RECT 117.190 94.010 117.360 94.180 ;
        RECT 117.550 94.010 117.720 94.180 ;
        RECT 117.910 94.010 118.080 94.180 ;
        RECT 118.270 94.010 118.440 94.180 ;
      LAYER L1M1_PR_C ;
        RECT 125.430 95.560 125.600 95.730 ;
      LAYER mcon ;
        RECT 119.260 94.010 119.430 94.180 ;
        RECT 119.700 94.010 119.870 94.180 ;
        RECT 120.140 94.010 120.310 94.180 ;
        RECT 120.550 94.010 120.720 94.180 ;
        RECT 121.560 94.010 121.730 94.180 ;
        RECT 121.920 94.010 122.090 94.180 ;
        RECT 122.280 94.010 122.450 94.180 ;
      LAYER L1M1_PR_C ;
        RECT 123.990 94.820 124.160 94.990 ;
      LAYER mcon ;
        RECT 123.120 94.010 123.290 94.180 ;
        RECT 123.480 94.010 123.650 94.180 ;
        RECT 123.840 94.010 124.010 94.180 ;
        RECT 124.680 94.010 124.850 94.180 ;
        RECT 125.040 94.010 125.210 94.180 ;
        RECT 125.400 94.010 125.570 94.180 ;
        RECT 126.460 94.010 126.630 94.180 ;
        RECT 126.900 94.010 127.070 94.180 ;
        RECT 127.340 94.010 127.510 94.180 ;
        RECT 127.750 94.010 127.920 94.180 ;
        RECT 128.710 94.010 128.880 94.180 ;
        RECT 129.070 94.010 129.240 94.180 ;
        RECT 129.430 94.010 129.600 94.180 ;
        RECT 129.790 94.010 129.960 94.180 ;
        RECT 131.310 94.000 131.480 94.170 ;
        RECT 131.750 94.000 131.920 94.170 ;
        RECT 132.160 94.000 132.330 94.170 ;
        RECT 132.590 94.000 132.760 94.170 ;
        RECT 133.030 94.000 133.200 94.170 ;
        RECT 133.440 94.000 133.610 94.170 ;
        RECT 135.150 94.000 135.320 94.170 ;
        RECT 135.590 94.000 135.760 94.170 ;
        RECT 136.000 94.000 136.170 94.170 ;
        RECT 136.430 94.000 136.600 94.170 ;
        RECT 136.870 94.000 137.040 94.170 ;
        RECT 137.280 94.000 137.450 94.170 ;
        RECT 138.990 94.000 139.160 94.170 ;
        RECT 139.430 94.000 139.600 94.170 ;
        RECT 139.840 94.000 140.010 94.170 ;
        RECT 140.270 94.000 140.440 94.170 ;
        RECT 140.710 94.000 140.880 94.170 ;
        RECT 141.120 94.000 141.290 94.170 ;
      LAYER L1M1_PR_C ;
        RECT 13.110 92.600 13.280 92.770 ;
        RECT 25.110 92.230 25.280 92.400 ;
        RECT 24.150 91.860 24.320 92.030 ;
        RECT 28.470 92.600 28.640 92.770 ;
        RECT 14.550 90.380 14.720 90.550 ;
        RECT 27.510 91.860 27.680 92.030 ;
        RECT 28.470 91.860 28.640 92.030 ;
        RECT 29.910 91.490 30.080 91.660 ;
        RECT 30.390 91.490 30.560 91.660 ;
        RECT 33.270 90.750 33.440 90.920 ;
        RECT 34.710 90.380 34.880 90.550 ;
        RECT 39.990 91.860 40.160 92.030 ;
        RECT 45.750 92.600 45.920 92.770 ;
        RECT 57.270 92.230 57.440 92.400 ;
        RECT 60.150 91.860 60.320 92.030 ;
        RECT 59.670 91.120 59.840 91.290 ;
        RECT 77.430 92.230 77.600 92.400 ;
        RECT 71.670 90.380 71.840 90.550 ;
        RECT 78.870 91.490 79.040 91.660 ;
        RECT 84.150 92.230 84.320 92.400 ;
        RECT 85.590 91.490 85.760 91.660 ;
        RECT 88.470 91.860 88.640 92.030 ;
        RECT 92.310 91.490 92.480 91.660 ;
        RECT 97.110 92.230 97.280 92.400 ;
        RECT 99.030 91.490 99.200 91.660 ;
        RECT 101.910 91.860 102.080 92.030 ;
        RECT 105.750 91.490 105.920 91.660 ;
        RECT 111.030 92.600 111.200 92.770 ;
        RECT 108.630 91.860 108.800 92.030 ;
        RECT 109.590 91.860 109.760 92.030 ;
        RECT 111.030 91.490 111.200 91.660 ;
        RECT 113.910 91.860 114.080 92.030 ;
        RECT 114.870 91.490 115.040 91.660 ;
        RECT 118.710 91.860 118.880 92.030 ;
        RECT 117.270 90.750 117.440 90.920 ;
        RECT 123.990 92.230 124.160 92.400 ;
        RECT 125.430 91.490 125.600 91.660 ;
      LAYER mcon ;
        RECT 6.510 85.860 6.680 86.030 ;
        RECT 6.950 85.860 7.120 86.030 ;
        RECT 7.360 85.860 7.530 86.030 ;
        RECT 7.790 85.860 7.960 86.030 ;
        RECT 8.230 85.860 8.400 86.030 ;
        RECT 8.640 85.860 8.810 86.030 ;
        RECT 10.350 85.860 10.520 86.030 ;
        RECT 10.790 85.860 10.960 86.030 ;
        RECT 11.200 85.860 11.370 86.030 ;
        RECT 11.630 85.860 11.800 86.030 ;
        RECT 12.070 85.860 12.240 86.030 ;
        RECT 12.480 85.860 12.650 86.030 ;
      LAYER L1M1_PR_C ;
        RECT 21.750 88.160 21.920 88.330 ;
        RECT 21.270 87.050 21.440 87.220 ;
      LAYER mcon ;
        RECT 14.190 85.860 14.360 86.030 ;
        RECT 14.630 85.860 14.800 86.030 ;
        RECT 15.040 85.860 15.210 86.030 ;
        RECT 15.470 85.860 15.640 86.030 ;
        RECT 15.910 85.860 16.080 86.030 ;
        RECT 16.320 85.860 16.490 86.030 ;
        RECT 17.500 85.870 17.670 86.040 ;
        RECT 17.940 85.870 18.110 86.040 ;
        RECT 18.380 85.870 18.550 86.040 ;
        RECT 18.790 85.870 18.960 86.040 ;
        RECT 20.760 85.870 20.930 86.040 ;
        RECT 21.120 85.870 21.290 86.040 ;
      LAYER L1M1_PR_C ;
        RECT 27.510 88.530 27.680 88.700 ;
        RECT 24.630 87.050 24.800 87.220 ;
      LAYER mcon ;
        RECT 22.300 85.870 22.470 86.040 ;
        RECT 22.740 85.870 22.910 86.040 ;
        RECT 23.180 85.870 23.350 86.040 ;
        RECT 23.590 85.870 23.760 86.040 ;
        RECT 24.120 85.870 24.290 86.040 ;
        RECT 24.480 85.870 24.650 86.040 ;
      LAYER L1M1_PR_C ;
        RECT 25.110 86.680 25.280 86.850 ;
        RECT 28.950 87.790 29.120 87.960 ;
      LAYER mcon ;
        RECT 25.660 85.870 25.830 86.040 ;
        RECT 26.100 85.870 26.270 86.040 ;
        RECT 26.540 85.870 26.710 86.040 ;
        RECT 26.950 85.870 27.120 86.040 ;
        RECT 27.910 85.870 28.080 86.040 ;
        RECT 28.270 85.870 28.440 86.040 ;
        RECT 28.630 85.870 28.800 86.040 ;
        RECT 28.990 85.870 29.160 86.040 ;
      LAYER L1M1_PR_C ;
        RECT 35.670 87.420 35.840 87.590 ;
        RECT 31.830 87.050 32.000 87.220 ;
      LAYER mcon ;
        RECT 29.980 85.870 30.150 86.040 ;
        RECT 30.420 85.870 30.590 86.040 ;
        RECT 30.860 85.870 31.030 86.040 ;
        RECT 31.270 85.870 31.440 86.040 ;
        RECT 31.800 85.870 31.970 86.040 ;
        RECT 32.160 85.870 32.330 86.040 ;
        RECT 32.520 85.870 32.690 86.040 ;
        RECT 33.360 85.870 33.530 86.040 ;
        RECT 33.720 85.870 33.890 86.040 ;
        RECT 34.080 85.870 34.250 86.040 ;
        RECT 34.920 85.870 35.090 86.040 ;
        RECT 35.280 85.870 35.450 86.040 ;
        RECT 35.640 85.870 35.810 86.040 ;
      LAYER L1M1_PR_C ;
        RECT 42.390 87.420 42.560 87.590 ;
        RECT 38.550 87.050 38.720 87.220 ;
      LAYER mcon ;
        RECT 36.700 85.870 36.870 86.040 ;
        RECT 37.140 85.870 37.310 86.040 ;
        RECT 37.580 85.870 37.750 86.040 ;
        RECT 37.990 85.870 38.160 86.040 ;
        RECT 38.520 85.870 38.690 86.040 ;
        RECT 38.880 85.870 39.050 86.040 ;
        RECT 39.240 85.870 39.410 86.040 ;
        RECT 40.080 85.870 40.250 86.040 ;
        RECT 40.440 85.870 40.610 86.040 ;
        RECT 40.800 85.870 40.970 86.040 ;
        RECT 41.640 85.870 41.810 86.040 ;
        RECT 42.000 85.870 42.170 86.040 ;
        RECT 42.360 85.870 42.530 86.040 ;
      LAYER L1M1_PR_C ;
        RECT 49.110 87.420 49.280 87.590 ;
      LAYER mcon ;
        RECT 43.420 85.870 43.590 86.040 ;
        RECT 43.860 85.870 44.030 86.040 ;
        RECT 44.300 85.870 44.470 86.040 ;
        RECT 44.710 85.870 44.880 86.040 ;
        RECT 45.240 85.870 45.410 86.040 ;
        RECT 45.600 85.870 45.770 86.040 ;
        RECT 45.960 85.870 46.130 86.040 ;
      LAYER L1M1_PR_C ;
        RECT 46.710 86.680 46.880 86.850 ;
      LAYER mcon ;
        RECT 46.800 85.870 46.970 86.040 ;
        RECT 47.160 85.870 47.330 86.040 ;
        RECT 47.520 85.870 47.690 86.040 ;
        RECT 48.360 85.870 48.530 86.040 ;
        RECT 48.720 85.870 48.890 86.040 ;
        RECT 49.080 85.870 49.250 86.040 ;
      LAYER L1M1_PR_C ;
        RECT 53.430 88.530 53.600 88.700 ;
        RECT 57.750 88.530 57.920 88.700 ;
        RECT 54.390 87.420 54.560 87.590 ;
        RECT 51.990 87.050 52.160 87.220 ;
        RECT 55.350 87.420 55.520 87.590 ;
        RECT 52.950 87.050 53.120 87.220 ;
      LAYER mcon ;
        RECT 50.140 85.870 50.310 86.040 ;
        RECT 50.580 85.870 50.750 86.040 ;
        RECT 51.020 85.870 51.190 86.040 ;
        RECT 51.430 85.870 51.600 86.040 ;
        RECT 54.040 85.870 54.210 86.040 ;
        RECT 54.400 85.870 54.570 86.040 ;
        RECT 54.760 85.870 54.930 86.040 ;
        RECT 55.900 85.870 56.070 86.040 ;
        RECT 56.340 85.870 56.510 86.040 ;
        RECT 56.780 85.870 56.950 86.040 ;
        RECT 57.190 85.870 57.360 86.040 ;
      LAYER L1M1_PR_C ;
        RECT 59.190 87.420 59.360 87.590 ;
        RECT 63.990 88.530 64.160 88.700 ;
        RECT 61.590 87.050 61.760 87.220 ;
      LAYER mcon ;
        RECT 58.200 85.870 58.370 86.040 ;
        RECT 58.710 85.870 58.880 86.040 ;
        RECT 60.390 85.870 60.560 86.040 ;
        RECT 60.750 85.870 60.920 86.040 ;
        RECT 61.110 85.870 61.280 86.040 ;
      LAYER L1M1_PR_C ;
        RECT 65.430 88.530 65.600 88.700 ;
      LAYER mcon ;
        RECT 62.140 85.870 62.310 86.040 ;
        RECT 62.580 85.870 62.750 86.040 ;
        RECT 63.020 85.870 63.190 86.040 ;
        RECT 63.430 85.870 63.600 86.040 ;
        RECT 64.390 85.870 64.560 86.040 ;
        RECT 64.750 85.870 64.920 86.040 ;
        RECT 65.110 85.870 65.280 86.040 ;
        RECT 65.470 85.870 65.640 86.040 ;
      LAYER L1M1_PR_C ;
        RECT 69.750 88.530 69.920 88.700 ;
        RECT 69.270 87.050 69.440 87.220 ;
      LAYER mcon ;
        RECT 66.460 85.870 66.630 86.040 ;
        RECT 66.900 85.870 67.070 86.040 ;
        RECT 67.340 85.870 67.510 86.040 ;
        RECT 67.750 85.870 67.920 86.040 ;
        RECT 68.760 85.870 68.930 86.040 ;
        RECT 69.120 85.870 69.290 86.040 ;
      LAYER L1M1_PR_C ;
        RECT 72.630 87.050 72.800 87.220 ;
      LAYER mcon ;
        RECT 70.300 85.870 70.470 86.040 ;
        RECT 70.740 85.870 70.910 86.040 ;
        RECT 71.180 85.870 71.350 86.040 ;
        RECT 71.590 85.870 71.760 86.040 ;
      LAYER L1M1_PR_C ;
        RECT 74.070 86.680 74.240 86.850 ;
        RECT 74.550 86.680 74.720 86.850 ;
        RECT 75.030 86.310 75.200 86.480 ;
        RECT 81.270 87.420 81.440 87.590 ;
      LAYER mcon ;
        RECT 72.100 85.870 72.270 86.040 ;
        RECT 72.460 85.870 72.630 86.040 ;
        RECT 72.820 85.870 72.990 86.040 ;
        RECT 73.180 85.870 73.350 86.040 ;
        RECT 73.540 85.870 73.710 86.040 ;
        RECT 75.580 85.870 75.750 86.040 ;
        RECT 76.020 85.870 76.190 86.040 ;
        RECT 76.460 85.870 76.630 86.040 ;
        RECT 76.870 85.870 77.040 86.040 ;
        RECT 77.400 85.870 77.570 86.040 ;
        RECT 77.760 85.870 77.930 86.040 ;
        RECT 78.120 85.870 78.290 86.040 ;
      LAYER L1M1_PR_C ;
        RECT 79.830 86.680 80.000 86.850 ;
      LAYER mcon ;
        RECT 78.960 85.870 79.130 86.040 ;
        RECT 79.320 85.870 79.490 86.040 ;
        RECT 79.680 85.870 79.850 86.040 ;
        RECT 80.520 85.870 80.690 86.040 ;
        RECT 80.880 85.870 81.050 86.040 ;
        RECT 81.240 85.870 81.410 86.040 ;
      LAYER L1M1_PR_C ;
        RECT 87.990 87.420 88.160 87.590 ;
        RECT 84.150 87.050 84.320 87.220 ;
      LAYER mcon ;
        RECT 82.300 85.870 82.470 86.040 ;
        RECT 82.740 85.870 82.910 86.040 ;
        RECT 83.180 85.870 83.350 86.040 ;
        RECT 83.590 85.870 83.760 86.040 ;
        RECT 84.120 85.870 84.290 86.040 ;
        RECT 84.480 85.870 84.650 86.040 ;
        RECT 84.840 85.870 85.010 86.040 ;
        RECT 85.680 85.870 85.850 86.040 ;
        RECT 86.040 85.870 86.210 86.040 ;
        RECT 86.400 85.870 86.570 86.040 ;
        RECT 87.240 85.870 87.410 86.040 ;
        RECT 87.600 85.870 87.770 86.040 ;
        RECT 87.960 85.870 88.130 86.040 ;
      LAYER L1M1_PR_C ;
        RECT 97.590 87.420 97.760 87.590 ;
        RECT 93.750 87.050 93.920 87.220 ;
      LAYER mcon ;
        RECT 89.550 85.860 89.720 86.030 ;
        RECT 89.990 85.860 90.160 86.030 ;
        RECT 90.400 85.860 90.570 86.030 ;
        RECT 90.830 85.860 91.000 86.030 ;
        RECT 91.270 85.860 91.440 86.030 ;
        RECT 91.680 85.860 91.850 86.030 ;
        RECT 93.720 85.870 93.890 86.040 ;
        RECT 94.080 85.870 94.250 86.040 ;
        RECT 94.440 85.870 94.610 86.040 ;
        RECT 95.280 85.870 95.450 86.040 ;
        RECT 95.640 85.870 95.810 86.040 ;
        RECT 96.000 85.870 96.170 86.040 ;
        RECT 96.840 85.870 97.010 86.040 ;
        RECT 97.200 85.870 97.370 86.040 ;
        RECT 97.560 85.870 97.730 86.040 ;
      LAYER L1M1_PR_C ;
        RECT 101.910 87.790 102.080 87.960 ;
        RECT 103.350 87.420 103.520 87.590 ;
      LAYER mcon ;
        RECT 98.620 85.870 98.790 86.040 ;
        RECT 99.060 85.870 99.230 86.040 ;
        RECT 99.500 85.870 99.670 86.040 ;
        RECT 99.910 85.870 100.080 86.040 ;
        RECT 102.360 85.870 102.530 86.040 ;
        RECT 102.720 85.870 102.890 86.040 ;
        RECT 103.080 85.870 103.250 86.040 ;
        RECT 103.440 85.870 103.610 86.040 ;
        RECT 103.800 85.870 103.970 86.040 ;
      LAYER L1M1_PR_C ;
        RECT 104.790 86.680 104.960 86.850 ;
      LAYER mcon ;
        RECT 104.850 85.870 105.020 86.040 ;
        RECT 105.210 85.870 105.380 86.040 ;
        RECT 105.570 85.870 105.740 86.040 ;
        RECT 105.930 85.870 106.100 86.040 ;
        RECT 106.290 85.870 106.460 86.040 ;
      LAYER L1M1_PR_C ;
        RECT 111.030 88.530 111.200 88.700 ;
        RECT 109.110 87.420 109.280 87.590 ;
        RECT 110.550 87.420 110.720 87.590 ;
      LAYER mcon ;
        RECT 107.260 85.870 107.430 86.040 ;
        RECT 107.700 85.870 107.870 86.040 ;
        RECT 108.140 85.870 108.310 86.040 ;
        RECT 108.550 85.870 108.720 86.040 ;
        RECT 109.070 85.870 109.240 86.040 ;
        RECT 109.430 85.870 109.600 86.040 ;
        RECT 109.790 85.870 109.960 86.040 ;
      LAYER L1M1_PR_C ;
        RECT 114.870 87.790 115.040 87.960 ;
      LAYER mcon ;
        RECT 110.710 85.870 110.880 86.040 ;
        RECT 111.070 85.870 111.240 86.040 ;
        RECT 111.580 85.870 111.750 86.040 ;
        RECT 112.020 85.870 112.190 86.040 ;
        RECT 112.460 85.870 112.630 86.040 ;
        RECT 112.870 85.870 113.040 86.040 ;
      LAYER L1M1_PR_C ;
        RECT 118.230 88.530 118.400 88.700 ;
        RECT 113.430 86.310 113.600 86.480 ;
      LAYER mcon ;
        RECT 113.830 85.870 114.000 86.040 ;
        RECT 114.190 85.870 114.360 86.040 ;
        RECT 114.550 85.870 114.720 86.040 ;
        RECT 114.910 85.870 115.080 86.040 ;
        RECT 115.900 85.870 116.070 86.040 ;
        RECT 116.340 85.870 116.510 86.040 ;
        RECT 116.780 85.870 116.950 86.040 ;
        RECT 117.190 85.870 117.360 86.040 ;
      LAYER L1M1_PR_C ;
        RECT 119.670 87.050 119.840 87.220 ;
      LAYER mcon ;
        RECT 118.630 85.870 118.800 86.040 ;
        RECT 118.990 85.870 119.160 86.040 ;
        RECT 119.350 85.870 119.520 86.040 ;
        RECT 119.710 85.870 119.880 86.040 ;
        RECT 121.230 85.860 121.400 86.030 ;
        RECT 121.670 85.860 121.840 86.030 ;
        RECT 122.080 85.860 122.250 86.030 ;
        RECT 122.510 85.860 122.680 86.030 ;
        RECT 122.950 85.860 123.120 86.030 ;
        RECT 123.360 85.860 123.530 86.030 ;
        RECT 125.070 85.860 125.240 86.030 ;
        RECT 125.510 85.860 125.680 86.030 ;
        RECT 125.920 85.860 126.090 86.030 ;
        RECT 126.350 85.860 126.520 86.030 ;
        RECT 126.790 85.860 126.960 86.030 ;
        RECT 127.200 85.860 127.370 86.030 ;
        RECT 128.910 85.860 129.080 86.030 ;
        RECT 129.350 85.860 129.520 86.030 ;
        RECT 129.760 85.860 129.930 86.030 ;
        RECT 130.190 85.860 130.360 86.030 ;
        RECT 130.630 85.860 130.800 86.030 ;
        RECT 131.040 85.860 131.210 86.030 ;
        RECT 132.220 85.870 132.390 86.040 ;
        RECT 132.660 85.870 132.830 86.040 ;
        RECT 133.100 85.870 133.270 86.040 ;
        RECT 133.510 85.870 133.680 86.040 ;
        RECT 136.000 85.870 136.170 86.040 ;
        RECT 136.360 85.870 136.530 86.040 ;
        RECT 137.550 85.860 137.720 86.030 ;
        RECT 137.990 85.860 138.160 86.030 ;
        RECT 138.400 85.860 138.570 86.030 ;
        RECT 138.830 85.860 139.000 86.030 ;
        RECT 139.270 85.860 139.440 86.030 ;
        RECT 139.680 85.860 139.850 86.030 ;
      LAYER L1M1_PR_C ;
        RECT 11.190 84.460 11.360 84.630 ;
        RECT 19.350 84.090 19.520 84.260 ;
        RECT 22.710 84.460 22.880 84.630 ;
        RECT 26.550 83.720 26.720 83.890 ;
        RECT 25.110 82.610 25.280 82.780 ;
        RECT 29.430 83.720 29.600 83.890 ;
        RECT 30.390 83.720 30.560 83.890 ;
        RECT 31.830 83.350 32.000 83.520 ;
        RECT 32.790 83.350 32.960 83.520 ;
        RECT 30.870 82.240 31.040 82.410 ;
        RECT 35.190 82.240 35.360 82.410 ;
        RECT 39.510 83.720 39.680 83.890 ;
        RECT 36.630 82.240 36.800 82.410 ;
        RECT 43.350 83.350 43.520 83.520 ;
        RECT 49.110 83.720 49.280 83.890 ;
        RECT 52.950 83.350 53.120 83.520 ;
        RECT 55.830 83.720 56.000 83.890 ;
        RECT 59.670 83.350 59.840 83.520 ;
        RECT 64.950 82.240 65.120 82.410 ;
        RECT 66.390 82.610 66.560 82.780 ;
        RECT 73.590 84.090 73.760 84.260 ;
        RECT 72.630 83.720 72.800 83.890 ;
        RECT 74.070 83.720 74.240 83.890 ;
        RECT 77.430 84.090 77.600 84.260 ;
        RECT 78.390 84.090 78.560 84.260 ;
        RECT 76.950 83.350 77.120 83.520 ;
        RECT 82.710 83.720 82.880 83.890 ;
        RECT 84.630 83.720 84.800 83.890 ;
        RECT 85.590 83.720 85.760 83.890 ;
        RECT 79.830 82.240 80.000 82.410 ;
        RECT 83.190 82.240 83.360 82.410 ;
        RECT 87.990 83.720 88.160 83.890 ;
        RECT 91.830 83.350 92.000 83.520 ;
        RECT 94.710 83.720 94.880 83.890 ;
        RECT 98.550 83.350 98.720 83.520 ;
        RECT 102.390 84.460 102.560 84.630 ;
        RECT 101.430 83.720 101.600 83.890 ;
        RECT 108.630 84.460 108.800 84.630 ;
        RECT 116.790 84.090 116.960 84.260 ;
        RECT 15.030 80.390 15.200 80.560 ;
      LAYER mcon ;
        RECT 6.510 77.720 6.680 77.890 ;
        RECT 6.950 77.720 7.120 77.890 ;
        RECT 7.360 77.720 7.530 77.890 ;
        RECT 7.790 77.720 7.960 77.890 ;
        RECT 8.230 77.720 8.400 77.890 ;
        RECT 8.640 77.720 8.810 77.890 ;
        RECT 10.350 77.720 10.520 77.890 ;
        RECT 10.790 77.720 10.960 77.890 ;
        RECT 11.200 77.720 11.370 77.890 ;
        RECT 11.630 77.720 11.800 77.890 ;
        RECT 12.070 77.720 12.240 77.890 ;
        RECT 12.480 77.720 12.650 77.890 ;
      LAYER L1M1_PR_C ;
        RECT 16.470 78.910 16.640 79.080 ;
      LAYER mcon ;
        RECT 15.430 77.730 15.600 77.900 ;
        RECT 15.790 77.730 15.960 77.900 ;
        RECT 16.150 77.730 16.320 77.900 ;
        RECT 16.510 77.730 16.680 77.900 ;
        RECT 18.030 77.720 18.200 77.890 ;
        RECT 18.470 77.720 18.640 77.890 ;
        RECT 18.880 77.720 19.050 77.890 ;
        RECT 19.310 77.720 19.480 77.890 ;
        RECT 19.750 77.720 19.920 77.890 ;
        RECT 20.160 77.720 20.330 77.890 ;
        RECT 21.340 77.730 21.510 77.900 ;
        RECT 21.780 77.730 21.950 77.900 ;
        RECT 22.220 77.730 22.390 77.900 ;
        RECT 22.630 77.730 22.800 77.900 ;
        RECT 23.630 77.730 23.800 77.900 ;
        RECT 23.990 77.730 24.160 77.900 ;
        RECT 24.350 77.730 24.520 77.900 ;
        RECT 25.270 77.730 25.440 77.900 ;
        RECT 25.630 77.730 25.800 77.900 ;
      LAYER L1M1_PR_C ;
        RECT 26.550 78.910 26.720 79.080 ;
      LAYER mcon ;
        RECT 30.230 77.730 30.400 77.900 ;
        RECT 30.590 77.730 30.760 77.900 ;
        RECT 30.950 77.730 31.120 77.900 ;
      LAYER L1M1_PR_C ;
        RECT 38.070 80.390 38.240 80.560 ;
      LAYER mcon ;
        RECT 34.200 77.730 34.370 77.900 ;
        RECT 34.560 77.730 34.730 77.900 ;
        RECT 34.920 77.730 35.090 77.900 ;
        RECT 36.810 77.730 36.980 77.900 ;
        RECT 37.170 77.730 37.340 77.900 ;
        RECT 37.530 77.730 37.700 77.900 ;
        RECT 39.150 77.720 39.320 77.890 ;
        RECT 39.590 77.720 39.760 77.890 ;
        RECT 40.000 77.720 40.170 77.890 ;
        RECT 40.430 77.720 40.600 77.890 ;
        RECT 40.870 77.720 41.040 77.890 ;
        RECT 41.280 77.720 41.450 77.890 ;
        RECT 42.830 77.730 43.000 77.900 ;
        RECT 43.190 77.730 43.360 77.900 ;
        RECT 43.550 77.730 43.720 77.900 ;
        RECT 44.470 77.730 44.640 77.900 ;
        RECT 44.830 77.730 45.000 77.900 ;
      LAYER L1M1_PR_C ;
        RECT 45.750 78.170 45.920 78.340 ;
      LAYER mcon ;
        RECT 49.430 77.730 49.600 77.900 ;
        RECT 49.790 77.730 49.960 77.900 ;
        RECT 50.150 77.730 50.320 77.900 ;
      LAYER L1M1_PR_C ;
        RECT 57.270 80.390 57.440 80.560 ;
      LAYER mcon ;
        RECT 53.400 77.730 53.570 77.900 ;
        RECT 53.760 77.730 53.930 77.900 ;
        RECT 54.120 77.730 54.290 77.900 ;
      LAYER L1M1_PR_C ;
        RECT 65.430 79.280 65.600 79.450 ;
        RECT 62.550 78.910 62.720 79.080 ;
      LAYER mcon ;
        RECT 56.010 77.730 56.180 77.900 ;
        RECT 56.370 77.730 56.540 77.900 ;
        RECT 56.730 77.730 56.900 77.900 ;
        RECT 58.350 77.720 58.520 77.890 ;
        RECT 58.790 77.720 58.960 77.890 ;
        RECT 59.200 77.720 59.370 77.890 ;
        RECT 59.630 77.720 59.800 77.890 ;
        RECT 60.070 77.720 60.240 77.890 ;
        RECT 60.480 77.720 60.650 77.890 ;
        RECT 61.560 77.730 61.730 77.900 ;
        RECT 61.920 77.730 62.090 77.900 ;
        RECT 62.280 77.730 62.450 77.900 ;
        RECT 63.120 77.730 63.290 77.900 ;
        RECT 63.480 77.730 63.650 77.900 ;
        RECT 63.840 77.730 64.010 77.900 ;
        RECT 64.680 77.730 64.850 77.900 ;
        RECT 65.040 77.730 65.210 77.900 ;
        RECT 65.400 77.730 65.570 77.900 ;
      LAYER L1M1_PR_C ;
        RECT 71.670 78.910 71.840 79.080 ;
      LAYER mcon ;
        RECT 66.990 77.720 67.160 77.890 ;
        RECT 67.430 77.720 67.600 77.890 ;
        RECT 67.840 77.720 68.010 77.890 ;
        RECT 68.270 77.720 68.440 77.890 ;
        RECT 68.710 77.720 68.880 77.890 ;
        RECT 69.120 77.720 69.290 77.890 ;
        RECT 72.120 77.730 72.290 77.900 ;
        RECT 72.480 77.730 72.650 77.900 ;
        RECT 72.840 77.730 73.010 77.900 ;
        RECT 73.200 77.730 73.370 77.900 ;
        RECT 73.560 77.730 73.730 77.900 ;
      LAYER L1M1_PR_C ;
        RECT 75.030 78.540 75.200 78.710 ;
        RECT 85.110 79.280 85.280 79.450 ;
      LAYER mcon ;
        RECT 74.610 77.730 74.780 77.900 ;
        RECT 74.970 77.730 75.140 77.900 ;
        RECT 75.330 77.730 75.500 77.900 ;
        RECT 75.690 77.730 75.860 77.900 ;
        RECT 76.050 77.730 76.220 77.900 ;
        RECT 77.550 77.720 77.720 77.890 ;
        RECT 77.990 77.720 78.160 77.890 ;
        RECT 78.400 77.720 78.570 77.890 ;
        RECT 78.830 77.720 79.000 77.890 ;
        RECT 79.270 77.720 79.440 77.890 ;
        RECT 79.680 77.720 79.850 77.890 ;
        RECT 81.240 77.730 81.410 77.900 ;
        RECT 81.600 77.730 81.770 77.900 ;
        RECT 81.960 77.730 82.130 77.900 ;
      LAYER L1M1_PR_C ;
        RECT 83.670 78.540 83.840 78.710 ;
      LAYER mcon ;
        RECT 82.800 77.730 82.970 77.900 ;
        RECT 83.160 77.730 83.330 77.900 ;
        RECT 83.520 77.730 83.690 77.900 ;
        RECT 84.360 77.730 84.530 77.900 ;
        RECT 84.720 77.730 84.890 77.900 ;
        RECT 85.080 77.730 85.250 77.900 ;
      LAYER L1M1_PR_C ;
        RECT 91.830 79.280 92.000 79.450 ;
      LAYER mcon ;
        RECT 86.140 77.730 86.310 77.900 ;
        RECT 86.580 77.730 86.750 77.900 ;
        RECT 87.020 77.730 87.190 77.900 ;
        RECT 87.430 77.730 87.600 77.900 ;
        RECT 87.960 77.730 88.130 77.900 ;
        RECT 88.320 77.730 88.490 77.900 ;
        RECT 88.680 77.730 88.850 77.900 ;
      LAYER L1M1_PR_C ;
        RECT 89.430 78.540 89.600 78.710 ;
      LAYER mcon ;
        RECT 89.520 77.730 89.690 77.900 ;
        RECT 89.880 77.730 90.050 77.900 ;
        RECT 90.240 77.730 90.410 77.900 ;
        RECT 91.080 77.730 91.250 77.900 ;
        RECT 91.440 77.730 91.610 77.900 ;
        RECT 91.800 77.730 91.970 77.900 ;
      LAYER L1M1_PR_C ;
        RECT 95.190 78.540 95.360 78.710 ;
        RECT 96.150 78.540 96.320 78.710 ;
      LAYER mcon ;
        RECT 92.860 77.730 93.030 77.900 ;
        RECT 93.300 77.730 93.470 77.900 ;
        RECT 93.740 77.730 93.910 77.900 ;
        RECT 94.150 77.730 94.320 77.900 ;
        RECT 94.660 77.730 94.830 77.900 ;
        RECT 95.020 77.730 95.190 77.900 ;
        RECT 95.380 77.730 95.550 77.900 ;
        RECT 96.630 77.730 96.800 77.900 ;
        RECT 96.990 77.730 97.160 77.900 ;
      LAYER L1M1_PR_C ;
        RECT 97.590 78.170 97.760 78.340 ;
        RECT 102.870 80.390 103.040 80.560 ;
        RECT 100.470 78.540 100.640 78.710 ;
        RECT 101.430 78.540 101.600 78.710 ;
      LAYER mcon ;
        RECT 98.140 77.730 98.310 77.900 ;
        RECT 98.580 77.730 98.750 77.900 ;
        RECT 99.020 77.730 99.190 77.900 ;
        RECT 99.430 77.730 99.600 77.900 ;
        RECT 99.940 77.730 100.110 77.900 ;
        RECT 100.300 77.730 100.470 77.900 ;
        RECT 100.660 77.730 100.830 77.900 ;
        RECT 101.910 77.730 102.080 77.900 ;
        RECT 102.270 77.730 102.440 77.900 ;
      LAYER L1M1_PR_C ;
        RECT 105.750 78.540 105.920 78.710 ;
        RECT 106.710 78.540 106.880 78.710 ;
      LAYER mcon ;
        RECT 103.420 77.730 103.590 77.900 ;
        RECT 103.860 77.730 104.030 77.900 ;
        RECT 104.300 77.730 104.470 77.900 ;
        RECT 104.710 77.730 104.880 77.900 ;
        RECT 105.220 77.730 105.390 77.900 ;
        RECT 105.580 77.730 105.750 77.900 ;
        RECT 105.940 77.730 106.110 77.900 ;
        RECT 107.190 77.730 107.360 77.900 ;
        RECT 107.550 77.730 107.720 77.900 ;
      LAYER L1M1_PR_C ;
        RECT 108.150 78.170 108.320 78.340 ;
        RECT 111.990 79.280 112.160 79.450 ;
      LAYER mcon ;
        RECT 108.700 77.730 108.870 77.900 ;
        RECT 109.140 77.730 109.310 77.900 ;
        RECT 109.580 77.730 109.750 77.900 ;
        RECT 109.990 77.730 110.160 77.900 ;
      LAYER L1M1_PR_C ;
        RECT 110.550 78.540 110.720 78.710 ;
      LAYER mcon ;
        RECT 110.950 77.730 111.120 77.900 ;
        RECT 111.310 77.730 111.480 77.900 ;
        RECT 111.670 77.730 111.840 77.900 ;
        RECT 112.030 77.730 112.200 77.900 ;
        RECT 113.020 77.730 113.190 77.900 ;
        RECT 113.460 77.730 113.630 77.900 ;
        RECT 113.900 77.730 114.070 77.900 ;
        RECT 114.310 77.730 114.480 77.900 ;
      LAYER L1M1_PR_C ;
        RECT 116.310 79.280 116.480 79.450 ;
        RECT 114.870 78.170 115.040 78.340 ;
      LAYER mcon ;
        RECT 115.270 77.730 115.440 77.900 ;
        RECT 115.630 77.730 115.800 77.900 ;
        RECT 115.990 77.730 116.160 77.900 ;
        RECT 116.350 77.730 116.520 77.900 ;
        RECT 117.340 77.730 117.510 77.900 ;
        RECT 117.780 77.730 117.950 77.900 ;
        RECT 118.220 77.730 118.390 77.900 ;
        RECT 118.630 77.730 118.800 77.900 ;
      LAYER L1M1_PR_C ;
        RECT 120.630 79.280 120.800 79.450 ;
        RECT 119.190 78.170 119.360 78.340 ;
      LAYER mcon ;
        RECT 119.590 77.730 119.760 77.900 ;
        RECT 119.950 77.730 120.120 77.900 ;
        RECT 120.310 77.730 120.480 77.900 ;
        RECT 120.670 77.730 120.840 77.900 ;
      LAYER L1M1_PR_C ;
        RECT 124.950 80.020 125.120 80.190 ;
      LAYER mcon ;
        RECT 121.660 77.730 121.830 77.900 ;
        RECT 122.100 77.730 122.270 77.900 ;
        RECT 122.540 77.730 122.710 77.900 ;
        RECT 122.950 77.730 123.120 77.900 ;
      LAYER L1M1_PR_C ;
        RECT 123.510 78.170 123.680 78.340 ;
      LAYER mcon ;
        RECT 123.910 77.730 124.080 77.900 ;
        RECT 124.270 77.730 124.440 77.900 ;
        RECT 124.630 77.730 124.800 77.900 ;
        RECT 124.990 77.730 125.160 77.900 ;
        RECT 126.510 77.720 126.680 77.890 ;
        RECT 126.950 77.720 127.120 77.890 ;
        RECT 127.360 77.720 127.530 77.890 ;
        RECT 127.790 77.720 127.960 77.890 ;
        RECT 128.230 77.720 128.400 77.890 ;
        RECT 128.640 77.720 128.810 77.890 ;
        RECT 130.350 77.720 130.520 77.890 ;
        RECT 130.790 77.720 130.960 77.890 ;
        RECT 131.200 77.720 131.370 77.890 ;
        RECT 131.630 77.720 131.800 77.890 ;
        RECT 132.070 77.720 132.240 77.890 ;
        RECT 132.480 77.720 132.650 77.890 ;
        RECT 134.190 77.720 134.360 77.890 ;
        RECT 134.630 77.720 134.800 77.890 ;
        RECT 135.040 77.720 135.210 77.890 ;
        RECT 135.470 77.720 135.640 77.890 ;
        RECT 135.910 77.720 136.080 77.890 ;
        RECT 136.320 77.720 136.490 77.890 ;
        RECT 138.030 77.720 138.200 77.890 ;
        RECT 138.470 77.720 138.640 77.890 ;
        RECT 138.880 77.720 139.050 77.890 ;
        RECT 139.310 77.720 139.480 77.890 ;
        RECT 139.750 77.720 139.920 77.890 ;
        RECT 140.160 77.720 140.330 77.890 ;
      LAYER L1M1_PR_C ;
        RECT 17.430 75.950 17.600 76.120 ;
        RECT 18.870 74.470 19.040 74.640 ;
        RECT 21.750 76.320 21.920 76.490 ;
        RECT 28.470 75.950 28.640 76.120 ;
        RECT 23.190 74.100 23.360 74.270 ;
        RECT 29.910 75.210 30.080 75.380 ;
        RECT 35.190 75.950 35.360 76.120 ;
        RECT 36.630 75.210 36.800 75.380 ;
        RECT 41.910 75.950 42.080 76.120 ;
        RECT 43.350 75.210 43.520 75.380 ;
        RECT 47.670 75.580 47.840 75.750 ;
        RECT 51.510 75.210 51.680 75.380 ;
        RECT 57.750 75.950 57.920 76.120 ;
        RECT 54.390 74.470 54.560 74.640 ;
        RECT 57.750 75.580 57.920 75.750 ;
        RECT 55.830 74.100 56.000 74.270 ;
        RECT 64.950 76.320 65.120 76.490 ;
        RECT 73.110 75.950 73.280 76.120 ;
        RECT 79.350 75.580 79.520 75.750 ;
        RECT 80.310 75.580 80.480 75.750 ;
        RECT 82.710 75.950 82.880 76.120 ;
        RECT 85.110 75.210 85.280 75.380 ;
        RECT 86.550 75.580 86.720 75.750 ;
        RECT 85.590 75.210 85.760 75.380 ;
        RECT 89.910 75.580 90.080 75.750 ;
        RECT 90.870 75.210 91.040 75.380 ;
        RECT 93.750 75.580 93.920 75.750 ;
        RECT 98.550 75.950 98.720 76.120 ;
        RECT 97.110 75.580 97.280 75.750 ;
        RECT 99.030 75.210 99.200 75.380 ;
        RECT 101.430 75.950 101.600 76.120 ;
        RECT 104.310 75.950 104.480 76.120 ;
        RECT 105.750 75.580 105.920 75.750 ;
        RECT 111.030 75.950 111.200 76.120 ;
        RECT 110.070 75.580 110.240 75.750 ;
        RECT 111.510 75.580 111.680 75.750 ;
        RECT 113.430 75.580 113.600 75.750 ;
        RECT 117.270 75.950 117.440 76.120 ;
        RECT 14.070 72.250 14.240 72.420 ;
      LAYER mcon ;
        RECT 6.510 69.580 6.680 69.750 ;
        RECT 6.950 69.580 7.120 69.750 ;
        RECT 7.360 69.580 7.530 69.750 ;
        RECT 7.790 69.580 7.960 69.750 ;
        RECT 8.230 69.580 8.400 69.750 ;
        RECT 8.640 69.580 8.810 69.750 ;
        RECT 9.820 69.590 9.990 69.760 ;
        RECT 10.260 69.590 10.430 69.760 ;
        RECT 10.700 69.590 10.870 69.760 ;
        RECT 11.110 69.590 11.280 69.760 ;
      LAYER L1M1_PR_C ;
        RECT 12.630 70.400 12.800 70.570 ;
        RECT 16.950 72.250 17.120 72.420 ;
      LAYER mcon ;
        RECT 13.030 69.590 13.200 69.760 ;
        RECT 13.390 69.590 13.560 69.760 ;
        RECT 13.750 69.590 13.920 69.760 ;
        RECT 14.110 69.590 14.280 69.760 ;
      LAYER L1M1_PR_C ;
        RECT 18.390 71.880 18.560 72.050 ;
      LAYER mcon ;
        RECT 15.100 69.590 15.270 69.760 ;
        RECT 15.540 69.590 15.710 69.760 ;
        RECT 15.980 69.590 16.150 69.760 ;
        RECT 16.390 69.590 16.560 69.760 ;
        RECT 17.350 69.590 17.520 69.760 ;
        RECT 17.710 69.590 17.880 69.760 ;
        RECT 18.070 69.590 18.240 69.760 ;
        RECT 18.430 69.590 18.600 69.760 ;
      LAYER L1M1_PR_C ;
        RECT 23.670 71.140 23.840 71.310 ;
        RECT 24.150 71.510 24.320 71.680 ;
        RECT 22.230 70.770 22.400 70.940 ;
        RECT 22.710 70.770 22.880 70.940 ;
      LAYER mcon ;
        RECT 19.420 69.590 19.590 69.760 ;
        RECT 19.860 69.590 20.030 69.760 ;
        RECT 20.300 69.590 20.470 69.760 ;
        RECT 20.710 69.590 20.880 69.760 ;
        RECT 21.500 69.590 21.670 69.760 ;
        RECT 21.860 69.590 22.030 69.760 ;
        RECT 22.220 69.590 22.390 69.760 ;
        RECT 22.580 69.590 22.750 69.760 ;
        RECT 22.940 69.590 23.110 69.760 ;
      LAYER L1M1_PR_C ;
        RECT 30.390 71.140 30.560 71.310 ;
        RECT 26.550 70.770 26.720 70.940 ;
      LAYER mcon ;
        RECT 23.830 69.590 24.000 69.760 ;
        RECT 24.190 69.590 24.360 69.760 ;
        RECT 24.700 69.590 24.870 69.760 ;
        RECT 25.140 69.590 25.310 69.760 ;
        RECT 25.580 69.590 25.750 69.760 ;
        RECT 25.990 69.590 26.160 69.760 ;
        RECT 26.520 69.590 26.690 69.760 ;
        RECT 26.880 69.590 27.050 69.760 ;
        RECT 27.240 69.590 27.410 69.760 ;
        RECT 28.080 69.590 28.250 69.760 ;
        RECT 28.440 69.590 28.610 69.760 ;
        RECT 28.800 69.590 28.970 69.760 ;
        RECT 29.640 69.590 29.810 69.760 ;
        RECT 30.000 69.590 30.170 69.760 ;
        RECT 30.360 69.590 30.530 69.760 ;
      LAYER L1M1_PR_C ;
        RECT 37.110 71.140 37.280 71.310 ;
        RECT 33.270 70.770 33.440 70.940 ;
      LAYER mcon ;
        RECT 31.420 69.590 31.590 69.760 ;
        RECT 31.860 69.590 32.030 69.760 ;
        RECT 32.300 69.590 32.470 69.760 ;
        RECT 32.710 69.590 32.880 69.760 ;
        RECT 33.240 69.590 33.410 69.760 ;
        RECT 33.600 69.590 33.770 69.760 ;
        RECT 33.960 69.590 34.130 69.760 ;
        RECT 34.800 69.590 34.970 69.760 ;
        RECT 35.160 69.590 35.330 69.760 ;
        RECT 35.520 69.590 35.690 69.760 ;
        RECT 36.360 69.590 36.530 69.760 ;
        RECT 36.720 69.590 36.890 69.760 ;
        RECT 37.080 69.590 37.250 69.760 ;
      LAYER L1M1_PR_C ;
        RECT 43.830 71.140 44.000 71.310 ;
        RECT 39.990 70.770 40.160 70.940 ;
      LAYER mcon ;
        RECT 38.140 69.590 38.310 69.760 ;
        RECT 38.580 69.590 38.750 69.760 ;
        RECT 39.020 69.590 39.190 69.760 ;
        RECT 39.430 69.590 39.600 69.760 ;
        RECT 39.960 69.590 40.130 69.760 ;
        RECT 40.320 69.590 40.490 69.760 ;
        RECT 40.680 69.590 40.850 69.760 ;
        RECT 41.520 69.590 41.690 69.760 ;
        RECT 41.880 69.590 42.050 69.760 ;
        RECT 42.240 69.590 42.410 69.760 ;
        RECT 43.080 69.590 43.250 69.760 ;
        RECT 43.440 69.590 43.610 69.760 ;
        RECT 43.800 69.590 43.970 69.760 ;
      LAYER L1M1_PR_C ;
        RECT 51.990 71.140 52.160 71.310 ;
      LAYER mcon ;
        RECT 44.860 69.590 45.030 69.760 ;
        RECT 45.300 69.590 45.470 69.760 ;
        RECT 45.740 69.590 45.910 69.760 ;
        RECT 46.150 69.590 46.320 69.760 ;
        RECT 48.120 69.590 48.290 69.760 ;
        RECT 48.480 69.590 48.650 69.760 ;
        RECT 48.840 69.590 49.010 69.760 ;
      LAYER L1M1_PR_C ;
        RECT 49.590 70.400 49.760 70.570 ;
      LAYER mcon ;
        RECT 49.680 69.590 49.850 69.760 ;
        RECT 50.040 69.590 50.210 69.760 ;
        RECT 50.400 69.590 50.570 69.760 ;
        RECT 51.240 69.590 51.410 69.760 ;
        RECT 51.600 69.590 51.770 69.760 ;
        RECT 51.960 69.590 52.130 69.760 ;
      LAYER L1M1_PR_C ;
        RECT 56.790 71.880 56.960 72.050 ;
        RECT 54.870 71.140 55.040 71.310 ;
        RECT 56.310 71.140 56.480 71.310 ;
      LAYER mcon ;
        RECT 53.020 69.590 53.190 69.760 ;
        RECT 53.460 69.590 53.630 69.760 ;
        RECT 53.900 69.590 54.070 69.760 ;
        RECT 54.310 69.590 54.480 69.760 ;
        RECT 54.830 69.590 55.000 69.760 ;
        RECT 55.190 69.590 55.360 69.760 ;
        RECT 55.550 69.590 55.720 69.760 ;
      LAYER L1M1_PR_C ;
        RECT 63.510 71.140 63.680 71.310 ;
      LAYER mcon ;
        RECT 56.470 69.590 56.640 69.760 ;
        RECT 56.830 69.590 57.000 69.760 ;
        RECT 57.340 69.590 57.510 69.760 ;
        RECT 57.780 69.590 57.950 69.760 ;
        RECT 58.220 69.590 58.390 69.760 ;
        RECT 58.630 69.590 58.800 69.760 ;
        RECT 59.640 69.590 59.810 69.760 ;
        RECT 60.000 69.590 60.170 69.760 ;
        RECT 60.360 69.590 60.530 69.760 ;
      LAYER L1M1_PR_C ;
        RECT 61.590 70.400 61.760 70.570 ;
      LAYER mcon ;
        RECT 61.200 69.590 61.370 69.760 ;
        RECT 61.560 69.590 61.730 69.760 ;
        RECT 61.920 69.590 62.090 69.760 ;
        RECT 62.760 69.590 62.930 69.760 ;
        RECT 63.120 69.590 63.290 69.760 ;
        RECT 63.480 69.590 63.650 69.760 ;
      LAYER L1M1_PR_C ;
        RECT 70.230 71.140 70.400 71.310 ;
        RECT 66.390 70.770 66.560 70.940 ;
      LAYER mcon ;
        RECT 64.540 69.590 64.710 69.760 ;
        RECT 64.980 69.590 65.150 69.760 ;
        RECT 65.420 69.590 65.590 69.760 ;
        RECT 65.830 69.590 66.000 69.760 ;
        RECT 66.360 69.590 66.530 69.760 ;
        RECT 66.720 69.590 66.890 69.760 ;
        RECT 67.080 69.590 67.250 69.760 ;
        RECT 67.920 69.590 68.090 69.760 ;
        RECT 68.280 69.590 68.450 69.760 ;
        RECT 68.640 69.590 68.810 69.760 ;
        RECT 69.480 69.590 69.650 69.760 ;
        RECT 69.840 69.590 70.010 69.760 ;
        RECT 70.200 69.590 70.370 69.760 ;
      LAYER L1M1_PR_C ;
        RECT 74.070 71.140 74.240 71.310 ;
        RECT 73.110 70.770 73.280 70.940 ;
      LAYER mcon ;
        RECT 71.260 69.590 71.430 69.760 ;
        RECT 71.700 69.590 71.870 69.760 ;
        RECT 72.140 69.590 72.310 69.760 ;
        RECT 72.550 69.590 72.720 69.760 ;
        RECT 73.080 69.590 73.250 69.760 ;
        RECT 73.440 69.590 73.610 69.760 ;
      LAYER L1M1_PR_C ;
        RECT 79.350 71.140 79.520 71.310 ;
        RECT 79.830 72.250 80.000 72.420 ;
        RECT 76.950 70.770 77.120 70.940 ;
      LAYER mcon ;
        RECT 74.620 69.590 74.790 69.760 ;
        RECT 75.060 69.590 75.230 69.760 ;
        RECT 75.500 69.590 75.670 69.760 ;
        RECT 75.910 69.590 76.080 69.760 ;
        RECT 77.180 69.590 77.350 69.760 ;
        RECT 77.540 69.590 77.710 69.760 ;
        RECT 77.900 69.590 78.070 69.760 ;
        RECT 78.260 69.590 78.430 69.760 ;
        RECT 78.620 69.590 78.790 69.760 ;
      LAYER L1M1_PR_C ;
        RECT 86.070 71.140 86.240 71.310 ;
      LAYER mcon ;
        RECT 79.510 69.590 79.680 69.760 ;
        RECT 79.870 69.590 80.040 69.760 ;
        RECT 80.380 69.590 80.550 69.760 ;
        RECT 80.820 69.590 80.990 69.760 ;
        RECT 81.260 69.590 81.430 69.760 ;
        RECT 81.670 69.590 81.840 69.760 ;
        RECT 82.200 69.590 82.370 69.760 ;
        RECT 82.560 69.590 82.730 69.760 ;
        RECT 82.920 69.590 83.090 69.760 ;
      LAYER L1M1_PR_C ;
        RECT 84.150 70.400 84.320 70.570 ;
      LAYER mcon ;
        RECT 83.760 69.590 83.930 69.760 ;
        RECT 84.120 69.590 84.290 69.760 ;
        RECT 84.480 69.590 84.650 69.760 ;
        RECT 85.320 69.590 85.490 69.760 ;
        RECT 85.680 69.590 85.850 69.760 ;
        RECT 86.040 69.590 86.210 69.760 ;
      LAYER L1M1_PR_C ;
        RECT 92.790 71.140 92.960 71.310 ;
      LAYER mcon ;
        RECT 87.100 69.590 87.270 69.760 ;
        RECT 87.540 69.590 87.710 69.760 ;
        RECT 87.980 69.590 88.150 69.760 ;
        RECT 88.390 69.590 88.560 69.760 ;
        RECT 88.920 69.590 89.090 69.760 ;
        RECT 89.280 69.590 89.450 69.760 ;
        RECT 89.640 69.590 89.810 69.760 ;
      LAYER L1M1_PR_C ;
        RECT 91.350 70.400 91.520 70.570 ;
      LAYER mcon ;
        RECT 90.480 69.590 90.650 69.760 ;
        RECT 90.840 69.590 91.010 69.760 ;
        RECT 91.200 69.590 91.370 69.760 ;
        RECT 92.040 69.590 92.210 69.760 ;
        RECT 92.400 69.590 92.570 69.760 ;
        RECT 92.760 69.590 92.930 69.760 ;
      LAYER L1M1_PR_C ;
        RECT 96.630 72.250 96.800 72.420 ;
      LAYER mcon ;
        RECT 93.820 69.590 93.990 69.760 ;
        RECT 94.260 69.590 94.430 69.760 ;
        RECT 94.700 69.590 94.870 69.760 ;
        RECT 95.110 69.590 95.280 69.760 ;
        RECT 95.640 69.590 95.810 69.760 ;
        RECT 96.000 69.590 96.170 69.760 ;
      LAYER L1M1_PR_C ;
        RECT 101.430 71.140 101.600 71.310 ;
        RECT 99.030 70.770 99.200 70.940 ;
        RECT 100.470 70.770 100.640 70.940 ;
        RECT 101.910 70.770 102.080 70.940 ;
      LAYER mcon ;
        RECT 97.180 69.590 97.350 69.760 ;
        RECT 97.620 69.590 97.790 69.760 ;
        RECT 98.060 69.590 98.230 69.760 ;
        RECT 98.470 69.590 98.640 69.760 ;
        RECT 99.260 69.590 99.430 69.760 ;
        RECT 99.620 69.590 99.790 69.760 ;
        RECT 99.980 69.590 100.150 69.760 ;
        RECT 100.340 69.590 100.510 69.760 ;
        RECT 100.700 69.590 100.870 69.760 ;
      LAYER L1M1_PR_C ;
        RECT 104.310 70.770 104.480 70.940 ;
        RECT 106.230 70.770 106.400 70.940 ;
      LAYER mcon ;
        RECT 101.590 69.590 101.760 69.760 ;
        RECT 101.950 69.590 102.120 69.760 ;
        RECT 102.460 69.590 102.630 69.760 ;
        RECT 102.900 69.590 103.070 69.760 ;
        RECT 103.340 69.590 103.510 69.760 ;
        RECT 103.750 69.590 103.920 69.760 ;
        RECT 104.280 69.590 104.450 69.760 ;
        RECT 104.640 69.590 104.810 69.760 ;
        RECT 105.000 69.590 105.170 69.760 ;
        RECT 105.360 69.590 105.530 69.760 ;
      LAYER L1M1_PR_C ;
        RECT 110.550 71.880 110.720 72.050 ;
        RECT 108.630 71.140 108.800 71.310 ;
        RECT 110.070 71.140 110.240 71.310 ;
        RECT 106.230 70.030 106.400 70.200 ;
      LAYER mcon ;
        RECT 106.780 69.590 106.950 69.760 ;
        RECT 107.220 69.590 107.390 69.760 ;
        RECT 107.660 69.590 107.830 69.760 ;
        RECT 108.070 69.590 108.240 69.760 ;
        RECT 108.590 69.590 108.760 69.760 ;
        RECT 108.950 69.590 109.120 69.760 ;
        RECT 109.310 69.590 109.480 69.760 ;
      LAYER L1M1_PR_C ;
        RECT 113.910 72.250 114.080 72.420 ;
        RECT 112.950 70.770 113.120 70.940 ;
      LAYER mcon ;
        RECT 110.230 69.590 110.400 69.760 ;
        RECT 110.590 69.590 110.760 69.760 ;
        RECT 111.100 69.590 111.270 69.760 ;
        RECT 111.540 69.590 111.710 69.760 ;
        RECT 111.980 69.590 112.150 69.760 ;
        RECT 112.390 69.590 112.560 69.760 ;
        RECT 112.920 69.590 113.090 69.760 ;
        RECT 113.280 69.590 113.450 69.760 ;
      LAYER L1M1_PR_C ;
        RECT 120.150 71.140 120.320 71.310 ;
      LAYER mcon ;
        RECT 114.460 69.590 114.630 69.760 ;
        RECT 114.900 69.590 115.070 69.760 ;
        RECT 115.340 69.590 115.510 69.760 ;
        RECT 115.750 69.590 115.920 69.760 ;
        RECT 116.280 69.590 116.450 69.760 ;
        RECT 116.640 69.590 116.810 69.760 ;
        RECT 117.000 69.590 117.170 69.760 ;
      LAYER L1M1_PR_C ;
        RECT 118.710 70.400 118.880 70.570 ;
      LAYER mcon ;
        RECT 117.840 69.590 118.010 69.760 ;
        RECT 118.200 69.590 118.370 69.760 ;
        RECT 118.560 69.590 118.730 69.760 ;
        RECT 119.400 69.590 119.570 69.760 ;
        RECT 119.760 69.590 119.930 69.760 ;
        RECT 120.120 69.590 120.290 69.760 ;
        RECT 121.180 69.590 121.350 69.760 ;
        RECT 121.620 69.590 121.790 69.760 ;
        RECT 122.060 69.590 122.230 69.760 ;
        RECT 122.470 69.590 122.640 69.760 ;
      LAYER L1M1_PR_C ;
        RECT 124.470 70.770 124.640 70.940 ;
        RECT 130.710 71.880 130.880 72.050 ;
        RECT 123.030 70.030 123.200 70.200 ;
      LAYER mcon ;
        RECT 123.430 69.590 123.600 69.760 ;
        RECT 123.790 69.590 123.960 69.760 ;
        RECT 124.150 69.590 124.320 69.760 ;
        RECT 124.510 69.590 124.680 69.760 ;
        RECT 126.030 69.580 126.200 69.750 ;
        RECT 126.470 69.580 126.640 69.750 ;
        RECT 126.880 69.580 127.050 69.750 ;
        RECT 127.310 69.580 127.480 69.750 ;
        RECT 127.750 69.580 127.920 69.750 ;
        RECT 128.160 69.580 128.330 69.750 ;
      LAYER L1M1_PR_C ;
        RECT 129.270 70.030 129.440 70.200 ;
      LAYER mcon ;
        RECT 129.670 69.590 129.840 69.760 ;
        RECT 130.030 69.590 130.200 69.760 ;
        RECT 130.390 69.590 130.560 69.760 ;
        RECT 130.750 69.590 130.920 69.760 ;
        RECT 132.270 69.580 132.440 69.750 ;
        RECT 132.710 69.580 132.880 69.750 ;
        RECT 133.120 69.580 133.290 69.750 ;
        RECT 133.550 69.580 133.720 69.750 ;
        RECT 133.990 69.580 134.160 69.750 ;
        RECT 134.400 69.580 134.570 69.750 ;
        RECT 136.110 69.580 136.280 69.750 ;
        RECT 136.550 69.580 136.720 69.750 ;
        RECT 136.960 69.580 137.130 69.750 ;
        RECT 137.390 69.580 137.560 69.750 ;
        RECT 137.830 69.580 138.000 69.750 ;
        RECT 138.240 69.580 138.410 69.750 ;
        RECT 139.420 69.590 139.590 69.760 ;
        RECT 139.860 69.590 140.030 69.760 ;
        RECT 140.300 69.590 140.470 69.760 ;
        RECT 140.710 69.590 140.880 69.760 ;
      LAYER L1M1_PR_C ;
        RECT 10.710 67.440 10.880 67.610 ;
        RECT 9.270 66.330 9.440 66.500 ;
        RECT 15.510 67.440 15.680 67.610 ;
        RECT 14.070 67.070 14.240 67.240 ;
        RECT 15.030 67.070 15.200 67.240 ;
        RECT 19.830 68.180 20.000 68.350 ;
        RECT 18.390 67.440 18.560 67.610 ;
        RECT 19.830 67.440 20.000 67.610 ;
        RECT 24.630 67.810 24.800 67.980 ;
        RECT 26.070 67.070 26.240 67.240 ;
        RECT 28.950 67.440 29.120 67.610 ;
        RECT 32.790 67.070 32.960 67.240 ;
        RECT 35.670 67.440 35.840 67.610 ;
        RECT 36.630 67.440 36.800 67.610 ;
        RECT 39.030 67.440 39.200 67.610 ;
        RECT 42.870 67.070 43.040 67.240 ;
        RECT 50.070 67.810 50.240 67.980 ;
        RECT 51.990 67.070 52.160 67.240 ;
        RECT 57.750 67.440 57.920 67.610 ;
        RECT 61.590 67.070 61.760 67.240 ;
        RECT 64.470 67.440 64.640 67.610 ;
        RECT 68.310 67.070 68.480 67.240 ;
        RECT 71.190 67.440 71.360 67.610 ;
        RECT 75.030 67.070 75.200 67.240 ;
        RECT 79.830 68.180 80.000 68.350 ;
        RECT 78.390 67.440 78.560 67.610 ;
        RECT 80.310 67.810 80.480 67.980 ;
        RECT 83.190 68.180 83.360 68.350 ;
        RECT 80.790 66.700 80.960 66.870 ;
        RECT 84.150 67.440 84.320 67.610 ;
        RECT 86.070 67.440 86.240 67.610 ;
        RECT 87.030 67.440 87.200 67.610 ;
        RECT 95.190 67.440 95.360 67.610 ;
        RECT 103.350 67.810 103.520 67.980 ;
        RECT 113.430 68.180 113.600 68.350 ;
        RECT 111.510 67.440 111.680 67.610 ;
        RECT 111.990 67.440 112.160 67.610 ;
        RECT 106.710 65.960 106.880 66.130 ;
        RECT 113.910 67.070 114.080 67.240 ;
        RECT 116.310 67.440 116.480 67.610 ;
        RECT 120.150 67.070 120.320 67.240 ;
        RECT 130.710 68.180 130.880 68.350 ;
        RECT 123.030 67.440 123.200 67.610 ;
        RECT 124.470 67.070 124.640 67.240 ;
        RECT 124.950 65.960 125.120 66.130 ;
        RECT 132.150 67.440 132.320 67.610 ;
        RECT 125.430 65.960 125.600 66.130 ;
        RECT 135.990 67.810 136.160 67.980 ;
        RECT 135.510 67.440 135.680 67.610 ;
        RECT 9.750 63.370 9.920 63.540 ;
        RECT 8.790 63.000 8.960 63.170 ;
        RECT 9.270 63.000 9.440 63.170 ;
      LAYER mcon ;
        RECT 5.980 61.450 6.150 61.620 ;
        RECT 6.420 61.450 6.590 61.620 ;
        RECT 6.860 61.450 7.030 61.620 ;
        RECT 7.270 61.450 7.440 61.620 ;
        RECT 7.790 61.450 7.960 61.620 ;
        RECT 8.150 61.450 8.320 61.620 ;
        RECT 8.510 61.450 8.680 61.620 ;
      LAYER L1M1_PR_C ;
        RECT 12.630 62.630 12.800 62.800 ;
        RECT 14.070 62.630 14.240 62.800 ;
      LAYER mcon ;
        RECT 9.430 61.450 9.600 61.620 ;
        RECT 9.790 61.450 9.960 61.620 ;
        RECT 10.300 61.450 10.470 61.620 ;
        RECT 10.740 61.450 10.910 61.620 ;
        RECT 11.180 61.450 11.350 61.620 ;
        RECT 11.590 61.450 11.760 61.620 ;
      LAYER L1M1_PR_C ;
        RECT 13.590 62.260 13.760 62.430 ;
      LAYER mcon ;
        RECT 12.120 61.450 12.290 61.620 ;
        RECT 12.480 61.450 12.650 61.620 ;
        RECT 12.840 61.450 13.010 61.620 ;
        RECT 13.200 61.450 13.370 61.620 ;
      LAYER L1M1_PR_C ;
        RECT 18.870 63.000 19.040 63.170 ;
        RECT 17.430 62.630 17.600 62.800 ;
        RECT 17.910 62.630 18.080 62.800 ;
        RECT 19.350 62.630 19.520 62.800 ;
      LAYER mcon ;
        RECT 14.620 61.450 14.790 61.620 ;
        RECT 15.060 61.450 15.230 61.620 ;
        RECT 15.500 61.450 15.670 61.620 ;
        RECT 15.910 61.450 16.080 61.620 ;
        RECT 16.700 61.450 16.870 61.620 ;
        RECT 17.060 61.450 17.230 61.620 ;
        RECT 17.420 61.450 17.590 61.620 ;
        RECT 17.780 61.450 17.950 61.620 ;
        RECT 18.140 61.450 18.310 61.620 ;
        RECT 19.030 61.450 19.200 61.620 ;
        RECT 19.390 61.450 19.560 61.620 ;
        RECT 19.900 61.450 20.070 61.620 ;
        RECT 20.340 61.450 20.510 61.620 ;
        RECT 20.780 61.450 20.950 61.620 ;
        RECT 21.190 61.450 21.360 61.620 ;
      LAYER L1M1_PR_C ;
        RECT 24.630 63.370 24.800 63.540 ;
      LAYER mcon ;
        RECT 22.190 61.450 22.360 61.620 ;
        RECT 22.550 61.450 22.720 61.620 ;
        RECT 22.910 61.450 23.080 61.620 ;
        RECT 23.830 61.450 24.000 61.620 ;
        RECT 24.190 61.450 24.360 61.620 ;
      LAYER L1M1_PR_C ;
        RECT 25.110 62.630 25.280 62.800 ;
      LAYER mcon ;
        RECT 28.790 61.450 28.960 61.620 ;
        RECT 29.150 61.450 29.320 61.620 ;
        RECT 29.510 61.450 29.680 61.620 ;
        RECT 32.760 61.450 32.930 61.620 ;
        RECT 33.120 61.450 33.290 61.620 ;
        RECT 33.480 61.450 33.650 61.620 ;
      LAYER L1M1_PR_C ;
        RECT 36.630 61.890 36.800 62.060 ;
        RECT 42.870 63.000 43.040 63.170 ;
      LAYER mcon ;
        RECT 35.370 61.450 35.540 61.620 ;
        RECT 35.730 61.450 35.900 61.620 ;
        RECT 36.090 61.450 36.260 61.620 ;
        RECT 37.180 61.450 37.350 61.620 ;
        RECT 37.620 61.450 37.790 61.620 ;
        RECT 38.060 61.450 38.230 61.620 ;
        RECT 38.470 61.450 38.640 61.620 ;
        RECT 39.000 61.450 39.170 61.620 ;
        RECT 39.360 61.450 39.530 61.620 ;
        RECT 39.720 61.450 39.890 61.620 ;
      LAYER L1M1_PR_C ;
        RECT 41.430 62.260 41.600 62.430 ;
      LAYER mcon ;
        RECT 40.560 61.450 40.730 61.620 ;
        RECT 40.920 61.450 41.090 61.620 ;
        RECT 41.280 61.450 41.450 61.620 ;
        RECT 42.120 61.450 42.290 61.620 ;
        RECT 42.480 61.450 42.650 61.620 ;
        RECT 42.840 61.450 43.010 61.620 ;
        RECT 43.900 61.450 44.070 61.620 ;
        RECT 44.340 61.450 44.510 61.620 ;
        RECT 44.780 61.450 44.950 61.620 ;
        RECT 45.190 61.450 45.360 61.620 ;
      LAYER L1M1_PR_C ;
        RECT 49.590 63.370 49.760 63.540 ;
      LAYER mcon ;
        RECT 47.150 61.450 47.320 61.620 ;
        RECT 47.510 61.450 47.680 61.620 ;
        RECT 47.870 61.450 48.040 61.620 ;
        RECT 48.790 61.450 48.960 61.620 ;
        RECT 49.150 61.450 49.320 61.620 ;
      LAYER L1M1_PR_C ;
        RECT 50.070 62.630 50.240 62.800 ;
      LAYER mcon ;
        RECT 53.750 61.450 53.920 61.620 ;
        RECT 54.110 61.450 54.280 61.620 ;
        RECT 54.470 61.450 54.640 61.620 ;
      LAYER L1M1_PR_C ;
        RECT 61.590 64.110 61.760 64.280 ;
      LAYER mcon ;
        RECT 57.720 61.450 57.890 61.620 ;
        RECT 58.080 61.450 58.250 61.620 ;
        RECT 58.440 61.450 58.610 61.620 ;
      LAYER L1M1_PR_C ;
        RECT 63.990 62.630 64.160 62.800 ;
        RECT 65.910 62.630 66.080 62.800 ;
      LAYER mcon ;
        RECT 60.330 61.450 60.500 61.620 ;
        RECT 60.690 61.450 60.860 61.620 ;
        RECT 61.050 61.450 61.220 61.620 ;
        RECT 62.140 61.450 62.310 61.620 ;
        RECT 62.580 61.450 62.750 61.620 ;
        RECT 63.020 61.450 63.190 61.620 ;
        RECT 63.430 61.450 63.600 61.620 ;
        RECT 63.960 61.450 64.130 61.620 ;
        RECT 64.320 61.450 64.490 61.620 ;
        RECT 64.680 61.450 64.850 61.620 ;
        RECT 65.040 61.450 65.210 61.620 ;
      LAYER L1M1_PR_C ;
        RECT 69.750 64.110 69.920 64.280 ;
        RECT 65.910 61.890 66.080 62.060 ;
      LAYER mcon ;
        RECT 66.460 61.450 66.630 61.620 ;
        RECT 66.900 61.450 67.070 61.620 ;
        RECT 67.340 61.450 67.510 61.620 ;
        RECT 67.750 61.450 67.920 61.620 ;
      LAYER L1M1_PR_C ;
        RECT 68.310 61.890 68.480 62.060 ;
      LAYER mcon ;
        RECT 68.760 61.450 68.930 61.620 ;
        RECT 69.120 61.450 69.290 61.620 ;
        RECT 69.480 61.450 69.650 61.620 ;
        RECT 69.840 61.450 70.010 61.620 ;
        RECT 70.200 61.450 70.370 61.620 ;
      LAYER L1M1_PR_C ;
        RECT 71.670 62.630 71.840 62.800 ;
        RECT 71.190 62.260 71.360 62.430 ;
      LAYER mcon ;
        RECT 71.250 61.450 71.420 61.620 ;
        RECT 71.610 61.450 71.780 61.620 ;
        RECT 71.970 61.450 72.140 61.620 ;
        RECT 72.330 61.450 72.500 61.620 ;
        RECT 72.690 61.450 72.860 61.620 ;
      LAYER L1M1_PR_C ;
        RECT 79.350 63.000 79.520 63.170 ;
        RECT 75.510 62.630 75.680 62.800 ;
      LAYER mcon ;
        RECT 73.660 61.450 73.830 61.620 ;
        RECT 74.100 61.450 74.270 61.620 ;
        RECT 74.540 61.450 74.710 61.620 ;
        RECT 74.950 61.450 75.120 61.620 ;
        RECT 75.480 61.450 75.650 61.620 ;
        RECT 75.840 61.450 76.010 61.620 ;
        RECT 76.200 61.450 76.370 61.620 ;
        RECT 77.040 61.450 77.210 61.620 ;
        RECT 77.400 61.450 77.570 61.620 ;
        RECT 77.760 61.450 77.930 61.620 ;
        RECT 78.600 61.450 78.770 61.620 ;
        RECT 78.960 61.450 79.130 61.620 ;
        RECT 79.320 61.450 79.490 61.620 ;
      LAYER L1M1_PR_C ;
        RECT 83.190 64.110 83.360 64.280 ;
        RECT 82.710 62.630 82.880 62.800 ;
      LAYER mcon ;
        RECT 80.380 61.450 80.550 61.620 ;
        RECT 80.820 61.450 80.990 61.620 ;
        RECT 81.260 61.450 81.430 61.620 ;
        RECT 81.670 61.450 81.840 61.620 ;
        RECT 82.200 61.450 82.370 61.620 ;
        RECT 82.560 61.450 82.730 61.620 ;
      LAYER L1M1_PR_C ;
        RECT 87.030 64.110 87.200 64.280 ;
        RECT 87.990 63.000 88.160 63.170 ;
        RECT 85.590 62.630 85.760 62.800 ;
        RECT 88.950 63.000 89.120 63.170 ;
        RECT 86.550 62.630 86.720 62.800 ;
      LAYER mcon ;
        RECT 83.740 61.450 83.910 61.620 ;
        RECT 84.180 61.450 84.350 61.620 ;
        RECT 84.620 61.450 84.790 61.620 ;
        RECT 85.030 61.450 85.200 61.620 ;
        RECT 87.640 61.450 87.810 61.620 ;
        RECT 88.000 61.450 88.170 61.620 ;
        RECT 88.360 61.450 88.530 61.620 ;
      LAYER L1M1_PR_C ;
        RECT 95.670 63.000 95.840 63.170 ;
      LAYER mcon ;
        RECT 89.500 61.450 89.670 61.620 ;
        RECT 89.940 61.450 90.110 61.620 ;
        RECT 90.380 61.450 90.550 61.620 ;
        RECT 90.790 61.450 90.960 61.620 ;
        RECT 91.800 61.450 91.970 61.620 ;
        RECT 92.160 61.450 92.330 61.620 ;
        RECT 92.520 61.450 92.690 61.620 ;
      LAYER L1M1_PR_C ;
        RECT 94.230 62.260 94.400 62.430 ;
      LAYER mcon ;
        RECT 93.360 61.450 93.530 61.620 ;
        RECT 93.720 61.450 93.890 61.620 ;
        RECT 94.080 61.450 94.250 61.620 ;
        RECT 94.920 61.450 95.090 61.620 ;
        RECT 95.280 61.450 95.450 61.620 ;
        RECT 95.640 61.450 95.810 61.620 ;
      LAYER L1M1_PR_C ;
        RECT 100.950 64.110 101.120 64.280 ;
        RECT 98.550 62.630 98.720 62.800 ;
        RECT 99.990 62.630 100.160 62.800 ;
        RECT 101.430 62.630 101.600 62.800 ;
      LAYER mcon ;
        RECT 96.700 61.450 96.870 61.620 ;
        RECT 97.140 61.450 97.310 61.620 ;
        RECT 97.580 61.450 97.750 61.620 ;
        RECT 97.990 61.450 98.160 61.620 ;
        RECT 98.780 61.450 98.950 61.620 ;
        RECT 99.140 61.450 99.310 61.620 ;
        RECT 99.500 61.450 99.670 61.620 ;
        RECT 99.860 61.450 100.030 61.620 ;
        RECT 100.220 61.450 100.390 61.620 ;
        RECT 101.110 61.450 101.280 61.620 ;
        RECT 101.470 61.450 101.640 61.620 ;
        RECT 102.510 61.440 102.680 61.610 ;
        RECT 102.950 61.440 103.120 61.610 ;
        RECT 103.360 61.440 103.530 61.610 ;
        RECT 103.790 61.440 103.960 61.610 ;
        RECT 104.230 61.440 104.400 61.610 ;
        RECT 104.640 61.440 104.810 61.610 ;
        RECT 106.670 61.450 106.840 61.620 ;
        RECT 107.030 61.450 107.200 61.620 ;
        RECT 107.390 61.450 107.560 61.620 ;
        RECT 108.310 61.450 108.480 61.620 ;
        RECT 108.670 61.450 108.840 61.620 ;
      LAYER L1M1_PR_C ;
        RECT 109.590 61.890 109.760 62.060 ;
      LAYER mcon ;
        RECT 113.270 61.450 113.440 61.620 ;
        RECT 113.630 61.450 113.800 61.620 ;
        RECT 113.990 61.450 114.160 61.620 ;
      LAYER L1M1_PR_C ;
        RECT 117.750 62.260 117.920 62.430 ;
        RECT 121.110 63.370 121.280 63.540 ;
      LAYER mcon ;
        RECT 117.240 61.450 117.410 61.620 ;
        RECT 117.600 61.450 117.770 61.620 ;
        RECT 117.960 61.450 118.130 61.620 ;
        RECT 119.850 61.450 120.020 61.620 ;
        RECT 120.210 61.450 120.380 61.620 ;
        RECT 120.570 61.450 120.740 61.620 ;
        RECT 121.660 61.450 121.830 61.620 ;
        RECT 122.100 61.450 122.270 61.620 ;
        RECT 122.540 61.450 122.710 61.620 ;
        RECT 122.950 61.450 123.120 61.620 ;
        RECT 123.950 61.450 124.120 61.620 ;
        RECT 124.310 61.450 124.480 61.620 ;
        RECT 124.670 61.450 124.840 61.620 ;
        RECT 125.590 61.450 125.760 61.620 ;
        RECT 125.950 61.450 126.120 61.620 ;
      LAYER L1M1_PR_C ;
        RECT 126.870 61.890 127.040 62.060 ;
      LAYER mcon ;
        RECT 130.550 61.450 130.720 61.620 ;
        RECT 130.910 61.450 131.080 61.620 ;
        RECT 131.270 61.450 131.440 61.620 ;
      LAYER L1M1_PR_C ;
        RECT 135.030 62.260 135.200 62.430 ;
        RECT 138.390 64.110 138.560 64.280 ;
      LAYER mcon ;
        RECT 134.520 61.450 134.690 61.620 ;
        RECT 134.880 61.450 135.050 61.620 ;
        RECT 135.240 61.450 135.410 61.620 ;
        RECT 137.130 61.450 137.300 61.620 ;
        RECT 137.490 61.450 137.660 61.620 ;
        RECT 137.850 61.450 138.020 61.620 ;
        RECT 138.940 61.450 139.110 61.620 ;
        RECT 139.380 61.450 139.550 61.620 ;
        RECT 139.820 61.450 139.990 61.620 ;
        RECT 140.230 61.450 140.400 61.620 ;
      LAYER L1M1_PR_C ;
        RECT 11.190 60.040 11.360 60.210 ;
        RECT 19.350 59.670 19.520 59.840 ;
        RECT 22.710 59.670 22.880 59.840 ;
        RECT 25.110 57.820 25.280 57.990 ;
        RECT 29.430 59.300 29.600 59.470 ;
        RECT 26.550 57.820 26.720 57.990 ;
        RECT 33.270 58.930 33.440 59.100 ;
        RECT 36.150 59.300 36.320 59.470 ;
        RECT 39.990 58.930 40.160 59.100 ;
        RECT 42.870 59.300 43.040 59.470 ;
        RECT 46.710 58.930 46.880 59.100 ;
        RECT 52.470 59.670 52.640 59.840 ;
        RECT 53.910 58.930 54.080 59.100 ;
        RECT 56.790 58.930 56.960 59.100 ;
        RECT 57.750 58.930 57.920 59.100 ;
        RECT 58.710 58.560 58.880 58.730 ;
        RECT 59.190 57.820 59.360 57.990 ;
        RECT 65.430 59.300 65.600 59.470 ;
        RECT 76.950 60.040 77.120 60.210 ;
        RECT 79.350 59.300 79.520 59.470 ;
        RECT 83.190 58.930 83.360 59.100 ;
        RECT 87.990 59.300 88.160 59.470 ;
        RECT 91.830 58.930 92.000 59.100 ;
        RECT 94.710 59.300 94.880 59.470 ;
        RECT 98.550 58.930 98.720 59.100 ;
        RECT 107.190 60.040 107.360 60.210 ;
        RECT 103.830 59.300 104.000 59.470 ;
        RECT 103.830 58.930 104.000 59.100 ;
        RECT 111.990 59.670 112.160 59.840 ;
        RECT 113.430 58.930 113.600 59.100 ;
        RECT 117.270 59.300 117.440 59.470 ;
        RECT 120.150 58.930 120.320 59.100 ;
        RECT 123.030 59.300 123.200 59.470 ;
        RECT 126.870 58.930 127.040 59.100 ;
        RECT 129.750 59.300 129.920 59.470 ;
        RECT 133.590 58.930 133.760 59.100 ;
        RECT 6.390 54.490 6.560 54.660 ;
      LAYER mcon ;
        RECT 5.880 53.310 6.050 53.480 ;
        RECT 6.240 53.310 6.410 53.480 ;
      LAYER L1M1_PR_C ;
        RECT 6.870 54.120 7.040 54.290 ;
        RECT 10.230 55.970 10.400 56.140 ;
        RECT 12.630 55.970 12.800 56.140 ;
        RECT 9.750 54.490 9.920 54.660 ;
      LAYER mcon ;
        RECT 7.420 53.310 7.590 53.480 ;
        RECT 7.860 53.310 8.030 53.480 ;
        RECT 8.300 53.310 8.470 53.480 ;
        RECT 8.710 53.310 8.880 53.480 ;
        RECT 9.240 53.310 9.410 53.480 ;
        RECT 9.600 53.310 9.770 53.480 ;
      LAYER L1M1_PR_C ;
        RECT 14.070 55.600 14.240 55.770 ;
      LAYER mcon ;
        RECT 10.780 53.310 10.950 53.480 ;
        RECT 11.220 53.310 11.390 53.480 ;
        RECT 11.660 53.310 11.830 53.480 ;
        RECT 12.070 53.310 12.240 53.480 ;
        RECT 13.030 53.310 13.200 53.480 ;
        RECT 13.390 53.310 13.560 53.480 ;
        RECT 13.750 53.310 13.920 53.480 ;
        RECT 14.110 53.310 14.280 53.480 ;
      LAYER L1M1_PR_C ;
        RECT 18.390 54.860 18.560 55.030 ;
        RECT 18.870 54.860 19.040 55.030 ;
        RECT 16.950 54.490 17.120 54.660 ;
      LAYER mcon ;
        RECT 15.100 53.310 15.270 53.480 ;
        RECT 15.540 53.310 15.710 53.480 ;
        RECT 15.980 53.310 16.150 53.480 ;
        RECT 16.390 53.310 16.560 53.480 ;
        RECT 16.920 53.310 17.090 53.480 ;
        RECT 17.280 53.310 17.450 53.480 ;
        RECT 18.190 53.310 18.360 53.480 ;
        RECT 18.550 53.310 18.720 53.480 ;
        RECT 18.910 53.310 19.080 53.480 ;
      LAYER L1M1_PR_C ;
        RECT 19.350 53.750 19.520 53.920 ;
        RECT 19.830 54.860 20.000 55.030 ;
        RECT 23.670 55.230 23.840 55.400 ;
        RECT 24.630 54.860 24.800 55.030 ;
        RECT 22.230 54.490 22.400 54.660 ;
        RECT 25.590 54.860 25.760 55.030 ;
        RECT 23.190 54.490 23.360 54.660 ;
      LAYER mcon ;
        RECT 20.380 53.310 20.550 53.480 ;
        RECT 20.820 53.310 20.990 53.480 ;
        RECT 21.260 53.310 21.430 53.480 ;
        RECT 21.670 53.310 21.840 53.480 ;
        RECT 24.280 53.310 24.450 53.480 ;
        RECT 24.640 53.310 24.810 53.480 ;
        RECT 25.000 53.310 25.170 53.480 ;
      LAYER L1M1_PR_C ;
        RECT 31.830 54.860 32.000 55.030 ;
      LAYER mcon ;
        RECT 26.140 53.310 26.310 53.480 ;
        RECT 26.580 53.310 26.750 53.480 ;
        RECT 27.020 53.310 27.190 53.480 ;
        RECT 27.430 53.310 27.600 53.480 ;
        RECT 27.960 53.310 28.130 53.480 ;
        RECT 28.320 53.310 28.490 53.480 ;
        RECT 28.680 53.310 28.850 53.480 ;
      LAYER L1M1_PR_C ;
        RECT 30.390 54.120 30.560 54.290 ;
      LAYER mcon ;
        RECT 29.520 53.310 29.690 53.480 ;
        RECT 29.880 53.310 30.050 53.480 ;
        RECT 30.240 53.310 30.410 53.480 ;
        RECT 31.080 53.310 31.250 53.480 ;
        RECT 31.440 53.310 31.610 53.480 ;
        RECT 31.800 53.310 31.970 53.480 ;
      LAYER L1M1_PR_C ;
        RECT 38.550 54.860 38.720 55.030 ;
        RECT 34.710 54.490 34.880 54.660 ;
      LAYER mcon ;
        RECT 32.860 53.310 33.030 53.480 ;
        RECT 33.300 53.310 33.470 53.480 ;
        RECT 33.740 53.310 33.910 53.480 ;
        RECT 34.150 53.310 34.320 53.480 ;
        RECT 34.680 53.310 34.850 53.480 ;
        RECT 35.040 53.310 35.210 53.480 ;
        RECT 35.400 53.310 35.570 53.480 ;
        RECT 36.240 53.310 36.410 53.480 ;
        RECT 36.600 53.310 36.770 53.480 ;
        RECT 36.960 53.310 37.130 53.480 ;
        RECT 37.800 53.310 37.970 53.480 ;
        RECT 38.160 53.310 38.330 53.480 ;
        RECT 38.520 53.310 38.690 53.480 ;
      LAYER L1M1_PR_C ;
        RECT 45.270 54.860 45.440 55.030 ;
      LAYER mcon ;
        RECT 39.580 53.310 39.750 53.480 ;
        RECT 40.020 53.310 40.190 53.480 ;
        RECT 40.460 53.310 40.630 53.480 ;
        RECT 40.870 53.310 41.040 53.480 ;
        RECT 41.400 53.310 41.570 53.480 ;
        RECT 41.760 53.310 41.930 53.480 ;
        RECT 42.120 53.310 42.290 53.480 ;
      LAYER L1M1_PR_C ;
        RECT 43.830 54.120 44.000 54.290 ;
      LAYER mcon ;
        RECT 42.960 53.310 43.130 53.480 ;
        RECT 43.320 53.310 43.490 53.480 ;
        RECT 43.680 53.310 43.850 53.480 ;
        RECT 44.520 53.310 44.690 53.480 ;
        RECT 44.880 53.310 45.050 53.480 ;
        RECT 45.240 53.310 45.410 53.480 ;
      LAYER L1M1_PR_C ;
        RECT 51.990 54.860 52.160 55.030 ;
        RECT 48.150 54.490 48.320 54.660 ;
      LAYER mcon ;
        RECT 46.300 53.310 46.470 53.480 ;
        RECT 46.740 53.310 46.910 53.480 ;
        RECT 47.180 53.310 47.350 53.480 ;
        RECT 47.590 53.310 47.760 53.480 ;
        RECT 48.120 53.310 48.290 53.480 ;
        RECT 48.480 53.310 48.650 53.480 ;
        RECT 48.840 53.310 49.010 53.480 ;
        RECT 49.680 53.310 49.850 53.480 ;
        RECT 50.040 53.310 50.210 53.480 ;
        RECT 50.400 53.310 50.570 53.480 ;
        RECT 51.240 53.310 51.410 53.480 ;
        RECT 51.600 53.310 51.770 53.480 ;
        RECT 51.960 53.310 52.130 53.480 ;
      LAYER L1M1_PR_C ;
        RECT 58.710 54.860 58.880 55.030 ;
      LAYER mcon ;
        RECT 53.020 53.310 53.190 53.480 ;
        RECT 53.460 53.310 53.630 53.480 ;
        RECT 53.900 53.310 54.070 53.480 ;
        RECT 54.310 53.310 54.480 53.480 ;
        RECT 54.840 53.310 55.010 53.480 ;
        RECT 55.200 53.310 55.370 53.480 ;
        RECT 55.560 53.310 55.730 53.480 ;
      LAYER L1M1_PR_C ;
        RECT 56.310 54.120 56.480 54.290 ;
      LAYER mcon ;
        RECT 56.400 53.310 56.570 53.480 ;
        RECT 56.760 53.310 56.930 53.480 ;
        RECT 57.120 53.310 57.290 53.480 ;
        RECT 57.960 53.310 58.130 53.480 ;
        RECT 58.320 53.310 58.490 53.480 ;
        RECT 58.680 53.310 58.850 53.480 ;
      LAYER L1M1_PR_C ;
        RECT 65.430 54.860 65.600 55.030 ;
        RECT 61.590 54.490 61.760 54.660 ;
      LAYER mcon ;
        RECT 59.740 53.310 59.910 53.480 ;
        RECT 60.180 53.310 60.350 53.480 ;
        RECT 60.620 53.310 60.790 53.480 ;
        RECT 61.030 53.310 61.200 53.480 ;
        RECT 61.560 53.310 61.730 53.480 ;
        RECT 61.920 53.310 62.090 53.480 ;
        RECT 62.280 53.310 62.450 53.480 ;
        RECT 63.120 53.310 63.290 53.480 ;
        RECT 63.480 53.310 63.650 53.480 ;
        RECT 63.840 53.310 64.010 53.480 ;
        RECT 64.680 53.310 64.850 53.480 ;
        RECT 65.040 53.310 65.210 53.480 ;
        RECT 65.400 53.310 65.570 53.480 ;
      LAYER L1M1_PR_C ;
        RECT 72.150 54.860 72.320 55.030 ;
        RECT 68.310 54.490 68.480 54.660 ;
      LAYER mcon ;
        RECT 66.460 53.310 66.630 53.480 ;
        RECT 66.900 53.310 67.070 53.480 ;
        RECT 67.340 53.310 67.510 53.480 ;
        RECT 67.750 53.310 67.920 53.480 ;
        RECT 68.280 53.310 68.450 53.480 ;
        RECT 68.640 53.310 68.810 53.480 ;
        RECT 69.000 53.310 69.170 53.480 ;
        RECT 69.840 53.310 70.010 53.480 ;
        RECT 70.200 53.310 70.370 53.480 ;
        RECT 70.560 53.310 70.730 53.480 ;
        RECT 71.400 53.310 71.570 53.480 ;
        RECT 71.760 53.310 71.930 53.480 ;
        RECT 72.120 53.310 72.290 53.480 ;
      LAYER L1M1_PR_C ;
        RECT 78.870 54.860 79.040 55.030 ;
        RECT 75.030 54.490 75.200 54.660 ;
      LAYER mcon ;
        RECT 73.180 53.310 73.350 53.480 ;
        RECT 73.620 53.310 73.790 53.480 ;
        RECT 74.060 53.310 74.230 53.480 ;
        RECT 74.470 53.310 74.640 53.480 ;
        RECT 75.000 53.310 75.170 53.480 ;
        RECT 75.360 53.310 75.530 53.480 ;
        RECT 75.720 53.310 75.890 53.480 ;
        RECT 76.560 53.310 76.730 53.480 ;
        RECT 76.920 53.310 77.090 53.480 ;
        RECT 77.280 53.310 77.450 53.480 ;
        RECT 78.120 53.310 78.290 53.480 ;
        RECT 78.480 53.310 78.650 53.480 ;
        RECT 78.840 53.310 79.010 53.480 ;
      LAYER L1M1_PR_C ;
        RECT 86.550 54.860 86.720 55.030 ;
        RECT 82.710 54.490 82.880 54.660 ;
      LAYER mcon ;
        RECT 79.900 53.310 80.070 53.480 ;
        RECT 80.340 53.310 80.510 53.480 ;
        RECT 80.780 53.310 80.950 53.480 ;
        RECT 81.190 53.310 81.360 53.480 ;
        RECT 82.680 53.310 82.850 53.480 ;
        RECT 83.040 53.310 83.210 53.480 ;
        RECT 83.400 53.310 83.570 53.480 ;
        RECT 84.240 53.310 84.410 53.480 ;
        RECT 84.600 53.310 84.770 53.480 ;
        RECT 84.960 53.310 85.130 53.480 ;
        RECT 85.800 53.310 85.970 53.480 ;
        RECT 86.160 53.310 86.330 53.480 ;
        RECT 86.520 53.310 86.690 53.480 ;
      LAYER L1M1_PR_C ;
        RECT 90.870 55.970 91.040 56.140 ;
        RECT 91.830 54.860 92.000 55.030 ;
        RECT 89.430 54.490 89.600 54.660 ;
        RECT 90.390 54.490 90.560 54.660 ;
      LAYER mcon ;
        RECT 87.580 53.310 87.750 53.480 ;
        RECT 88.020 53.310 88.190 53.480 ;
        RECT 88.460 53.310 88.630 53.480 ;
        RECT 88.870 53.310 89.040 53.480 ;
        RECT 91.480 53.310 91.650 53.480 ;
        RECT 91.840 53.310 92.010 53.480 ;
        RECT 92.200 53.310 92.370 53.480 ;
      LAYER L1M1_PR_C ;
        RECT 96.150 55.970 96.320 56.140 ;
        RECT 95.190 54.490 95.360 54.660 ;
      LAYER mcon ;
        RECT 93.340 53.310 93.510 53.480 ;
        RECT 93.780 53.310 93.950 53.480 ;
        RECT 94.220 53.310 94.390 53.480 ;
        RECT 94.630 53.310 94.800 53.480 ;
      LAYER L1M1_PR_C ;
        RECT 96.630 54.490 96.800 54.660 ;
        RECT 97.110 54.490 97.280 54.660 ;
        RECT 98.070 54.490 98.240 54.660 ;
      LAYER mcon ;
        RECT 95.160 53.310 95.330 53.480 ;
        RECT 95.520 53.310 95.690 53.480 ;
      LAYER L1M1_PR_C ;
        RECT 106.230 54.860 106.400 55.030 ;
      LAYER mcon ;
        RECT 97.180 53.310 97.350 53.480 ;
        RECT 97.540 53.310 97.710 53.480 ;
        RECT 97.900 53.310 98.070 53.480 ;
        RECT 98.260 53.310 98.430 53.480 ;
        RECT 98.620 53.310 98.790 53.480 ;
        RECT 99.100 53.310 99.270 53.480 ;
        RECT 99.540 53.310 99.710 53.480 ;
        RECT 99.980 53.310 100.150 53.480 ;
        RECT 100.390 53.310 100.560 53.480 ;
        RECT 102.360 53.310 102.530 53.480 ;
        RECT 102.720 53.310 102.890 53.480 ;
        RECT 103.080 53.310 103.250 53.480 ;
      LAYER L1M1_PR_C ;
        RECT 104.790 54.120 104.960 54.290 ;
      LAYER mcon ;
        RECT 103.920 53.310 104.090 53.480 ;
        RECT 104.280 53.310 104.450 53.480 ;
        RECT 104.640 53.310 104.810 53.480 ;
        RECT 105.480 53.310 105.650 53.480 ;
        RECT 105.840 53.310 106.010 53.480 ;
        RECT 106.200 53.310 106.370 53.480 ;
      LAYER L1M1_PR_C ;
        RECT 112.950 54.860 113.120 55.030 ;
        RECT 110.070 54.490 110.240 54.660 ;
      LAYER mcon ;
        RECT 107.260 53.310 107.430 53.480 ;
        RECT 107.700 53.310 107.870 53.480 ;
        RECT 108.140 53.310 108.310 53.480 ;
        RECT 108.550 53.310 108.720 53.480 ;
        RECT 109.080 53.310 109.250 53.480 ;
        RECT 109.440 53.310 109.610 53.480 ;
        RECT 109.800 53.310 109.970 53.480 ;
        RECT 110.640 53.310 110.810 53.480 ;
        RECT 111.000 53.310 111.170 53.480 ;
        RECT 111.360 53.310 111.530 53.480 ;
        RECT 112.200 53.310 112.370 53.480 ;
        RECT 112.560 53.310 112.730 53.480 ;
        RECT 112.920 53.310 113.090 53.480 ;
      LAYER L1M1_PR_C ;
        RECT 120.150 54.860 120.320 55.030 ;
      LAYER mcon ;
        RECT 113.980 53.310 114.150 53.480 ;
        RECT 114.420 53.310 114.590 53.480 ;
        RECT 114.860 53.310 115.030 53.480 ;
        RECT 115.270 53.310 115.440 53.480 ;
        RECT 116.280 53.310 116.450 53.480 ;
        RECT 116.640 53.310 116.810 53.480 ;
        RECT 117.000 53.310 117.170 53.480 ;
      LAYER L1M1_PR_C ;
        RECT 118.230 54.120 118.400 54.290 ;
      LAYER mcon ;
        RECT 117.840 53.310 118.010 53.480 ;
        RECT 118.200 53.310 118.370 53.480 ;
        RECT 118.560 53.310 118.730 53.480 ;
        RECT 119.400 53.310 119.570 53.480 ;
        RECT 119.760 53.310 119.930 53.480 ;
        RECT 120.120 53.310 120.290 53.480 ;
      LAYER L1M1_PR_C ;
        RECT 126.870 54.860 127.040 55.030 ;
        RECT 123.030 54.490 123.200 54.660 ;
      LAYER mcon ;
        RECT 121.180 53.310 121.350 53.480 ;
        RECT 121.620 53.310 121.790 53.480 ;
        RECT 122.060 53.310 122.230 53.480 ;
        RECT 122.470 53.310 122.640 53.480 ;
        RECT 123.000 53.310 123.170 53.480 ;
        RECT 123.360 53.310 123.530 53.480 ;
        RECT 123.720 53.310 123.890 53.480 ;
        RECT 124.560 53.310 124.730 53.480 ;
        RECT 124.920 53.310 125.090 53.480 ;
        RECT 125.280 53.310 125.450 53.480 ;
        RECT 126.120 53.310 126.290 53.480 ;
        RECT 126.480 53.310 126.650 53.480 ;
        RECT 126.840 53.310 127.010 53.480 ;
      LAYER L1M1_PR_C ;
        RECT 133.590 54.860 133.760 55.030 ;
        RECT 130.230 54.490 130.400 54.660 ;
      LAYER mcon ;
        RECT 127.900 53.310 128.070 53.480 ;
        RECT 128.340 53.310 128.510 53.480 ;
        RECT 128.780 53.310 128.950 53.480 ;
        RECT 129.190 53.310 129.360 53.480 ;
        RECT 129.720 53.310 129.890 53.480 ;
        RECT 130.080 53.310 130.250 53.480 ;
        RECT 130.440 53.310 130.610 53.480 ;
        RECT 131.280 53.310 131.450 53.480 ;
        RECT 131.640 53.310 131.810 53.480 ;
        RECT 132.000 53.310 132.170 53.480 ;
        RECT 132.840 53.310 133.010 53.480 ;
        RECT 133.200 53.310 133.370 53.480 ;
        RECT 133.560 53.310 133.730 53.480 ;
      LAYER L1M1_PR_C ;
        RECT 137.910 55.970 138.080 56.140 ;
        RECT 138.870 54.860 139.040 55.030 ;
        RECT 136.470 54.490 136.640 54.660 ;
        RECT 139.350 54.860 139.520 55.030 ;
        RECT 137.430 54.490 137.600 54.660 ;
      LAYER mcon ;
        RECT 134.620 53.310 134.790 53.480 ;
        RECT 135.060 53.310 135.230 53.480 ;
        RECT 135.500 53.310 135.670 53.480 ;
        RECT 135.910 53.310 136.080 53.480 ;
        RECT 138.520 53.310 138.690 53.480 ;
        RECT 138.880 53.310 139.050 53.480 ;
        RECT 139.240 53.310 139.410 53.480 ;
        RECT 140.380 53.310 140.550 53.480 ;
        RECT 140.820 53.310 140.990 53.480 ;
        RECT 141.260 53.310 141.430 53.480 ;
        RECT 141.670 53.310 141.840 53.480 ;
      LAYER L1M1_PR_C ;
        RECT 13.110 51.160 13.280 51.330 ;
        RECT 11.670 50.420 11.840 50.590 ;
        RECT 9.270 50.050 9.440 50.220 ;
        RECT 17.430 51.530 17.600 51.700 ;
        RECT 16.470 51.160 16.640 51.330 ;
        RECT 17.910 51.160 18.080 51.330 ;
        RECT 20.790 51.160 20.960 51.330 ;
        RECT 21.750 51.160 21.920 51.330 ;
        RECT 22.710 51.160 22.880 51.330 ;
        RECT 23.670 51.160 23.840 51.330 ;
        RECT 21.270 50.790 21.440 50.960 ;
        RECT 26.070 51.530 26.240 51.700 ;
        RECT 27.030 50.790 27.200 50.960 ;
        RECT 29.910 51.160 30.080 51.330 ;
        RECT 32.310 51.160 32.480 51.330 ;
        RECT 36.150 50.790 36.320 50.960 ;
        RECT 39.030 51.160 39.200 51.330 ;
        RECT 42.870 50.790 43.040 50.960 ;
        RECT 50.070 51.530 50.240 51.700 ;
        RECT 51.990 50.790 52.160 50.960 ;
        RECT 60.150 51.530 60.320 51.700 ;
        RECT 61.590 50.790 61.760 50.960 ;
        RECT 64.470 51.160 64.640 51.330 ;
        RECT 68.310 50.790 68.480 50.960 ;
        RECT 72.630 51.530 72.800 51.700 ;
        RECT 75.030 50.790 75.200 50.960 ;
        RECT 78.870 51.530 79.040 51.700 ;
        RECT 77.910 51.160 78.080 51.330 ;
        RECT 84.150 51.530 84.320 51.700 ;
        RECT 85.590 50.790 85.760 50.960 ;
        RECT 88.470 51.160 88.640 51.330 ;
        RECT 92.310 50.790 92.480 50.960 ;
        RECT 95.670 51.160 95.840 51.330 ;
        RECT 99.510 51.160 99.680 51.330 ;
        RECT 96.150 49.680 96.320 49.850 ;
        RECT 102.390 50.790 102.560 50.960 ;
        RECT 108.630 51.160 108.800 51.330 ;
        RECT 111.510 50.790 111.680 50.960 ;
        RECT 116.310 51.530 116.480 51.700 ;
        RECT 118.230 50.790 118.400 50.960 ;
        RECT 124.950 51.160 125.120 51.330 ;
        RECT 128.310 51.160 128.480 51.330 ;
        RECT 126.390 50.790 126.560 50.960 ;
        RECT 133.110 51.530 133.280 51.700 ;
        RECT 134.550 50.790 134.720 50.960 ;
        RECT 139.350 51.160 139.520 51.330 ;
        RECT 137.430 50.790 137.600 50.960 ;
        RECT 138.870 50.790 139.040 50.960 ;
      LAYER mcon ;
        RECT 6.510 45.160 6.680 45.330 ;
        RECT 6.950 45.160 7.120 45.330 ;
        RECT 7.360 45.160 7.530 45.330 ;
        RECT 7.790 45.160 7.960 45.330 ;
        RECT 8.230 45.160 8.400 45.330 ;
        RECT 8.640 45.160 8.810 45.330 ;
      LAYER L1M1_PR_C ;
        RECT 12.630 47.090 12.800 47.260 ;
      LAYER mcon ;
        RECT 10.190 45.170 10.360 45.340 ;
        RECT 10.550 45.170 10.720 45.340 ;
        RECT 10.910 45.170 11.080 45.340 ;
        RECT 11.830 45.170 12.000 45.340 ;
        RECT 12.190 45.170 12.360 45.340 ;
      LAYER L1M1_PR_C ;
        RECT 13.110 45.980 13.280 46.150 ;
      LAYER mcon ;
        RECT 16.790 45.170 16.960 45.340 ;
        RECT 17.150 45.170 17.320 45.340 ;
        RECT 17.510 45.170 17.680 45.340 ;
      LAYER L1M1_PR_C ;
        RECT 24.630 46.720 24.800 46.890 ;
      LAYER mcon ;
        RECT 20.760 45.170 20.930 45.340 ;
        RECT 21.120 45.170 21.290 45.340 ;
        RECT 21.480 45.170 21.650 45.340 ;
      LAYER L1M1_PR_C ;
        RECT 28.470 46.720 28.640 46.890 ;
      LAYER mcon ;
        RECT 23.370 45.170 23.540 45.340 ;
        RECT 23.730 45.170 23.900 45.340 ;
        RECT 24.090 45.170 24.260 45.340 ;
        RECT 25.180 45.170 25.350 45.340 ;
        RECT 25.620 45.170 25.790 45.340 ;
        RECT 26.060 45.170 26.230 45.340 ;
        RECT 26.470 45.170 26.640 45.340 ;
      LAYER L1M1_PR_C ;
        RECT 27.030 45.980 27.200 46.150 ;
        RECT 29.430 46.720 29.600 46.890 ;
        RECT 29.910 46.350 30.080 46.520 ;
        RECT 30.870 46.350 31.040 46.520 ;
        RECT 36.150 47.460 36.320 47.630 ;
        RECT 35.670 46.720 35.840 46.890 ;
        RECT 36.630 47.830 36.800 48.000 ;
        RECT 34.230 46.350 34.400 46.520 ;
      LAYER mcon ;
        RECT 27.440 45.170 27.610 45.340 ;
        RECT 27.800 45.170 27.970 45.340 ;
        RECT 28.160 45.170 28.330 45.340 ;
        RECT 30.800 45.170 30.970 45.340 ;
        RECT 31.160 45.170 31.330 45.340 ;
        RECT 31.520 45.170 31.690 45.340 ;
        RECT 31.880 45.170 32.050 45.340 ;
        RECT 32.380 45.170 32.550 45.340 ;
        RECT 32.820 45.170 32.990 45.340 ;
        RECT 33.260 45.170 33.430 45.340 ;
        RECT 33.670 45.170 33.840 45.340 ;
        RECT 34.200 45.170 34.370 45.340 ;
        RECT 34.560 45.170 34.730 45.340 ;
        RECT 35.470 45.170 35.640 45.340 ;
        RECT 35.830 45.170 36.000 45.340 ;
        RECT 36.190 45.170 36.360 45.340 ;
      LAYER L1M1_PR_C ;
        RECT 43.350 46.720 43.520 46.890 ;
      LAYER mcon ;
        RECT 37.660 45.170 37.830 45.340 ;
        RECT 38.100 45.170 38.270 45.340 ;
        RECT 38.540 45.170 38.710 45.340 ;
        RECT 38.950 45.170 39.120 45.340 ;
        RECT 39.480 45.170 39.650 45.340 ;
        RECT 39.840 45.170 40.010 45.340 ;
        RECT 40.200 45.170 40.370 45.340 ;
      LAYER L1M1_PR_C ;
        RECT 41.910 45.980 42.080 46.150 ;
      LAYER mcon ;
        RECT 41.040 45.170 41.210 45.340 ;
        RECT 41.400 45.170 41.570 45.340 ;
        RECT 41.760 45.170 41.930 45.340 ;
        RECT 42.600 45.170 42.770 45.340 ;
        RECT 42.960 45.170 43.130 45.340 ;
        RECT 43.320 45.170 43.490 45.340 ;
      LAYER L1M1_PR_C ;
        RECT 46.710 46.350 46.880 46.520 ;
        RECT 48.150 46.350 48.320 46.520 ;
      LAYER mcon ;
        RECT 44.380 45.170 44.550 45.340 ;
        RECT 44.820 45.170 44.990 45.340 ;
        RECT 45.260 45.170 45.430 45.340 ;
        RECT 45.670 45.170 45.840 45.340 ;
        RECT 46.200 45.170 46.370 45.340 ;
        RECT 46.560 45.170 46.730 45.340 ;
        RECT 46.920 45.170 47.090 45.340 ;
        RECT 47.280 45.170 47.450 45.340 ;
      LAYER L1M1_PR_C ;
        RECT 54.870 46.720 55.040 46.890 ;
        RECT 48.150 45.610 48.320 45.780 ;
      LAYER mcon ;
        RECT 48.700 45.170 48.870 45.340 ;
        RECT 49.140 45.170 49.310 45.340 ;
        RECT 49.580 45.170 49.750 45.340 ;
        RECT 49.990 45.170 50.160 45.340 ;
        RECT 51.000 45.170 51.170 45.340 ;
        RECT 51.360 45.170 51.530 45.340 ;
        RECT 51.720 45.170 51.890 45.340 ;
      LAYER L1M1_PR_C ;
        RECT 53.430 45.980 53.600 46.150 ;
      LAYER mcon ;
        RECT 52.560 45.170 52.730 45.340 ;
        RECT 52.920 45.170 53.090 45.340 ;
        RECT 53.280 45.170 53.450 45.340 ;
        RECT 54.120 45.170 54.290 45.340 ;
        RECT 54.480 45.170 54.650 45.340 ;
        RECT 54.840 45.170 55.010 45.340 ;
      LAYER L1M1_PR_C ;
        RECT 61.590 46.720 61.760 46.890 ;
      LAYER mcon ;
        RECT 55.900 45.170 56.070 45.340 ;
        RECT 56.340 45.170 56.510 45.340 ;
        RECT 56.780 45.170 56.950 45.340 ;
        RECT 57.190 45.170 57.360 45.340 ;
        RECT 57.720 45.170 57.890 45.340 ;
        RECT 58.080 45.170 58.250 45.340 ;
        RECT 58.440 45.170 58.610 45.340 ;
      LAYER L1M1_PR_C ;
        RECT 59.190 45.980 59.360 46.150 ;
      LAYER mcon ;
        RECT 59.280 45.170 59.450 45.340 ;
        RECT 59.640 45.170 59.810 45.340 ;
        RECT 60.000 45.170 60.170 45.340 ;
        RECT 60.840 45.170 61.010 45.340 ;
        RECT 61.200 45.170 61.370 45.340 ;
        RECT 61.560 45.170 61.730 45.340 ;
      LAYER L1M1_PR_C ;
        RECT 65.430 46.720 65.600 46.890 ;
        RECT 65.910 46.720 66.080 46.890 ;
        RECT 66.390 46.350 66.560 46.520 ;
      LAYER mcon ;
        RECT 62.620 45.170 62.790 45.340 ;
        RECT 63.060 45.170 63.230 45.340 ;
        RECT 63.500 45.170 63.670 45.340 ;
        RECT 63.910 45.170 64.080 45.340 ;
        RECT 64.430 45.170 64.600 45.340 ;
        RECT 64.790 45.170 64.960 45.340 ;
        RECT 65.150 45.170 65.320 45.340 ;
        RECT 66.070 45.170 66.240 45.340 ;
        RECT 66.430 45.170 66.600 45.340 ;
        RECT 66.940 45.170 67.110 45.340 ;
        RECT 67.380 45.170 67.550 45.340 ;
        RECT 67.820 45.170 67.990 45.340 ;
        RECT 68.230 45.170 68.400 45.340 ;
      LAYER L1M1_PR_C ;
        RECT 71.670 47.090 71.840 47.260 ;
      LAYER mcon ;
        RECT 69.230 45.170 69.400 45.340 ;
        RECT 69.590 45.170 69.760 45.340 ;
        RECT 69.950 45.170 70.120 45.340 ;
        RECT 70.870 45.170 71.040 45.340 ;
        RECT 71.230 45.170 71.400 45.340 ;
      LAYER L1M1_PR_C ;
        RECT 72.150 45.610 72.320 45.780 ;
      LAYER mcon ;
        RECT 75.830 45.170 76.000 45.340 ;
        RECT 76.190 45.170 76.360 45.340 ;
        RECT 76.550 45.170 76.720 45.340 ;
        RECT 79.800 45.170 79.970 45.340 ;
        RECT 80.160 45.170 80.330 45.340 ;
        RECT 80.520 45.170 80.690 45.340 ;
      LAYER L1M1_PR_C ;
        RECT 83.670 45.610 83.840 45.780 ;
        RECT 89.910 46.720 90.080 46.890 ;
      LAYER mcon ;
        RECT 82.410 45.170 82.580 45.340 ;
        RECT 82.770 45.170 82.940 45.340 ;
        RECT 83.130 45.170 83.300 45.340 ;
        RECT 84.220 45.170 84.390 45.340 ;
        RECT 84.660 45.170 84.830 45.340 ;
        RECT 85.100 45.170 85.270 45.340 ;
        RECT 85.510 45.170 85.680 45.340 ;
        RECT 86.040 45.170 86.210 45.340 ;
        RECT 86.400 45.170 86.570 45.340 ;
        RECT 86.760 45.170 86.930 45.340 ;
      LAYER L1M1_PR_C ;
        RECT 88.470 45.980 88.640 46.150 ;
      LAYER mcon ;
        RECT 87.600 45.170 87.770 45.340 ;
        RECT 87.960 45.170 88.130 45.340 ;
        RECT 88.320 45.170 88.490 45.340 ;
        RECT 89.160 45.170 89.330 45.340 ;
        RECT 89.520 45.170 89.690 45.340 ;
        RECT 89.880 45.170 90.050 45.340 ;
        RECT 91.470 45.160 91.640 45.330 ;
        RECT 91.910 45.160 92.080 45.330 ;
        RECT 92.320 45.160 92.490 45.330 ;
        RECT 92.750 45.160 92.920 45.330 ;
        RECT 93.190 45.160 93.360 45.330 ;
        RECT 93.600 45.160 93.770 45.330 ;
      LAYER L1M1_PR_C ;
        RECT 96.630 46.720 96.800 46.890 ;
        RECT 95.190 45.610 95.360 45.780 ;
        RECT 97.590 46.720 97.760 46.890 ;
        RECT 98.070 46.350 98.240 46.520 ;
        RECT 98.550 46.350 98.720 46.520 ;
        RECT 104.790 46.720 104.960 46.890 ;
        RECT 102.390 46.350 102.560 46.520 ;
        RECT 105.270 46.720 105.440 46.890 ;
        RECT 103.350 46.350 103.520 46.520 ;
      LAYER mcon ;
        RECT 95.600 45.170 95.770 45.340 ;
        RECT 95.960 45.170 96.130 45.340 ;
        RECT 96.320 45.170 96.490 45.340 ;
        RECT 98.960 45.170 99.130 45.340 ;
        RECT 99.320 45.170 99.490 45.340 ;
        RECT 99.680 45.170 99.850 45.340 ;
        RECT 100.040 45.170 100.210 45.340 ;
        RECT 100.540 45.170 100.710 45.340 ;
        RECT 100.980 45.170 101.150 45.340 ;
        RECT 101.420 45.170 101.590 45.340 ;
        RECT 101.830 45.170 102.000 45.340 ;
      LAYER L1M1_PR_C ;
        RECT 103.350 45.610 103.520 45.780 ;
      LAYER mcon ;
        RECT 104.440 45.170 104.610 45.340 ;
        RECT 104.800 45.170 104.970 45.340 ;
        RECT 105.160 45.170 105.330 45.340 ;
      LAYER L1M1_PR_C ;
        RECT 112.470 46.720 112.640 46.890 ;
        RECT 108.630 46.350 108.800 46.520 ;
      LAYER mcon ;
        RECT 106.300 45.170 106.470 45.340 ;
        RECT 106.740 45.170 106.910 45.340 ;
        RECT 107.180 45.170 107.350 45.340 ;
        RECT 107.590 45.170 107.760 45.340 ;
        RECT 108.600 45.170 108.770 45.340 ;
        RECT 108.960 45.170 109.130 45.340 ;
        RECT 109.320 45.170 109.490 45.340 ;
        RECT 110.160 45.170 110.330 45.340 ;
        RECT 110.520 45.170 110.690 45.340 ;
        RECT 110.880 45.170 111.050 45.340 ;
        RECT 111.720 45.170 111.890 45.340 ;
        RECT 112.080 45.170 112.250 45.340 ;
        RECT 112.440 45.170 112.610 45.340 ;
      LAYER L1M1_PR_C ;
        RECT 120.150 46.720 120.320 46.890 ;
      LAYER mcon ;
        RECT 113.500 45.170 113.670 45.340 ;
        RECT 113.940 45.170 114.110 45.340 ;
        RECT 114.380 45.170 114.550 45.340 ;
        RECT 114.790 45.170 114.960 45.340 ;
        RECT 116.280 45.170 116.450 45.340 ;
        RECT 116.640 45.170 116.810 45.340 ;
        RECT 117.000 45.170 117.170 45.340 ;
      LAYER L1M1_PR_C ;
        RECT 117.750 45.980 117.920 46.150 ;
      LAYER mcon ;
        RECT 117.840 45.170 118.010 45.340 ;
        RECT 118.200 45.170 118.370 45.340 ;
        RECT 118.560 45.170 118.730 45.340 ;
        RECT 119.400 45.170 119.570 45.340 ;
        RECT 119.760 45.170 119.930 45.340 ;
        RECT 120.120 45.170 120.290 45.340 ;
        RECT 121.710 45.160 121.880 45.330 ;
        RECT 122.150 45.160 122.320 45.330 ;
        RECT 122.560 45.160 122.730 45.330 ;
        RECT 122.990 45.160 123.160 45.330 ;
        RECT 123.430 45.160 123.600 45.330 ;
        RECT 123.840 45.160 124.010 45.330 ;
        RECT 125.390 45.170 125.560 45.340 ;
        RECT 125.750 45.170 125.920 45.340 ;
        RECT 126.110 45.170 126.280 45.340 ;
        RECT 127.030 45.170 127.200 45.340 ;
        RECT 127.390 45.170 127.560 45.340 ;
      LAYER L1M1_PR_C ;
        RECT 128.310 46.350 128.480 46.520 ;
      LAYER mcon ;
        RECT 131.990 45.170 132.160 45.340 ;
        RECT 132.350 45.170 132.520 45.340 ;
        RECT 132.710 45.170 132.880 45.340 ;
      LAYER L1M1_PR_C ;
        RECT 136.470 45.980 136.640 46.150 ;
      LAYER mcon ;
        RECT 135.960 45.170 136.130 45.340 ;
        RECT 136.320 45.170 136.490 45.340 ;
        RECT 136.680 45.170 136.850 45.340 ;
      LAYER L1M1_PR_C ;
        RECT 139.830 45.610 140.000 45.780 ;
      LAYER mcon ;
        RECT 138.570 45.170 138.740 45.340 ;
        RECT 138.930 45.170 139.100 45.340 ;
        RECT 139.290 45.170 139.460 45.340 ;
        RECT 140.380 45.170 140.550 45.340 ;
        RECT 140.820 45.170 140.990 45.340 ;
        RECT 141.260 45.170 141.430 45.340 ;
        RECT 141.670 45.170 141.840 45.340 ;
      LAYER L1M1_PR_C ;
        RECT 13.110 43.020 13.280 43.190 ;
        RECT 15.990 43.760 16.160 43.930 ;
        RECT 13.590 41.910 13.760 42.080 ;
        RECT 20.310 43.020 20.480 43.190 ;
        RECT 21.270 43.020 21.440 43.190 ;
        RECT 17.430 41.540 17.600 41.710 ;
        RECT 23.190 42.650 23.360 42.820 ;
        RECT 21.750 42.280 21.920 42.450 ;
        RECT 25.590 43.020 25.760 43.190 ;
        RECT 27.030 43.020 27.200 43.190 ;
        RECT 28.470 42.650 28.640 42.820 ;
        RECT 27.030 41.540 27.200 41.710 ;
        RECT 30.870 43.020 31.040 43.190 ;
        RECT 34.710 42.650 34.880 42.820 ;
        RECT 38.070 43.020 38.240 43.190 ;
        RECT 40.950 43.020 41.120 43.190 ;
        RECT 38.550 41.540 38.720 41.710 ;
        RECT 44.790 42.650 44.960 42.820 ;
        RECT 50.070 43.390 50.240 43.560 ;
        RECT 51.510 42.650 51.680 42.820 ;
        RECT 54.390 43.020 54.560 43.190 ;
        RECT 58.230 42.650 58.400 42.820 ;
        RECT 61.110 43.020 61.280 43.190 ;
        RECT 64.950 42.650 65.120 42.820 ;
        RECT 67.830 43.020 68.000 43.190 ;
        RECT 71.670 42.650 71.840 42.820 ;
        RECT 75.510 43.020 75.680 43.190 ;
        RECT 78.390 42.650 78.560 42.820 ;
        RECT 82.230 43.020 82.400 43.190 ;
        RECT 85.110 42.650 85.280 42.820 ;
        RECT 87.990 43.020 88.160 43.190 ;
        RECT 91.830 42.650 92.000 42.820 ;
        RECT 94.710 43.020 94.880 43.190 ;
        RECT 95.670 43.020 95.840 43.190 ;
        RECT 97.110 42.650 97.280 42.820 ;
        RECT 98.070 42.650 98.240 42.820 ;
        RECT 96.150 42.280 96.320 42.450 ;
        RECT 102.390 43.020 102.560 43.190 ;
        RECT 100.470 42.280 100.640 42.450 ;
        RECT 105.270 42.650 105.440 42.820 ;
        RECT 110.550 43.390 110.720 43.560 ;
        RECT 111.990 42.650 112.160 42.820 ;
        RECT 117.270 43.020 117.440 43.190 ;
        RECT 120.150 42.650 120.320 42.820 ;
        RECT 123.990 43.020 124.160 43.190 ;
        RECT 126.870 42.650 127.040 42.820 ;
        RECT 129.750 43.020 129.920 43.190 ;
        RECT 133.590 42.650 133.760 42.820 ;
        RECT 136.470 43.020 136.640 43.190 ;
        RECT 137.910 43.020 138.080 43.190 ;
        RECT 139.350 43.020 139.520 43.190 ;
        RECT 138.870 41.540 139.040 41.710 ;
        RECT 15.990 39.690 16.160 39.860 ;
        RECT 15.510 38.210 15.680 38.380 ;
      LAYER mcon ;
        RECT 6.510 37.020 6.680 37.190 ;
        RECT 6.950 37.020 7.120 37.190 ;
        RECT 7.360 37.020 7.530 37.190 ;
        RECT 7.790 37.020 7.960 37.190 ;
        RECT 8.230 37.020 8.400 37.190 ;
        RECT 8.640 37.020 8.810 37.190 ;
        RECT 10.350 37.020 10.520 37.190 ;
        RECT 10.790 37.020 10.960 37.190 ;
        RECT 11.200 37.020 11.370 37.190 ;
        RECT 11.630 37.020 11.800 37.190 ;
        RECT 12.070 37.020 12.240 37.190 ;
        RECT 12.480 37.020 12.650 37.190 ;
        RECT 15.000 37.030 15.170 37.200 ;
        RECT 15.360 37.030 15.530 37.200 ;
      LAYER L1M1_PR_C ;
        RECT 18.870 38.580 19.040 38.750 ;
        RECT 19.830 38.580 20.000 38.750 ;
        RECT 20.310 38.580 20.480 38.750 ;
      LAYER mcon ;
        RECT 16.540 37.030 16.710 37.200 ;
        RECT 16.980 37.030 17.150 37.200 ;
        RECT 17.420 37.030 17.590 37.200 ;
        RECT 17.830 37.030 18.000 37.200 ;
        RECT 18.350 37.030 18.520 37.200 ;
        RECT 18.710 37.030 18.880 37.200 ;
        RECT 19.070 37.030 19.240 37.200 ;
      LAYER L1M1_PR_C ;
        RECT 24.630 39.690 24.800 39.860 ;
        RECT 23.670 38.580 23.840 38.750 ;
        RECT 24.150 38.580 24.320 38.750 ;
      LAYER mcon ;
        RECT 19.990 37.030 20.160 37.200 ;
        RECT 20.350 37.030 20.520 37.200 ;
        RECT 20.860 37.030 21.030 37.200 ;
        RECT 21.300 37.030 21.470 37.200 ;
        RECT 21.740 37.030 21.910 37.200 ;
        RECT 22.150 37.030 22.320 37.200 ;
        RECT 22.670 37.030 22.840 37.200 ;
        RECT 23.030 37.030 23.200 37.200 ;
        RECT 23.390 37.030 23.560 37.200 ;
      LAYER L1M1_PR_C ;
        RECT 28.470 38.580 28.640 38.750 ;
        RECT 28.950 38.580 29.120 38.750 ;
        RECT 27.030 38.210 27.200 38.380 ;
      LAYER mcon ;
        RECT 24.310 37.030 24.480 37.200 ;
        RECT 24.670 37.030 24.840 37.200 ;
        RECT 25.180 37.030 25.350 37.200 ;
        RECT 25.620 37.030 25.790 37.200 ;
        RECT 26.060 37.030 26.230 37.200 ;
        RECT 26.470 37.030 26.640 37.200 ;
        RECT 27.000 37.030 27.170 37.200 ;
        RECT 27.360 37.030 27.530 37.200 ;
        RECT 28.270 37.030 28.440 37.200 ;
        RECT 28.630 37.030 28.800 37.200 ;
        RECT 28.990 37.030 29.160 37.200 ;
      LAYER L1M1_PR_C ;
        RECT 29.430 37.470 29.600 37.640 ;
        RECT 34.230 39.690 34.400 39.860 ;
        RECT 33.270 38.580 33.440 38.750 ;
        RECT 34.710 38.950 34.880 39.120 ;
        RECT 32.310 38.210 32.480 38.380 ;
      LAYER mcon ;
        RECT 30.460 37.030 30.630 37.200 ;
        RECT 30.900 37.030 31.070 37.200 ;
        RECT 31.340 37.030 31.510 37.200 ;
        RECT 31.750 37.030 31.920 37.200 ;
        RECT 32.280 37.030 32.450 37.200 ;
        RECT 32.640 37.030 32.810 37.200 ;
        RECT 33.550 37.030 33.720 37.200 ;
        RECT 33.910 37.030 34.080 37.200 ;
        RECT 34.270 37.030 34.440 37.200 ;
      LAYER L1M1_PR_C ;
        RECT 41.430 38.580 41.600 38.750 ;
      LAYER mcon ;
        RECT 35.740 37.030 35.910 37.200 ;
        RECT 36.180 37.030 36.350 37.200 ;
        RECT 36.620 37.030 36.790 37.200 ;
        RECT 37.030 37.030 37.200 37.200 ;
        RECT 37.560 37.030 37.730 37.200 ;
        RECT 37.920 37.030 38.090 37.200 ;
        RECT 38.280 37.030 38.450 37.200 ;
      LAYER L1M1_PR_C ;
        RECT 39.990 37.840 40.160 38.010 ;
      LAYER mcon ;
        RECT 39.120 37.030 39.290 37.200 ;
        RECT 39.480 37.030 39.650 37.200 ;
        RECT 39.840 37.030 40.010 37.200 ;
        RECT 40.680 37.030 40.850 37.200 ;
        RECT 41.040 37.030 41.210 37.200 ;
        RECT 41.400 37.030 41.570 37.200 ;
      LAYER L1M1_PR_C ;
        RECT 48.150 38.580 48.320 38.750 ;
        RECT 44.790 38.210 44.960 38.380 ;
      LAYER mcon ;
        RECT 42.460 37.030 42.630 37.200 ;
        RECT 42.900 37.030 43.070 37.200 ;
        RECT 43.340 37.030 43.510 37.200 ;
        RECT 43.750 37.030 43.920 37.200 ;
        RECT 44.280 37.030 44.450 37.200 ;
        RECT 44.640 37.030 44.810 37.200 ;
        RECT 45.000 37.030 45.170 37.200 ;
        RECT 45.840 37.030 46.010 37.200 ;
        RECT 46.200 37.030 46.370 37.200 ;
        RECT 46.560 37.030 46.730 37.200 ;
        RECT 47.400 37.030 47.570 37.200 ;
        RECT 47.760 37.030 47.930 37.200 ;
        RECT 48.120 37.030 48.290 37.200 ;
      LAYER L1M1_PR_C ;
        RECT 54.870 38.580 55.040 38.750 ;
      LAYER mcon ;
        RECT 49.180 37.030 49.350 37.200 ;
        RECT 49.620 37.030 49.790 37.200 ;
        RECT 50.060 37.030 50.230 37.200 ;
        RECT 50.470 37.030 50.640 37.200 ;
        RECT 51.000 37.030 51.170 37.200 ;
        RECT 51.360 37.030 51.530 37.200 ;
        RECT 51.720 37.030 51.890 37.200 ;
      LAYER L1M1_PR_C ;
        RECT 53.430 37.840 53.600 38.010 ;
      LAYER mcon ;
        RECT 52.560 37.030 52.730 37.200 ;
        RECT 52.920 37.030 53.090 37.200 ;
        RECT 53.280 37.030 53.450 37.200 ;
        RECT 54.120 37.030 54.290 37.200 ;
        RECT 54.480 37.030 54.650 37.200 ;
        RECT 54.840 37.030 55.010 37.200 ;
      LAYER L1M1_PR_C ;
        RECT 61.590 38.580 61.760 38.750 ;
        RECT 57.750 38.210 57.920 38.380 ;
      LAYER mcon ;
        RECT 55.900 37.030 56.070 37.200 ;
        RECT 56.340 37.030 56.510 37.200 ;
        RECT 56.780 37.030 56.950 37.200 ;
        RECT 57.190 37.030 57.360 37.200 ;
        RECT 57.720 37.030 57.890 37.200 ;
        RECT 58.080 37.030 58.250 37.200 ;
        RECT 58.440 37.030 58.610 37.200 ;
        RECT 59.280 37.030 59.450 37.200 ;
        RECT 59.640 37.030 59.810 37.200 ;
        RECT 60.000 37.030 60.170 37.200 ;
        RECT 60.840 37.030 61.010 37.200 ;
        RECT 61.200 37.030 61.370 37.200 ;
        RECT 61.560 37.030 61.730 37.200 ;
      LAYER L1M1_PR_C ;
        RECT 68.310 38.580 68.480 38.750 ;
        RECT 64.470 38.210 64.640 38.380 ;
      LAYER mcon ;
        RECT 62.620 37.030 62.790 37.200 ;
        RECT 63.060 37.030 63.230 37.200 ;
        RECT 63.500 37.030 63.670 37.200 ;
        RECT 63.910 37.030 64.080 37.200 ;
        RECT 64.440 37.030 64.610 37.200 ;
        RECT 64.800 37.030 64.970 37.200 ;
        RECT 65.160 37.030 65.330 37.200 ;
        RECT 66.000 37.030 66.170 37.200 ;
        RECT 66.360 37.030 66.530 37.200 ;
        RECT 66.720 37.030 66.890 37.200 ;
        RECT 67.560 37.030 67.730 37.200 ;
        RECT 67.920 37.030 68.090 37.200 ;
        RECT 68.280 37.030 68.450 37.200 ;
      LAYER L1M1_PR_C ;
        RECT 75.030 38.580 75.200 38.750 ;
        RECT 71.190 38.210 71.360 38.380 ;
        RECT 78.390 39.690 78.560 39.860 ;
      LAYER mcon ;
        RECT 69.340 37.030 69.510 37.200 ;
        RECT 69.780 37.030 69.950 37.200 ;
        RECT 70.220 37.030 70.390 37.200 ;
        RECT 70.630 37.030 70.800 37.200 ;
        RECT 71.160 37.030 71.330 37.200 ;
        RECT 71.520 37.030 71.690 37.200 ;
        RECT 71.880 37.030 72.050 37.200 ;
        RECT 72.720 37.030 72.890 37.200 ;
        RECT 73.080 37.030 73.250 37.200 ;
        RECT 73.440 37.030 73.610 37.200 ;
        RECT 74.280 37.030 74.450 37.200 ;
        RECT 74.640 37.030 74.810 37.200 ;
        RECT 75.000 37.030 75.170 37.200 ;
      LAYER L1M1_PR_C ;
        RECT 79.830 39.690 80.000 39.860 ;
      LAYER mcon ;
        RECT 76.060 37.030 76.230 37.200 ;
        RECT 76.500 37.030 76.670 37.200 ;
        RECT 76.940 37.030 77.110 37.200 ;
        RECT 77.350 37.030 77.520 37.200 ;
        RECT 78.790 37.030 78.960 37.200 ;
        RECT 79.150 37.030 79.320 37.200 ;
        RECT 79.510 37.030 79.680 37.200 ;
        RECT 79.870 37.030 80.040 37.200 ;
      LAYER L1M1_PR_C ;
        RECT 86.550 38.580 86.720 38.750 ;
      LAYER mcon ;
        RECT 80.860 37.030 81.030 37.200 ;
        RECT 81.300 37.030 81.470 37.200 ;
        RECT 81.740 37.030 81.910 37.200 ;
        RECT 82.150 37.030 82.320 37.200 ;
        RECT 82.680 37.030 82.850 37.200 ;
        RECT 83.040 37.030 83.210 37.200 ;
        RECT 83.400 37.030 83.570 37.200 ;
      LAYER L1M1_PR_C ;
        RECT 84.630 37.840 84.800 38.010 ;
      LAYER mcon ;
        RECT 84.240 37.030 84.410 37.200 ;
        RECT 84.600 37.030 84.770 37.200 ;
        RECT 84.960 37.030 85.130 37.200 ;
        RECT 85.800 37.030 85.970 37.200 ;
        RECT 86.160 37.030 86.330 37.200 ;
        RECT 86.520 37.030 86.690 37.200 ;
      LAYER L1M1_PR_C ;
        RECT 93.270 38.580 93.440 38.750 ;
        RECT 89.430 38.210 89.600 38.380 ;
      LAYER mcon ;
        RECT 87.580 37.030 87.750 37.200 ;
        RECT 88.020 37.030 88.190 37.200 ;
        RECT 88.460 37.030 88.630 37.200 ;
        RECT 88.870 37.030 89.040 37.200 ;
        RECT 89.400 37.030 89.570 37.200 ;
        RECT 89.760 37.030 89.930 37.200 ;
        RECT 90.120 37.030 90.290 37.200 ;
        RECT 90.960 37.030 91.130 37.200 ;
        RECT 91.320 37.030 91.490 37.200 ;
        RECT 91.680 37.030 91.850 37.200 ;
        RECT 92.520 37.030 92.690 37.200 ;
        RECT 92.880 37.030 93.050 37.200 ;
        RECT 93.240 37.030 93.410 37.200 ;
      LAYER L1M1_PR_C ;
        RECT 97.590 39.690 97.760 39.860 ;
        RECT 98.550 38.580 98.720 38.750 ;
        RECT 96.150 38.210 96.320 38.380 ;
        RECT 99.510 38.580 99.680 38.750 ;
        RECT 97.110 38.210 97.280 38.380 ;
      LAYER mcon ;
        RECT 94.300 37.030 94.470 37.200 ;
        RECT 94.740 37.030 94.910 37.200 ;
        RECT 95.180 37.030 95.350 37.200 ;
        RECT 95.590 37.030 95.760 37.200 ;
        RECT 98.200 37.030 98.370 37.200 ;
        RECT 98.560 37.030 98.730 37.200 ;
        RECT 98.920 37.030 99.090 37.200 ;
      LAYER L1M1_PR_C ;
        RECT 103.830 39.690 104.000 39.860 ;
        RECT 102.390 38.580 102.560 38.750 ;
        RECT 101.910 38.210 102.080 38.380 ;
        RECT 104.790 39.320 104.960 39.490 ;
      LAYER mcon ;
        RECT 100.060 37.030 100.230 37.200 ;
        RECT 100.500 37.030 100.670 37.200 ;
        RECT 100.940 37.030 101.110 37.200 ;
        RECT 101.350 37.030 101.520 37.200 ;
        RECT 101.880 37.030 102.050 37.200 ;
        RECT 102.240 37.030 102.410 37.200 ;
        RECT 103.150 37.030 103.320 37.200 ;
        RECT 103.510 37.030 103.680 37.200 ;
        RECT 103.870 37.030 104.040 37.200 ;
      LAYER L1M1_PR_C ;
        RECT 104.310 37.470 104.480 37.640 ;
        RECT 108.150 38.950 108.320 39.120 ;
        RECT 107.190 38.210 107.360 38.380 ;
      LAYER mcon ;
        RECT 105.340 37.030 105.510 37.200 ;
        RECT 105.780 37.030 105.950 37.200 ;
        RECT 106.220 37.030 106.390 37.200 ;
        RECT 106.630 37.030 106.800 37.200 ;
        RECT 107.160 37.030 107.330 37.200 ;
        RECT 107.520 37.030 107.690 37.200 ;
      LAYER L1M1_PR_C ;
        RECT 114.870 38.580 115.040 38.750 ;
        RECT 111.030 38.210 111.200 38.380 ;
      LAYER mcon ;
        RECT 108.700 37.030 108.870 37.200 ;
        RECT 109.140 37.030 109.310 37.200 ;
        RECT 109.580 37.030 109.750 37.200 ;
        RECT 109.990 37.030 110.160 37.200 ;
        RECT 111.000 37.030 111.170 37.200 ;
        RECT 111.360 37.030 111.530 37.200 ;
        RECT 111.720 37.030 111.890 37.200 ;
        RECT 112.560 37.030 112.730 37.200 ;
        RECT 112.920 37.030 113.090 37.200 ;
        RECT 113.280 37.030 113.450 37.200 ;
        RECT 114.120 37.030 114.290 37.200 ;
        RECT 114.480 37.030 114.650 37.200 ;
        RECT 114.840 37.030 115.010 37.200 ;
      LAYER L1M1_PR_C ;
        RECT 124.470 38.580 124.640 38.750 ;
        RECT 127.350 39.690 127.520 39.860 ;
      LAYER mcon ;
        RECT 116.430 37.020 116.600 37.190 ;
        RECT 116.870 37.020 117.040 37.190 ;
        RECT 117.280 37.020 117.450 37.190 ;
        RECT 117.710 37.020 117.880 37.190 ;
        RECT 118.150 37.020 118.320 37.190 ;
        RECT 118.560 37.020 118.730 37.190 ;
        RECT 120.600 37.030 120.770 37.200 ;
        RECT 120.960 37.030 121.130 37.200 ;
        RECT 121.320 37.030 121.490 37.200 ;
      LAYER L1M1_PR_C ;
        RECT 123.030 37.840 123.200 38.010 ;
      LAYER mcon ;
        RECT 122.160 37.030 122.330 37.200 ;
        RECT 122.520 37.030 122.690 37.200 ;
        RECT 122.880 37.030 123.050 37.200 ;
        RECT 123.720 37.030 123.890 37.200 ;
        RECT 124.080 37.030 124.250 37.200 ;
        RECT 124.440 37.030 124.610 37.200 ;
        RECT 125.500 37.030 125.670 37.200 ;
        RECT 125.940 37.030 126.110 37.200 ;
        RECT 126.380 37.030 126.550 37.200 ;
        RECT 126.790 37.030 126.960 37.200 ;
      LAYER L1M1_PR_C ;
        RECT 128.790 38.580 128.960 38.750 ;
        RECT 133.590 39.690 133.760 39.860 ;
        RECT 131.190 38.210 131.360 38.380 ;
      LAYER mcon ;
        RECT 127.800 37.030 127.970 37.200 ;
        RECT 128.310 37.030 128.480 37.200 ;
        RECT 129.990 37.030 130.160 37.200 ;
        RECT 130.350 37.030 130.520 37.200 ;
        RECT 130.710 37.030 130.880 37.200 ;
      LAYER L1M1_PR_C ;
        RECT 135.030 39.320 135.200 39.490 ;
      LAYER mcon ;
        RECT 131.740 37.030 131.910 37.200 ;
        RECT 132.180 37.030 132.350 37.200 ;
        RECT 132.620 37.030 132.790 37.200 ;
        RECT 133.030 37.030 133.200 37.200 ;
        RECT 133.990 37.030 134.160 37.200 ;
        RECT 134.350 37.030 134.520 37.200 ;
        RECT 134.710 37.030 134.880 37.200 ;
        RECT 135.070 37.030 135.240 37.200 ;
        RECT 136.060 37.030 136.230 37.200 ;
        RECT 136.500 37.030 136.670 37.200 ;
        RECT 136.940 37.030 137.110 37.200 ;
        RECT 137.350 37.030 137.520 37.200 ;
        RECT 139.360 37.030 139.530 37.200 ;
        RECT 139.720 37.030 139.890 37.200 ;
        RECT 140.380 37.030 140.550 37.200 ;
        RECT 140.820 37.030 140.990 37.200 ;
        RECT 141.260 37.030 141.430 37.200 ;
        RECT 141.670 37.030 141.840 37.200 ;
      LAYER L1M1_PR_C ;
        RECT 10.710 34.880 10.880 35.050 ;
        RECT 11.670 33.770 11.840 33.940 ;
        RECT 14.070 33.400 14.240 33.570 ;
        RECT 22.710 35.250 22.880 35.420 ;
        RECT 21.750 34.880 21.920 35.050 ;
        RECT 15.510 33.400 15.680 33.570 ;
        RECT 23.190 34.880 23.360 35.050 ;
        RECT 25.590 34.880 25.760 35.050 ;
        RECT 26.550 34.880 26.720 35.050 ;
        RECT 27.990 34.510 28.160 34.680 ;
        RECT 28.950 34.510 29.120 34.680 ;
        RECT 27.030 33.400 27.200 33.570 ;
        RECT 31.350 34.140 31.520 34.310 ;
        RECT 34.230 34.880 34.400 35.050 ;
        RECT 33.750 34.510 33.920 34.680 ;
        RECT 35.190 34.880 35.360 35.050 ;
        RECT 41.910 34.880 42.080 35.050 ;
        RECT 44.790 34.510 44.960 34.680 ;
        RECT 50.070 35.250 50.240 35.420 ;
        RECT 51.510 34.510 51.680 34.680 ;
        RECT 54.390 34.880 54.560 35.050 ;
        RECT 58.230 34.510 58.400 34.680 ;
        RECT 64.470 34.880 64.640 35.050 ;
        RECT 63.990 34.140 64.160 34.310 ;
        RECT 78.870 34.880 79.040 35.050 ;
        RECT 84.150 35.250 84.320 35.420 ;
        RECT 75.990 33.400 76.160 33.570 ;
        RECT 79.350 33.400 79.520 33.570 ;
        RECT 85.590 34.510 85.760 34.680 ;
        RECT 90.390 34.880 90.560 35.050 ;
        RECT 93.270 34.510 93.440 34.680 ;
        RECT 97.110 35.620 97.280 35.790 ;
        RECT 96.150 34.880 96.320 35.050 ;
        RECT 97.110 34.880 97.280 35.050 ;
        RECT 98.550 34.510 98.720 34.680 ;
        RECT 99.510 34.510 99.680 34.680 ;
        RECT 105.270 35.250 105.440 35.420 ;
        RECT 106.230 35.250 106.400 35.420 ;
        RECT 112.470 35.620 112.640 35.790 ;
        RECT 110.070 34.510 110.240 34.680 ;
        RECT 111.030 34.510 111.200 34.680 ;
        RECT 107.670 33.400 107.840 33.570 ;
        RECT 111.990 33.400 112.160 33.570 ;
        RECT 115.830 35.620 116.000 35.790 ;
        RECT 117.270 34.880 117.440 35.050 ;
        RECT 120.150 34.510 120.320 34.680 ;
        RECT 123.990 35.250 124.160 35.420 ;
        RECT 124.950 35.250 125.120 35.420 ;
        RECT 126.390 35.620 126.560 35.790 ;
        RECT 123.990 33.400 124.160 33.570 ;
        RECT 135.990 35.620 136.160 35.790 ;
        RECT 128.790 34.510 128.960 34.680 ;
        RECT 130.230 34.510 130.400 34.680 ;
        RECT 135.510 34.880 135.680 35.050 ;
        RECT 139.350 35.250 139.520 35.420 ;
        RECT 130.710 33.400 130.880 33.570 ;
        RECT 138.390 34.880 138.560 35.050 ;
        RECT 9.750 30.810 9.920 30.980 ;
      LAYER mcon ;
        RECT 7.310 28.890 7.480 29.060 ;
        RECT 7.670 28.890 7.840 29.060 ;
        RECT 8.030 28.890 8.200 29.060 ;
        RECT 8.950 28.890 9.120 29.060 ;
        RECT 9.310 28.890 9.480 29.060 ;
      LAYER L1M1_PR_C ;
        RECT 10.230 30.070 10.400 30.240 ;
      LAYER mcon ;
        RECT 13.910 28.890 14.080 29.060 ;
        RECT 14.270 28.890 14.440 29.060 ;
        RECT 14.630 28.890 14.800 29.060 ;
      LAYER L1M1_PR_C ;
        RECT 21.750 30.070 21.920 30.240 ;
      LAYER mcon ;
        RECT 17.880 28.890 18.050 29.060 ;
        RECT 18.240 28.890 18.410 29.060 ;
        RECT 18.600 28.890 18.770 29.060 ;
      LAYER L1M1_PR_C ;
        RECT 24.150 30.070 24.320 30.240 ;
      LAYER mcon ;
        RECT 20.490 28.890 20.660 29.060 ;
        RECT 20.850 28.890 21.020 29.060 ;
        RECT 21.210 28.890 21.380 29.060 ;
        RECT 22.300 28.890 22.470 29.060 ;
        RECT 22.740 28.890 22.910 29.060 ;
        RECT 23.180 28.890 23.350 29.060 ;
        RECT 23.590 28.890 23.760 29.060 ;
        RECT 24.120 28.890 24.290 29.060 ;
        RECT 24.480 28.890 24.650 29.060 ;
      LAYER L1M1_PR_C ;
        RECT 25.110 29.330 25.280 29.500 ;
        RECT 29.910 31.550 30.080 31.720 ;
        RECT 27.510 30.070 27.680 30.240 ;
        RECT 28.950 30.070 29.120 30.240 ;
        RECT 30.390 30.070 30.560 30.240 ;
      LAYER mcon ;
        RECT 25.660 28.890 25.830 29.060 ;
        RECT 26.100 28.890 26.270 29.060 ;
        RECT 26.540 28.890 26.710 29.060 ;
        RECT 26.950 28.890 27.120 29.060 ;
        RECT 27.740 28.890 27.910 29.060 ;
        RECT 28.100 28.890 28.270 29.060 ;
        RECT 28.460 28.890 28.630 29.060 ;
        RECT 28.820 28.890 28.990 29.060 ;
        RECT 29.180 28.890 29.350 29.060 ;
      LAYER L1M1_PR_C ;
        RECT 35.190 30.440 35.360 30.610 ;
        RECT 35.670 31.550 35.840 31.720 ;
        RECT 33.750 30.070 33.920 30.240 ;
        RECT 34.230 30.070 34.400 30.240 ;
      LAYER mcon ;
        RECT 30.070 28.890 30.240 29.060 ;
        RECT 30.430 28.890 30.600 29.060 ;
        RECT 30.940 28.890 31.110 29.060 ;
        RECT 31.380 28.890 31.550 29.060 ;
        RECT 31.820 28.890 31.990 29.060 ;
        RECT 32.230 28.890 32.400 29.060 ;
        RECT 33.020 28.890 33.190 29.060 ;
        RECT 33.380 28.890 33.550 29.060 ;
        RECT 33.740 28.890 33.910 29.060 ;
        RECT 34.100 28.890 34.270 29.060 ;
        RECT 34.460 28.890 34.630 29.060 ;
      LAYER L1M1_PR_C ;
        RECT 41.430 30.440 41.600 30.610 ;
        RECT 39.030 30.070 39.200 30.240 ;
        RECT 42.390 30.440 42.560 30.610 ;
        RECT 39.990 30.070 40.160 30.240 ;
      LAYER mcon ;
        RECT 35.350 28.890 35.520 29.060 ;
        RECT 35.710 28.890 35.880 29.060 ;
        RECT 36.220 28.890 36.390 29.060 ;
        RECT 36.660 28.890 36.830 29.060 ;
        RECT 37.100 28.890 37.270 29.060 ;
        RECT 37.510 28.890 37.680 29.060 ;
      LAYER L1M1_PR_C ;
        RECT 39.990 29.330 40.160 29.500 ;
      LAYER mcon ;
        RECT 41.080 28.890 41.250 29.060 ;
        RECT 41.440 28.890 41.610 29.060 ;
        RECT 41.800 28.890 41.970 29.060 ;
      LAYER L1M1_PR_C ;
        RECT 48.630 30.440 48.800 30.610 ;
      LAYER mcon ;
        RECT 42.940 28.890 43.110 29.060 ;
        RECT 43.380 28.890 43.550 29.060 ;
        RECT 43.820 28.890 43.990 29.060 ;
        RECT 44.230 28.890 44.400 29.060 ;
        RECT 44.760 28.890 44.930 29.060 ;
        RECT 45.120 28.890 45.290 29.060 ;
        RECT 45.480 28.890 45.650 29.060 ;
      LAYER L1M1_PR_C ;
        RECT 47.190 29.700 47.360 29.870 ;
      LAYER mcon ;
        RECT 46.320 28.890 46.490 29.060 ;
        RECT 46.680 28.890 46.850 29.060 ;
        RECT 47.040 28.890 47.210 29.060 ;
        RECT 47.880 28.890 48.050 29.060 ;
        RECT 48.240 28.890 48.410 29.060 ;
        RECT 48.600 28.890 48.770 29.060 ;
      LAYER L1M1_PR_C ;
        RECT 55.350 30.440 55.520 30.610 ;
        RECT 51.510 30.070 51.680 30.240 ;
      LAYER mcon ;
        RECT 49.660 28.890 49.830 29.060 ;
        RECT 50.100 28.890 50.270 29.060 ;
        RECT 50.540 28.890 50.710 29.060 ;
        RECT 50.950 28.890 51.120 29.060 ;
        RECT 51.480 28.890 51.650 29.060 ;
        RECT 51.840 28.890 52.010 29.060 ;
        RECT 52.200 28.890 52.370 29.060 ;
        RECT 53.040 28.890 53.210 29.060 ;
        RECT 53.400 28.890 53.570 29.060 ;
        RECT 53.760 28.890 53.930 29.060 ;
        RECT 54.600 28.890 54.770 29.060 ;
        RECT 54.960 28.890 55.130 29.060 ;
        RECT 55.320 28.890 55.490 29.060 ;
      LAYER L1M1_PR_C ;
        RECT 63.990 30.440 64.160 30.610 ;
      LAYER mcon ;
        RECT 56.910 28.880 57.080 29.050 ;
        RECT 57.350 28.880 57.520 29.050 ;
        RECT 57.760 28.880 57.930 29.050 ;
        RECT 58.190 28.880 58.360 29.050 ;
        RECT 58.630 28.880 58.800 29.050 ;
        RECT 59.040 28.880 59.210 29.050 ;
        RECT 60.120 28.890 60.290 29.060 ;
        RECT 60.480 28.890 60.650 29.060 ;
        RECT 60.840 28.890 61.010 29.060 ;
      LAYER L1M1_PR_C ;
        RECT 62.550 29.700 62.720 29.870 ;
      LAYER mcon ;
        RECT 61.680 28.890 61.850 29.060 ;
        RECT 62.040 28.890 62.210 29.060 ;
        RECT 62.400 28.890 62.570 29.060 ;
        RECT 63.240 28.890 63.410 29.060 ;
        RECT 63.600 28.890 63.770 29.060 ;
        RECT 63.960 28.890 64.130 29.060 ;
      LAYER L1M1_PR_C ;
        RECT 70.710 30.440 70.880 30.610 ;
        RECT 66.870 30.070 67.040 30.240 ;
      LAYER mcon ;
        RECT 65.020 28.890 65.190 29.060 ;
        RECT 65.460 28.890 65.630 29.060 ;
        RECT 65.900 28.890 66.070 29.060 ;
        RECT 66.310 28.890 66.480 29.060 ;
        RECT 66.840 28.890 67.010 29.060 ;
        RECT 67.200 28.890 67.370 29.060 ;
        RECT 67.560 28.890 67.730 29.060 ;
        RECT 68.400 28.890 68.570 29.060 ;
        RECT 68.760 28.890 68.930 29.060 ;
        RECT 69.120 28.890 69.290 29.060 ;
        RECT 69.960 28.890 70.130 29.060 ;
        RECT 70.320 28.890 70.490 29.060 ;
        RECT 70.680 28.890 70.850 29.060 ;
      LAYER L1M1_PR_C ;
        RECT 77.430 30.440 77.600 30.610 ;
        RECT 73.590 30.070 73.760 30.240 ;
      LAYER mcon ;
        RECT 71.740 28.890 71.910 29.060 ;
        RECT 72.180 28.890 72.350 29.060 ;
        RECT 72.620 28.890 72.790 29.060 ;
        RECT 73.030 28.890 73.200 29.060 ;
        RECT 73.560 28.890 73.730 29.060 ;
        RECT 73.920 28.890 74.090 29.060 ;
        RECT 74.280 28.890 74.450 29.060 ;
        RECT 75.120 28.890 75.290 29.060 ;
        RECT 75.480 28.890 75.650 29.060 ;
        RECT 75.840 28.890 76.010 29.060 ;
        RECT 76.680 28.890 76.850 29.060 ;
        RECT 77.040 28.890 77.210 29.060 ;
        RECT 77.400 28.890 77.570 29.060 ;
      LAYER L1M1_PR_C ;
        RECT 82.710 30.440 82.880 30.610 ;
        RECT 80.310 30.070 80.480 30.240 ;
        RECT 83.670 30.440 83.840 30.610 ;
        RECT 81.270 30.070 81.440 30.240 ;
      LAYER mcon ;
        RECT 78.460 28.890 78.630 29.060 ;
        RECT 78.900 28.890 79.070 29.060 ;
        RECT 79.340 28.890 79.510 29.060 ;
        RECT 79.750 28.890 79.920 29.060 ;
      LAYER L1M1_PR_C ;
        RECT 81.270 29.330 81.440 29.500 ;
      LAYER mcon ;
        RECT 82.360 28.890 82.530 29.060 ;
        RECT 82.720 28.890 82.890 29.060 ;
        RECT 83.080 28.890 83.250 29.060 ;
      LAYER L1M1_PR_C ;
        RECT 88.470 30.440 88.640 30.610 ;
        RECT 86.070 30.070 86.240 30.240 ;
        RECT 89.430 30.440 89.600 30.610 ;
        RECT 87.030 30.070 87.200 30.240 ;
      LAYER mcon ;
        RECT 84.220 28.890 84.390 29.060 ;
        RECT 84.660 28.890 84.830 29.060 ;
        RECT 85.100 28.890 85.270 29.060 ;
        RECT 85.510 28.890 85.680 29.060 ;
      LAYER L1M1_PR_C ;
        RECT 87.030 29.330 87.200 29.500 ;
      LAYER mcon ;
        RECT 88.120 28.890 88.290 29.060 ;
        RECT 88.480 28.890 88.650 29.060 ;
        RECT 88.840 28.890 89.010 29.060 ;
      LAYER L1M1_PR_C ;
        RECT 91.830 30.070 92.000 30.240 ;
      LAYER mcon ;
        RECT 89.980 28.890 90.150 29.060 ;
        RECT 90.420 28.890 90.590 29.060 ;
        RECT 90.860 28.890 91.030 29.060 ;
        RECT 91.270 28.890 91.440 29.060 ;
      LAYER L1M1_PR_C ;
        RECT 94.230 30.440 94.400 30.610 ;
        RECT 94.710 30.440 94.880 30.610 ;
        RECT 95.190 30.070 95.360 30.240 ;
        RECT 101.910 30.810 102.080 30.980 ;
      LAYER mcon ;
        RECT 92.240 28.890 92.410 29.060 ;
        RECT 92.600 28.890 92.770 29.060 ;
        RECT 92.960 28.890 93.130 29.060 ;
      LAYER L1M1_PR_C ;
        RECT 99.510 29.700 99.680 29.870 ;
        RECT 100.470 29.700 100.640 29.870 ;
      LAYER mcon ;
        RECT 95.600 28.890 95.770 29.060 ;
        RECT 95.960 28.890 96.130 29.060 ;
        RECT 96.320 28.890 96.490 29.060 ;
        RECT 96.680 28.890 96.850 29.060 ;
        RECT 97.180 28.890 97.350 29.060 ;
        RECT 97.620 28.890 97.790 29.060 ;
        RECT 98.060 28.890 98.230 29.060 ;
        RECT 98.470 28.890 98.640 29.060 ;
        RECT 98.980 28.890 99.150 29.060 ;
        RECT 99.340 28.890 99.510 29.060 ;
        RECT 99.700 28.890 99.870 29.060 ;
        RECT 100.950 28.890 101.120 29.060 ;
        RECT 101.310 28.890 101.480 29.060 ;
      LAYER L1M1_PR_C ;
        RECT 107.190 30.440 107.360 30.610 ;
        RECT 104.790 30.070 104.960 30.240 ;
        RECT 108.150 30.440 108.320 30.610 ;
        RECT 105.750 30.070 105.920 30.240 ;
      LAYER mcon ;
        RECT 102.460 28.890 102.630 29.060 ;
        RECT 102.900 28.890 103.070 29.060 ;
        RECT 103.340 28.890 103.510 29.060 ;
        RECT 103.750 28.890 103.920 29.060 ;
      LAYER L1M1_PR_C ;
        RECT 105.750 29.330 105.920 29.500 ;
      LAYER mcon ;
        RECT 106.840 28.890 107.010 29.060 ;
        RECT 107.200 28.890 107.370 29.060 ;
        RECT 107.560 28.890 107.730 29.060 ;
      LAYER L1M1_PR_C ;
        RECT 110.550 30.070 110.720 30.240 ;
      LAYER mcon ;
        RECT 108.700 28.890 108.870 29.060 ;
        RECT 109.140 28.890 109.310 29.060 ;
        RECT 109.580 28.890 109.750 29.060 ;
        RECT 109.990 28.890 110.160 29.060 ;
      LAYER L1M1_PR_C ;
        RECT 112.950 30.440 113.120 30.610 ;
        RECT 113.430 30.440 113.600 30.610 ;
        RECT 114.390 30.070 114.560 30.240 ;
        RECT 113.910 29.700 114.080 29.870 ;
        RECT 122.310 30.440 122.480 30.610 ;
        RECT 120.150 30.070 120.320 30.240 ;
        RECT 123.030 30.440 123.200 30.610 ;
        RECT 121.110 30.070 121.280 30.240 ;
      LAYER mcon ;
        RECT 110.960 28.890 111.130 29.060 ;
        RECT 111.320 28.890 111.490 29.060 ;
        RECT 111.680 28.890 111.850 29.060 ;
        RECT 114.320 28.890 114.490 29.060 ;
        RECT 114.680 28.890 114.850 29.060 ;
        RECT 115.040 28.890 115.210 29.060 ;
        RECT 115.400 28.890 115.570 29.060 ;
        RECT 116.430 28.880 116.600 29.050 ;
        RECT 116.870 28.880 117.040 29.050 ;
        RECT 117.280 28.880 117.450 29.050 ;
        RECT 117.710 28.880 117.880 29.050 ;
        RECT 118.150 28.880 118.320 29.050 ;
        RECT 118.560 28.880 118.730 29.050 ;
      LAYER L1M1_PR_C ;
        RECT 121.110 29.330 121.280 29.500 ;
      LAYER mcon ;
        RECT 122.200 28.890 122.370 29.060 ;
        RECT 122.560 28.890 122.730 29.060 ;
        RECT 122.920 28.890 123.090 29.060 ;
      LAYER L1M1_PR_C ;
        RECT 125.910 30.070 126.080 30.240 ;
        RECT 127.830 30.070 128.000 30.240 ;
      LAYER mcon ;
        RECT 124.060 28.890 124.230 29.060 ;
        RECT 124.500 28.890 124.670 29.060 ;
        RECT 124.940 28.890 125.110 29.060 ;
        RECT 125.350 28.890 125.520 29.060 ;
      LAYER L1M1_PR_C ;
        RECT 127.350 29.700 127.520 29.870 ;
        RECT 133.590 30.440 133.760 30.610 ;
        RECT 133.110 30.070 133.280 30.240 ;
      LAYER mcon ;
        RECT 125.880 28.890 126.050 29.060 ;
        RECT 126.240 28.890 126.410 29.060 ;
        RECT 126.600 28.890 126.770 29.060 ;
        RECT 126.960 28.890 127.130 29.060 ;
        RECT 128.910 28.880 129.080 29.050 ;
        RECT 129.350 28.880 129.520 29.050 ;
        RECT 129.760 28.880 129.930 29.050 ;
        RECT 130.190 28.880 130.360 29.050 ;
        RECT 130.630 28.880 130.800 29.050 ;
        RECT 131.040 28.880 131.210 29.050 ;
        RECT 132.600 28.890 132.770 29.060 ;
        RECT 132.960 28.890 133.130 29.060 ;
        RECT 134.670 28.880 134.840 29.050 ;
        RECT 135.110 28.880 135.280 29.050 ;
        RECT 135.520 28.880 135.690 29.050 ;
        RECT 135.950 28.880 136.120 29.050 ;
        RECT 136.390 28.880 136.560 29.050 ;
        RECT 136.800 28.880 136.970 29.050 ;
        RECT 138.510 28.880 138.680 29.050 ;
        RECT 138.950 28.880 139.120 29.050 ;
        RECT 139.360 28.880 139.530 29.050 ;
        RECT 139.790 28.880 139.960 29.050 ;
        RECT 140.230 28.880 140.400 29.050 ;
        RECT 140.640 28.880 140.810 29.050 ;
      LAYER L1M1_PR_C ;
        RECT 15.990 27.480 16.160 27.650 ;
        RECT 15.510 26.740 15.680 26.910 ;
        RECT 19.350 26.370 19.520 26.540 ;
        RECT 19.830 26.370 20.000 26.540 ;
        RECT 20.310 25.260 20.480 25.430 ;
        RECT 22.710 25.630 22.880 25.800 ;
        RECT 24.150 26.000 24.320 26.170 ;
        RECT 28.950 26.740 29.120 26.910 ;
        RECT 27.030 26.370 27.200 26.540 ;
        RECT 28.470 26.370 28.640 26.540 ;
        RECT 33.270 27.110 33.440 27.280 ;
        RECT 31.350 26.740 31.520 26.910 ;
        RECT 33.750 27.480 33.920 27.650 ;
        RECT 41.910 27.480 42.080 27.650 ;
        RECT 38.070 26.740 38.240 26.910 ;
        RECT 34.230 25.260 34.400 25.430 ;
        RECT 39.510 26.370 39.680 26.540 ;
        RECT 40.470 26.370 40.640 26.540 ;
        RECT 41.430 26.000 41.600 26.170 ;
        RECT 45.270 27.110 45.440 27.280 ;
        RECT 46.710 27.110 46.880 27.280 ;
        RECT 48.150 26.740 48.320 26.910 ;
        RECT 45.270 25.260 45.440 25.430 ;
        RECT 54.870 27.110 55.040 27.280 ;
        RECT 56.790 26.370 56.960 26.540 ;
        RECT 60.630 26.740 60.800 26.910 ;
        RECT 63.510 26.370 63.680 26.540 ;
        RECT 68.790 27.110 68.960 27.280 ;
        RECT 70.230 26.370 70.400 26.540 ;
        RECT 73.110 26.740 73.280 26.910 ;
        RECT 76.950 26.370 77.120 26.540 ;
        RECT 83.670 26.740 83.840 26.910 ;
        RECT 82.230 25.260 82.400 25.430 ;
        RECT 89.910 26.370 90.080 26.540 ;
        RECT 90.390 26.370 90.560 26.540 ;
        RECT 96.150 27.110 96.320 27.280 ;
        RECT 95.190 26.740 95.360 26.910 ;
        RECT 90.870 25.630 91.040 25.800 ;
        RECT 96.630 26.740 96.800 26.910 ;
        RECT 99.030 26.740 99.200 26.910 ;
        RECT 102.390 27.480 102.560 27.650 ;
        RECT 99.990 26.000 100.160 26.170 ;
        RECT 103.830 26.740 104.000 26.910 ;
        RECT 106.710 27.480 106.880 27.650 ;
        RECT 108.150 26.740 108.320 26.910 ;
        RECT 112.470 27.110 112.640 27.280 ;
        RECT 111.510 26.740 111.680 26.910 ;
        RECT 112.950 26.740 113.120 26.910 ;
        RECT 117.750 27.110 117.920 27.280 ;
        RECT 115.350 26.370 115.520 26.540 ;
        RECT 116.790 26.370 116.960 26.540 ;
        RECT 117.270 26.370 117.440 26.540 ;
        RECT 121.590 26.740 121.760 26.910 ;
        RECT 122.070 26.740 122.240 26.910 ;
        RECT 123.510 26.740 123.680 26.910 ;
        RECT 123.030 25.630 123.200 25.800 ;
        RECT 126.870 27.480 127.040 27.650 ;
        RECT 125.910 26.740 126.080 26.910 ;
        RECT 130.710 26.740 130.880 26.910 ;
        RECT 129.270 25.260 129.440 25.430 ;
      LAYER mcon ;
        RECT 6.510 20.740 6.680 20.910 ;
        RECT 6.950 20.740 7.120 20.910 ;
        RECT 7.360 20.740 7.530 20.910 ;
        RECT 7.790 20.740 7.960 20.910 ;
        RECT 8.230 20.740 8.400 20.910 ;
        RECT 8.640 20.740 8.810 20.910 ;
        RECT 12.160 20.750 12.330 20.920 ;
        RECT 12.520 20.750 12.690 20.920 ;
        RECT 13.710 20.740 13.880 20.910 ;
        RECT 14.150 20.740 14.320 20.910 ;
        RECT 14.560 20.740 14.730 20.910 ;
        RECT 14.990 20.740 15.160 20.910 ;
        RECT 15.430 20.740 15.600 20.910 ;
        RECT 15.840 20.740 16.010 20.910 ;
        RECT 18.880 20.750 19.050 20.920 ;
        RECT 19.240 20.750 19.410 20.920 ;
        RECT 19.900 20.750 20.070 20.920 ;
        RECT 20.340 20.750 20.510 20.920 ;
        RECT 20.780 20.750 20.950 20.920 ;
        RECT 21.190 20.750 21.360 20.920 ;
        RECT 23.200 20.750 23.370 20.920 ;
        RECT 23.560 20.750 23.730 20.920 ;
        RECT 24.220 20.750 24.390 20.920 ;
        RECT 24.660 20.750 24.830 20.920 ;
        RECT 25.100 20.750 25.270 20.920 ;
        RECT 25.510 20.750 25.680 20.920 ;
        RECT 26.510 20.750 26.680 20.920 ;
        RECT 26.870 20.750 27.040 20.920 ;
        RECT 27.230 20.750 27.400 20.920 ;
        RECT 28.150 20.750 28.320 20.920 ;
        RECT 28.510 20.750 28.680 20.920 ;
      LAYER L1M1_PR_C ;
        RECT 29.430 21.930 29.600 22.100 ;
      LAYER mcon ;
        RECT 33.110 20.750 33.280 20.920 ;
        RECT 33.470 20.750 33.640 20.920 ;
        RECT 33.830 20.750 34.000 20.920 ;
      LAYER L1M1_PR_C ;
        RECT 40.950 23.040 41.120 23.210 ;
      LAYER mcon ;
        RECT 37.080 20.750 37.250 20.920 ;
        RECT 37.440 20.750 37.610 20.920 ;
        RECT 37.800 20.750 37.970 20.920 ;
        RECT 39.690 20.750 39.860 20.920 ;
        RECT 40.050 20.750 40.220 20.920 ;
        RECT 40.410 20.750 40.580 20.920 ;
        RECT 42.030 20.740 42.200 20.910 ;
        RECT 42.470 20.740 42.640 20.910 ;
        RECT 42.880 20.740 43.050 20.910 ;
        RECT 43.310 20.740 43.480 20.910 ;
        RECT 43.750 20.740 43.920 20.910 ;
        RECT 44.160 20.740 44.330 20.910 ;
        RECT 45.720 20.750 45.890 20.920 ;
        RECT 46.080 20.750 46.250 20.920 ;
      LAYER L1M1_PR_C ;
        RECT 47.670 21.930 47.840 22.100 ;
      LAYER mcon ;
        RECT 47.590 20.750 47.760 20.920 ;
        RECT 47.950 20.750 48.120 20.920 ;
        RECT 50.010 20.750 50.180 20.920 ;
        RECT 50.370 20.750 50.540 20.920 ;
        RECT 50.730 20.750 50.900 20.920 ;
      LAYER L1M1_PR_C ;
        RECT 59.670 23.040 59.840 23.210 ;
        RECT 53.430 21.190 53.600 21.360 ;
      LAYER mcon ;
        RECT 51.950 20.750 52.120 20.920 ;
        RECT 52.310 20.750 52.480 20.920 ;
        RECT 52.670 20.750 52.840 20.920 ;
        RECT 56.490 20.750 56.660 20.920 ;
        RECT 56.850 20.750 57.020 20.920 ;
        RECT 58.410 20.750 58.580 20.920 ;
        RECT 58.770 20.750 58.940 20.920 ;
        RECT 59.130 20.750 59.300 20.920 ;
        RECT 60.750 20.740 60.920 20.910 ;
        RECT 61.190 20.740 61.360 20.910 ;
        RECT 61.600 20.740 61.770 20.910 ;
        RECT 62.030 20.740 62.200 20.910 ;
        RECT 62.470 20.740 62.640 20.910 ;
        RECT 62.880 20.740 63.050 20.910 ;
        RECT 64.430 20.750 64.600 20.920 ;
        RECT 64.790 20.750 64.960 20.920 ;
        RECT 65.150 20.750 65.320 20.920 ;
        RECT 66.070 20.750 66.240 20.920 ;
        RECT 66.430 20.750 66.600 20.920 ;
      LAYER L1M1_PR_C ;
        RECT 67.350 21.930 67.520 22.100 ;
      LAYER mcon ;
        RECT 71.030 20.750 71.200 20.920 ;
        RECT 71.390 20.750 71.560 20.920 ;
        RECT 71.750 20.750 71.920 20.920 ;
      LAYER L1M1_PR_C ;
        RECT 78.870 23.410 79.040 23.580 ;
      LAYER mcon ;
        RECT 75.000 20.750 75.170 20.920 ;
        RECT 75.360 20.750 75.530 20.920 ;
        RECT 75.720 20.750 75.890 20.920 ;
      LAYER L1M1_PR_C ;
        RECT 81.270 23.040 81.440 23.210 ;
        RECT 82.710 23.410 82.880 23.580 ;
      LAYER mcon ;
        RECT 77.610 20.750 77.780 20.920 ;
        RECT 77.970 20.750 78.140 20.920 ;
        RECT 78.330 20.750 78.500 20.920 ;
        RECT 79.420 20.750 79.590 20.920 ;
        RECT 79.860 20.750 80.030 20.920 ;
        RECT 80.300 20.750 80.470 20.920 ;
        RECT 80.710 20.750 80.880 20.920 ;
        RECT 81.670 20.750 81.840 20.920 ;
        RECT 82.030 20.750 82.200 20.920 ;
        RECT 82.390 20.750 82.560 20.920 ;
        RECT 82.750 20.750 82.920 20.920 ;
      LAYER L1M1_PR_C ;
        RECT 87.030 23.410 87.200 23.580 ;
      LAYER mcon ;
        RECT 83.740 20.750 83.910 20.920 ;
        RECT 84.180 20.750 84.350 20.920 ;
        RECT 84.620 20.750 84.790 20.920 ;
        RECT 85.030 20.750 85.200 20.920 ;
      LAYER L1M1_PR_C ;
        RECT 85.590 21.190 85.760 21.360 ;
      LAYER mcon ;
        RECT 85.990 20.750 86.160 20.920 ;
        RECT 86.350 20.750 86.520 20.920 ;
        RECT 86.710 20.750 86.880 20.920 ;
        RECT 87.070 20.750 87.240 20.920 ;
      LAYER L1M1_PR_C ;
        RECT 92.790 23.410 92.960 23.580 ;
        RECT 91.830 22.300 92.000 22.470 ;
        RECT 92.310 22.300 92.480 22.470 ;
      LAYER mcon ;
        RECT 88.060 20.750 88.230 20.920 ;
        RECT 88.500 20.750 88.670 20.920 ;
        RECT 88.940 20.750 89.110 20.920 ;
        RECT 89.350 20.750 89.520 20.920 ;
        RECT 90.830 20.750 91.000 20.920 ;
        RECT 91.190 20.750 91.360 20.920 ;
        RECT 91.550 20.750 91.720 20.920 ;
        RECT 92.470 20.750 92.640 20.920 ;
        RECT 92.830 20.750 93.000 20.920 ;
        RECT 93.340 20.750 93.510 20.920 ;
        RECT 93.780 20.750 93.950 20.920 ;
        RECT 94.220 20.750 94.390 20.920 ;
        RECT 94.630 20.750 94.800 20.920 ;
      LAYER L1M1_PR_C ;
        RECT 96.630 22.300 96.800 22.470 ;
        RECT 95.190 21.190 95.360 21.360 ;
      LAYER mcon ;
        RECT 95.590 20.750 95.760 20.920 ;
        RECT 95.950 20.750 96.120 20.920 ;
        RECT 96.310 20.750 96.480 20.920 ;
        RECT 96.670 20.750 96.840 20.920 ;
      LAYER L1M1_PR_C ;
        RECT 99.030 22.670 99.200 22.840 ;
        RECT 99.510 21.930 99.680 22.100 ;
        RECT 101.430 21.930 101.600 22.100 ;
      LAYER mcon ;
        RECT 97.660 20.750 97.830 20.920 ;
        RECT 98.100 20.750 98.270 20.920 ;
        RECT 98.540 20.750 98.710 20.920 ;
        RECT 98.950 20.750 99.120 20.920 ;
      LAYER L1M1_PR_C ;
        RECT 100.950 21.560 101.120 21.730 ;
      LAYER mcon ;
        RECT 99.480 20.750 99.650 20.920 ;
        RECT 99.840 20.750 100.010 20.920 ;
        RECT 100.200 20.750 100.370 20.920 ;
        RECT 100.560 20.750 100.730 20.920 ;
      LAYER L1M1_PR_C ;
        RECT 103.830 21.930 104.000 22.100 ;
        RECT 105.750 21.930 105.920 22.100 ;
      LAYER mcon ;
        RECT 101.980 20.750 102.150 20.920 ;
        RECT 102.420 20.750 102.590 20.920 ;
        RECT 102.860 20.750 103.030 20.920 ;
        RECT 103.270 20.750 103.440 20.920 ;
      LAYER L1M1_PR_C ;
        RECT 105.270 21.560 105.440 21.730 ;
      LAYER mcon ;
        RECT 103.800 20.750 103.970 20.920 ;
        RECT 104.160 20.750 104.330 20.920 ;
        RECT 104.520 20.750 104.690 20.920 ;
        RECT 104.880 20.750 105.050 20.920 ;
      LAYER L1M1_PR_C ;
        RECT 108.630 22.670 108.800 22.840 ;
      LAYER mcon ;
        RECT 106.300 20.750 106.470 20.920 ;
        RECT 106.740 20.750 106.910 20.920 ;
        RECT 107.180 20.750 107.350 20.920 ;
        RECT 107.590 20.750 107.760 20.920 ;
      LAYER L1M1_PR_C ;
        RECT 110.550 22.300 110.720 22.470 ;
        RECT 109.110 21.190 109.280 21.360 ;
      LAYER mcon ;
        RECT 109.510 20.750 109.680 20.920 ;
        RECT 109.870 20.750 110.040 20.920 ;
        RECT 110.230 20.750 110.400 20.920 ;
        RECT 110.590 20.750 110.760 20.920 ;
      LAYER L1M1_PR_C ;
        RECT 114.390 22.300 114.560 22.470 ;
        RECT 114.870 22.300 115.040 22.470 ;
        RECT 115.350 21.930 115.520 22.100 ;
      LAYER mcon ;
        RECT 111.580 20.750 111.750 20.920 ;
        RECT 112.020 20.750 112.190 20.920 ;
        RECT 112.460 20.750 112.630 20.920 ;
        RECT 112.870 20.750 113.040 20.920 ;
        RECT 113.390 20.750 113.560 20.920 ;
        RECT 113.750 20.750 113.920 20.920 ;
        RECT 114.110 20.750 114.280 20.920 ;
      LAYER L1M1_PR_C ;
        RECT 119.670 23.410 119.840 23.580 ;
        RECT 118.230 22.300 118.400 22.470 ;
        RECT 119.190 22.300 119.360 22.470 ;
      LAYER mcon ;
        RECT 115.030 20.750 115.200 20.920 ;
        RECT 115.390 20.750 115.560 20.920 ;
        RECT 115.900 20.750 116.070 20.920 ;
        RECT 116.340 20.750 116.510 20.920 ;
        RECT 116.780 20.750 116.950 20.920 ;
        RECT 117.190 20.750 117.360 20.920 ;
        RECT 117.710 20.750 117.880 20.920 ;
        RECT 118.070 20.750 118.240 20.920 ;
        RECT 118.430 20.750 118.600 20.920 ;
        RECT 119.350 20.750 119.520 20.920 ;
        RECT 119.710 20.750 119.880 20.920 ;
        RECT 120.220 20.750 120.390 20.920 ;
        RECT 120.660 20.750 120.830 20.920 ;
        RECT 121.100 20.750 121.270 20.920 ;
        RECT 121.510 20.750 121.680 20.920 ;
      LAYER L1M1_PR_C ;
        RECT 124.950 22.670 125.120 22.840 ;
      LAYER mcon ;
        RECT 122.510 20.750 122.680 20.920 ;
        RECT 122.870 20.750 123.040 20.920 ;
        RECT 123.230 20.750 123.400 20.920 ;
        RECT 124.150 20.750 124.320 20.920 ;
        RECT 124.510 20.750 124.680 20.920 ;
      LAYER L1M1_PR_C ;
        RECT 125.430 21.930 125.600 22.100 ;
      LAYER mcon ;
        RECT 129.110 20.750 129.280 20.920 ;
        RECT 129.470 20.750 129.640 20.920 ;
        RECT 129.830 20.750 130.000 20.920 ;
      LAYER L1M1_PR_C ;
        RECT 136.950 23.410 137.120 23.580 ;
      LAYER mcon ;
        RECT 133.080 20.750 133.250 20.920 ;
        RECT 133.440 20.750 133.610 20.920 ;
        RECT 133.800 20.750 133.970 20.920 ;
        RECT 135.690 20.750 135.860 20.920 ;
        RECT 136.050 20.750 136.220 20.920 ;
        RECT 136.410 20.750 136.580 20.920 ;
        RECT 138.030 20.740 138.200 20.910 ;
        RECT 138.470 20.740 138.640 20.910 ;
        RECT 138.880 20.740 139.050 20.910 ;
        RECT 139.310 20.740 139.480 20.910 ;
        RECT 139.750 20.740 139.920 20.910 ;
        RECT 140.160 20.740 140.330 20.910 ;
      LAYER L1M1_PR_C ;
        RECT 24.630 19.340 24.800 19.510 ;
        RECT 28.950 18.970 29.120 19.140 ;
        RECT 26.070 17.120 26.240 17.290 ;
        RECT 33.270 18.230 33.440 18.400 ;
        RECT 30.390 17.120 30.560 17.290 ;
        RECT 34.710 17.490 34.880 17.660 ;
        RECT 38.070 18.600 38.240 18.770 ;
        RECT 41.430 18.230 41.600 18.400 ;
        RECT 39.030 17.120 39.200 17.290 ;
        RECT 42.870 17.490 43.040 17.660 ;
        RECT 45.750 18.230 45.920 18.400 ;
        RECT 46.230 18.230 46.400 18.400 ;
        RECT 47.670 17.490 47.840 17.660 ;
        RECT 48.150 17.860 48.320 18.030 ;
        RECT 48.630 18.230 48.800 18.400 ;
        RECT 51.030 18.230 51.200 18.400 ;
        RECT 51.510 18.230 51.680 18.400 ;
        RECT 52.950 18.230 53.120 18.400 ;
        RECT 57.270 19.340 57.440 19.510 ;
        RECT 56.790 18.600 56.960 18.770 ;
        RECT 53.430 17.120 53.600 17.290 ;
        RECT 59.670 18.600 59.840 18.770 ;
        RECT 63.510 18.230 63.680 18.400 ;
        RECT 67.350 19.340 67.520 19.510 ;
        RECT 66.390 18.600 66.560 18.770 ;
        RECT 67.350 18.600 67.520 18.770 ;
        RECT 72.150 19.340 72.320 19.510 ;
        RECT 68.790 18.230 68.960 18.400 ;
        RECT 69.750 18.230 69.920 18.400 ;
        RECT 76.470 19.340 76.640 19.510 ;
        RECT 77.910 18.600 78.080 18.770 ;
        RECT 86.070 19.340 86.240 19.510 ;
        RECT 94.230 18.970 94.400 19.140 ;
        RECT 97.590 19.340 97.760 19.510 ;
        RECT 106.230 19.340 106.400 19.510 ;
        RECT 114.390 18.970 114.560 19.140 ;
        RECT 117.750 19.340 117.920 19.510 ;
      LAYER met1 ;
        RECT 108.090 144.920 108.380 144.970 ;
        RECT 117.200 144.920 117.520 144.980 ;
        RECT 95.690 144.780 117.520 144.920 ;
      LAYER met1 ;
        RECT 62.500 144.560 62.790 144.600 ;
        RECT 64.900 144.560 65.190 144.600 ;
        RECT 70.180 144.560 70.470 144.600 ;
        RECT 62.500 144.420 70.470 144.560 ;
        RECT 62.500 144.370 62.790 144.420 ;
        RECT 64.900 144.370 65.190 144.420 ;
        RECT 70.180 144.370 70.470 144.420 ;
      LAYER met1 ;
        RECT 20.730 144.180 21.020 144.230 ;
        RECT 32.720 144.180 33.040 144.240 ;
        RECT 20.730 144.040 33.040 144.180 ;
        RECT 20.730 144.000 21.020 144.040 ;
        RECT 32.720 143.980 33.040 144.040 ;
        RECT 38.010 144.180 38.300 144.230 ;
        RECT 49.520 144.180 49.840 144.240 ;
        RECT 51.930 144.180 52.220 144.230 ;
        RECT 38.010 144.040 52.220 144.180 ;
        RECT 38.010 144.000 38.300 144.040 ;
        RECT 49.520 143.980 49.840 144.040 ;
        RECT 51.930 144.000 52.220 144.040 ;
        RECT 61.050 144.180 61.340 144.230 ;
        RECT 77.840 144.180 78.160 144.240 ;
        RECT 61.050 144.040 65.110 144.180 ;
        RECT 77.640 144.040 78.160 144.180 ;
        RECT 61.050 144.000 61.340 144.040 ;
        RECT 64.970 143.870 65.110 144.040 ;
        RECT 77.840 143.980 78.160 144.040 ;
        RECT 87.450 144.180 87.740 144.230 ;
        RECT 95.690 144.180 95.830 144.780 ;
        RECT 108.090 144.740 108.380 144.780 ;
        RECT 117.200 144.720 117.520 144.780 ;
        RECT 99.440 144.180 99.760 144.240 ;
        RECT 87.450 144.040 95.830 144.180 ;
        RECT 99.240 144.040 99.760 144.180 ;
        RECT 87.450 144.000 87.740 144.040 ;
        RECT 64.880 143.610 65.200 143.870 ;
        RECT 72.090 143.810 72.380 143.860 ;
        RECT 87.530 143.810 87.670 144.000 ;
        RECT 99.440 143.980 99.760 144.040 ;
        RECT 72.090 143.670 87.670 143.810 ;
        RECT 72.090 143.630 72.380 143.670 ;
        RECT 28.890 143.440 29.180 143.490 ;
        RECT 30.800 143.440 31.120 143.500 ;
        RECT 36.560 143.440 36.880 143.500 ;
        RECT 28.890 143.300 31.120 143.440 ;
        RECT 36.360 143.300 36.880 143.440 ;
        RECT 28.890 143.260 29.180 143.300 ;
        RECT 30.800 143.240 31.120 143.300 ;
        RECT 36.560 143.240 36.880 143.300 ;
        RECT 50.000 143.440 50.320 143.500 ;
        RECT 50.490 143.440 50.780 143.490 ;
        RECT 50.000 143.300 50.780 143.440 ;
        RECT 50.000 143.240 50.320 143.300 ;
        RECT 50.490 143.260 50.780 143.300 ;
        RECT 63.930 143.440 64.220 143.490 ;
        RECT 70.640 143.440 70.960 143.500 ;
        RECT 86.000 143.440 86.320 143.500 ;
        RECT 63.930 143.300 70.960 143.440 ;
        RECT 85.800 143.300 86.320 143.440 ;
        RECT 63.930 143.260 64.220 143.300 ;
        RECT 70.640 143.240 70.960 143.300 ;
        RECT 86.000 143.240 86.320 143.300 ;
        RECT 98.010 143.440 98.300 143.490 ;
        RECT 98.480 143.440 98.800 143.500 ;
        RECT 106.640 143.440 106.960 143.500 ;
        RECT 98.010 143.300 98.800 143.440 ;
        RECT 106.440 143.300 106.960 143.440 ;
        RECT 98.010 143.260 98.300 143.300 ;
        RECT 98.480 143.240 98.800 143.300 ;
        RECT 106.640 143.240 106.960 143.300 ;
        RECT 5.760 142.710 142.080 143.080 ;
        RECT 33.210 141.590 33.500 141.640 ;
        RECT 36.560 141.590 36.880 141.650 ;
        RECT 33.210 141.450 36.880 141.590 ;
        RECT 33.210 141.410 33.500 141.450 ;
        RECT 36.560 141.390 36.880 141.450 ;
        RECT 50.000 141.590 50.320 141.650 ;
        RECT 50.490 141.590 50.780 141.640 ;
        RECT 50.000 141.450 50.780 141.590 ;
        RECT 50.000 141.390 50.320 141.450 ;
        RECT 50.490 141.410 50.780 141.450 ;
        RECT 64.880 141.590 65.200 141.650 ;
        RECT 81.690 141.590 81.980 141.640 ;
        RECT 86.000 141.590 86.320 141.650 ;
        RECT 64.880 141.450 65.400 141.590 ;
        RECT 81.690 141.450 86.320 141.590 ;
        RECT 64.880 141.390 65.200 141.450 ;
        RECT 81.690 141.410 81.980 141.450 ;
        RECT 86.000 141.390 86.320 141.450 ;
        RECT 98.480 141.220 98.800 141.280 ;
        RECT 98.280 141.080 98.800 141.220 ;
        RECT 98.480 141.020 98.800 141.080 ;
        RECT 106.640 141.220 106.960 141.280 ;
        RECT 109.530 141.220 109.820 141.270 ;
        RECT 106.640 141.080 109.820 141.220 ;
        RECT 106.640 141.020 106.960 141.080 ;
        RECT 109.530 141.040 109.820 141.080 ;
        RECT 33.680 140.850 34.000 140.910 ;
        RECT 33.480 140.710 34.000 140.850 ;
        RECT 33.680 140.650 34.000 140.710 ;
        RECT 44.240 140.850 44.560 140.910 ;
        RECT 50.970 140.850 51.260 140.900 ;
        RECT 44.240 140.710 51.260 140.850 ;
        RECT 44.240 140.650 44.560 140.710 ;
        RECT 50.970 140.670 51.260 140.710 ;
        RECT 71.610 140.850 71.900 140.900 ;
        RECT 77.840 140.850 78.160 140.910 ;
        RECT 71.610 140.710 78.160 140.850 ;
        RECT 71.610 140.670 71.900 140.710 ;
        RECT 77.840 140.650 78.160 140.710 ;
        RECT 82.170 140.850 82.460 140.900 ;
        RECT 86.960 140.850 87.280 140.910 ;
        RECT 101.360 140.850 101.680 140.910 ;
        RECT 82.170 140.710 87.280 140.850 ;
        RECT 101.160 140.710 101.680 140.850 ;
        RECT 82.170 140.670 82.460 140.710 ;
        RECT 86.960 140.650 87.280 140.710 ;
        RECT 101.360 140.650 101.680 140.710 ;
      LAYER met1 ;
        RECT 32.260 140.480 32.550 140.530 ;
        RECT 34.660 140.480 34.950 140.530 ;
        RECT 39.940 140.480 40.230 140.530 ;
        RECT 32.260 140.340 40.230 140.480 ;
        RECT 32.260 140.300 32.550 140.340 ;
        RECT 34.660 140.300 34.950 140.340 ;
        RECT 39.940 140.300 40.230 140.340 ;
        RECT 49.540 140.480 49.830 140.530 ;
        RECT 51.940 140.480 52.230 140.530 ;
        RECT 57.220 140.480 57.510 140.530 ;
        RECT 49.540 140.340 57.510 140.480 ;
        RECT 49.540 140.300 49.830 140.340 ;
        RECT 51.940 140.300 52.230 140.340 ;
        RECT 57.220 140.300 57.510 140.340 ;
      LAYER met1 ;
        RECT 74.490 140.480 74.780 140.530 ;
        RECT 79.290 140.480 79.580 140.530 ;
        RECT 74.490 140.340 79.580 140.480 ;
        RECT 74.490 140.300 74.780 140.340 ;
        RECT 79.290 140.300 79.580 140.340 ;
      LAYER met1 ;
        RECT 80.740 140.480 81.030 140.530 ;
        RECT 83.140 140.480 83.430 140.530 ;
        RECT 88.420 140.480 88.710 140.530 ;
        RECT 80.740 140.340 88.710 140.480 ;
        RECT 80.740 140.300 81.030 140.340 ;
        RECT 83.140 140.300 83.430 140.340 ;
        RECT 88.420 140.300 88.710 140.340 ;
        RECT 99.940 140.480 100.230 140.530 ;
        RECT 102.340 140.480 102.630 140.530 ;
        RECT 107.620 140.480 107.910 140.530 ;
        RECT 99.940 140.340 107.910 140.480 ;
        RECT 99.940 140.300 100.230 140.340 ;
        RECT 102.340 140.300 102.630 140.340 ;
        RECT 107.620 140.300 107.910 140.340 ;
      LAYER met1 ;
        RECT 72.090 139.740 72.380 139.790 ;
        RECT 78.320 139.740 78.640 139.800 ;
        RECT 99.440 139.740 99.760 139.800 ;
        RECT 72.090 139.600 78.640 139.740 ;
        RECT 72.090 139.560 72.380 139.600 ;
        RECT 78.320 139.540 78.640 139.600 ;
        RECT 92.810 139.600 99.760 139.740 ;
        RECT 66.320 139.370 66.640 139.430 ;
        RECT 66.120 139.230 66.640 139.370 ;
        RECT 66.320 139.170 66.640 139.230 ;
        RECT 74.960 139.370 75.280 139.430 ;
        RECT 75.930 139.370 76.220 139.420 ;
        RECT 92.810 139.370 92.950 139.600 ;
        RECT 99.440 139.540 99.760 139.600 ;
        RECT 93.680 139.370 94.000 139.430 ;
        RECT 74.960 139.230 92.950 139.370 ;
        RECT 93.480 139.230 94.000 139.370 ;
        RECT 74.960 139.170 75.280 139.230 ;
        RECT 75.930 139.190 76.220 139.230 ;
        RECT 93.680 139.170 94.000 139.230 ;
        RECT 100.880 139.370 101.200 139.430 ;
        RECT 112.890 139.370 113.180 139.420 ;
        RECT 100.880 139.230 113.180 139.370 ;
        RECT 100.880 139.170 101.200 139.230 ;
        RECT 112.890 139.190 113.180 139.230 ;
        RECT 63.930 137.520 64.220 137.570 ;
        RECT 66.320 137.520 66.640 137.580 ;
        RECT 63.930 137.380 66.640 137.520 ;
        RECT 63.930 137.340 64.220 137.380 ;
        RECT 66.320 137.320 66.640 137.380 ;
        RECT 99.440 137.150 99.760 137.210 ;
        RECT 99.440 137.010 102.070 137.150 ;
        RECT 99.440 136.950 99.760 137.010 ;
        RECT 30.800 136.780 31.120 136.840 ;
        RECT 30.600 136.640 31.120 136.780 ;
        RECT 30.800 136.580 31.120 136.640 ;
        RECT 70.640 136.780 70.960 136.840 ;
        RECT 76.890 136.780 77.180 136.830 ;
        RECT 86.960 136.780 87.280 136.840 ;
        RECT 98.490 136.780 98.780 136.830 ;
        RECT 101.360 136.780 101.680 136.840 ;
        RECT 70.640 136.640 77.180 136.780 ;
        RECT 86.760 136.640 87.280 136.780 ;
        RECT 70.640 136.580 70.960 136.640 ;
        RECT 76.890 136.600 77.180 136.640 ;
        RECT 86.960 136.580 87.280 136.640 ;
        RECT 88.970 136.640 98.230 136.780 ;
        RECT 32.250 136.410 32.540 136.460 ;
        RECT 49.520 136.410 49.840 136.470 ;
        RECT 32.250 136.270 49.840 136.410 ;
        RECT 32.250 136.230 32.540 136.270 ;
        RECT 49.520 136.210 49.840 136.270 ;
        RECT 77.850 136.230 78.140 136.460 ;
        RECT 78.320 136.410 78.640 136.470 ;
        RECT 78.320 136.270 78.840 136.410 ;
        RECT 75.450 135.860 75.740 136.090 ;
        RECT 76.410 136.040 76.700 136.090 ;
        RECT 77.360 136.040 77.680 136.100 ;
        RECT 76.410 135.900 77.680 136.040 ;
        RECT 77.930 136.040 78.070 136.230 ;
        RECT 78.320 136.210 78.640 136.270 ;
        RECT 85.040 136.040 85.360 136.100 ;
        RECT 88.970 136.040 89.110 136.640 ;
        RECT 89.370 136.410 89.660 136.460 ;
        RECT 93.680 136.410 94.000 136.470 ;
        RECT 89.370 136.270 94.000 136.410 ;
        RECT 89.370 136.230 89.660 136.270 ;
        RECT 93.680 136.210 94.000 136.270 ;
        RECT 89.850 136.040 90.140 136.090 ;
        RECT 77.930 135.900 90.140 136.040 ;
        RECT 76.410 135.860 76.700 135.900 ;
        RECT 36.080 135.300 36.400 135.360 ;
        RECT 35.880 135.160 36.400 135.300 ;
        RECT 75.530 135.300 75.670 135.860 ;
        RECT 77.360 135.840 77.680 135.900 ;
        RECT 85.040 135.840 85.360 135.900 ;
        RECT 89.850 135.860 90.140 135.900 ;
        RECT 90.810 136.040 91.100 136.090 ;
        RECT 94.160 136.040 94.480 136.100 ;
        RECT 90.810 135.900 94.480 136.040 ;
        RECT 98.090 136.040 98.230 136.640 ;
        RECT 98.490 136.640 101.680 136.780 ;
        RECT 101.930 136.780 102.070 137.010 ;
        RECT 110.010 136.780 110.300 136.830 ;
        RECT 110.960 136.780 111.280 136.840 ;
        RECT 101.930 136.640 111.280 136.780 ;
        RECT 98.490 136.600 98.780 136.640 ;
        RECT 101.360 136.580 101.680 136.640 ;
        RECT 110.010 136.600 110.300 136.640 ;
        RECT 110.960 136.580 111.280 136.640 ;
        RECT 100.880 136.410 101.200 136.470 ;
        RECT 102.800 136.410 103.120 136.470 ;
        RECT 100.680 136.270 101.200 136.410 ;
        RECT 100.880 136.210 101.200 136.270 ;
        RECT 101.450 136.270 103.120 136.410 ;
        RECT 101.450 136.090 101.590 136.270 ;
        RECT 102.800 136.210 103.120 136.270 ;
        RECT 101.370 136.040 101.660 136.090 ;
        RECT 98.090 135.900 101.660 136.040 ;
        RECT 90.810 135.860 91.100 135.900 ;
        RECT 94.160 135.840 94.480 135.900 ;
        RECT 101.370 135.860 101.660 135.900 ;
        RECT 101.840 136.040 102.160 136.100 ;
        RECT 111.440 136.040 111.760 136.100 ;
        RECT 101.840 135.900 102.360 136.040 ;
        RECT 111.240 135.900 111.760 136.040 ;
        RECT 101.840 135.840 102.160 135.900 ;
        RECT 111.440 135.840 111.760 135.900 ;
        RECT 117.200 136.040 117.520 136.100 ;
        RECT 118.640 136.040 118.960 136.100 ;
        RECT 119.610 136.040 119.900 136.090 ;
        RECT 117.200 135.900 119.900 136.040 ;
        RECT 117.200 135.840 117.520 135.900 ;
        RECT 118.640 135.840 118.960 135.900 ;
        RECT 119.610 135.860 119.900 135.900 ;
        RECT 90.330 135.670 90.620 135.720 ;
        RECT 101.370 135.670 101.660 135.720 ;
        RECT 102.320 135.670 102.640 135.730 ;
        RECT 90.330 135.530 102.640 135.670 ;
        RECT 90.330 135.490 90.620 135.530 ;
        RECT 101.370 135.490 101.660 135.530 ;
        RECT 102.320 135.470 102.640 135.530 ;
        RECT 107.600 135.300 107.920 135.360 ;
        RECT 118.160 135.300 118.480 135.360 ;
        RECT 75.530 135.160 107.920 135.300 ;
        RECT 117.960 135.160 118.480 135.300 ;
        RECT 36.080 135.100 36.400 135.160 ;
        RECT 107.600 135.100 107.920 135.160 ;
        RECT 118.160 135.100 118.480 135.160 ;
        RECT 5.760 134.570 142.080 134.940 ;
        RECT 32.720 133.450 33.040 133.510 ;
        RECT 32.520 133.310 33.040 133.450 ;
        RECT 32.720 133.250 33.040 133.310 ;
        RECT 85.050 133.450 85.340 133.500 ;
        RECT 101.840 133.450 102.160 133.510 ;
        RECT 107.600 133.450 107.920 133.510 ;
        RECT 85.050 133.310 102.160 133.450 ;
        RECT 107.400 133.310 107.920 133.450 ;
        RECT 85.050 133.270 85.340 133.310 ;
        RECT 101.840 133.250 102.160 133.310 ;
        RECT 107.600 133.250 107.920 133.310 ;
        RECT 113.850 133.450 114.140 133.500 ;
        RECT 118.160 133.450 118.480 133.510 ;
        RECT 113.850 133.310 118.480 133.450 ;
        RECT 113.850 133.270 114.140 133.310 ;
        RECT 118.160 133.250 118.480 133.310 ;
        RECT 74.490 133.080 74.780 133.130 ;
        RECT 125.850 133.080 126.140 133.130 ;
        RECT 74.490 132.940 79.510 133.080 ;
        RECT 74.490 132.900 74.780 132.940 ;
        RECT 29.360 132.710 29.680 132.770 ;
        RECT 31.770 132.710 32.060 132.760 ;
        RECT 29.360 132.570 32.060 132.710 ;
        RECT 29.360 132.510 29.680 132.570 ;
        RECT 31.770 132.530 32.060 132.570 ;
        RECT 32.730 132.710 33.020 132.760 ;
        RECT 39.440 132.710 39.760 132.770 ;
        RECT 32.730 132.570 39.760 132.710 ;
        RECT 32.730 132.530 33.020 132.570 ;
        RECT 39.440 132.510 39.760 132.570 ;
        RECT 79.370 132.400 79.510 132.940 ;
        RECT 100.490 132.940 126.140 133.080 ;
        RECT 88.890 132.530 89.180 132.760 ;
        RECT 89.370 132.710 89.660 132.760 ;
        RECT 93.680 132.710 94.000 132.770 ;
        RECT 89.370 132.570 94.000 132.710 ;
        RECT 89.370 132.530 89.660 132.570 ;
        RECT 34.170 132.160 34.460 132.390 ;
        RECT 35.130 132.340 35.420 132.390 ;
        RECT 36.080 132.340 36.400 132.400 ;
        RECT 78.810 132.340 79.100 132.390 ;
        RECT 35.130 132.200 79.100 132.340 ;
        RECT 35.130 132.160 35.420 132.200 ;
        RECT 34.250 131.970 34.390 132.160 ;
        RECT 36.080 132.140 36.400 132.200 ;
        RECT 78.810 132.160 79.100 132.200 ;
        RECT 79.280 132.340 79.600 132.400 ;
        RECT 80.240 132.340 80.560 132.400 ;
        RECT 87.450 132.340 87.740 132.390 ;
        RECT 79.280 132.200 79.800 132.340 ;
        RECT 80.240 132.200 87.740 132.340 ;
        RECT 79.280 132.140 79.600 132.200 ;
        RECT 80.240 132.140 80.560 132.200 ;
        RECT 87.450 132.160 87.740 132.200 ;
        RECT 87.920 132.340 88.240 132.400 ;
        RECT 88.970 132.340 89.110 132.530 ;
        RECT 93.680 132.510 94.000 132.570 ;
        RECT 99.920 132.340 100.240 132.400 ;
        RECT 100.490 132.390 100.630 132.940 ;
        RECT 101.360 132.710 101.680 132.770 ;
        RECT 102.320 132.710 102.640 132.770 ;
        RECT 105.770 132.760 105.910 132.940 ;
        RECT 125.850 132.900 126.140 132.940 ;
        RECT 101.160 132.570 101.680 132.710 ;
        RECT 102.120 132.570 102.640 132.710 ;
        RECT 101.360 132.510 101.680 132.570 ;
        RECT 102.320 132.510 102.640 132.570 ;
        RECT 105.690 132.530 105.980 132.760 ;
        RECT 106.170 132.530 106.460 132.760 ;
        RECT 114.330 132.710 114.620 132.760 ;
        RECT 106.730 132.570 114.620 132.710 ;
        RECT 87.920 132.200 88.440 132.340 ;
        RECT 88.970 132.200 100.240 132.340 ;
        RECT 87.920 132.140 88.240 132.200 ;
        RECT 99.920 132.140 100.240 132.200 ;
        RECT 100.410 132.160 100.700 132.390 ;
        RECT 100.890 132.340 101.180 132.390 ;
        RECT 102.800 132.340 103.120 132.400 ;
        RECT 100.890 132.200 103.120 132.340 ;
        RECT 100.890 132.160 101.180 132.200 ;
        RECT 102.800 132.140 103.120 132.200 ;
        RECT 103.280 132.340 103.600 132.400 ;
        RECT 106.250 132.340 106.390 132.530 ;
        RECT 103.280 132.200 106.390 132.340 ;
        RECT 103.280 132.140 103.600 132.200 ;
        RECT 36.560 131.970 36.880 132.030 ;
        RECT 34.250 131.830 36.880 131.970 ;
        RECT 36.560 131.770 36.880 131.830 ;
        RECT 98.010 131.970 98.300 132.020 ;
        RECT 98.010 131.830 103.030 131.970 ;
        RECT 98.010 131.790 98.300 131.830 ;
        RECT 80.730 131.600 81.020 131.650 ;
        RECT 83.600 131.600 83.920 131.660 ;
        RECT 80.730 131.460 83.920 131.600 ;
        RECT 102.890 131.600 103.030 131.830 ;
        RECT 106.730 131.600 106.870 132.570 ;
        RECT 114.330 132.530 114.620 132.570 ;
        RECT 107.600 132.340 107.920 132.400 ;
        RECT 107.400 132.200 107.920 132.340 ;
        RECT 107.600 132.140 107.920 132.200 ;
        RECT 110.960 132.340 111.280 132.400 ;
        RECT 111.450 132.340 111.740 132.390 ;
        RECT 110.960 132.200 111.740 132.340 ;
        RECT 110.960 132.140 111.280 132.200 ;
        RECT 111.450 132.160 111.740 132.200 ;
      LAYER met1 ;
        RECT 112.900 132.340 113.190 132.390 ;
        RECT 115.300 132.340 115.590 132.390 ;
        RECT 120.580 132.340 120.870 132.390 ;
        RECT 112.900 132.200 120.870 132.340 ;
        RECT 112.900 132.160 113.190 132.200 ;
        RECT 115.300 132.160 115.590 132.200 ;
        RECT 120.580 132.160 120.870 132.200 ;
      LAYER met1 ;
        RECT 102.890 131.460 106.870 131.600 ;
        RECT 80.730 131.420 81.020 131.460 ;
        RECT 83.600 131.400 83.920 131.460 ;
        RECT 76.400 131.230 76.720 131.290 ;
        RECT 76.200 131.090 76.720 131.230 ;
        RECT 76.400 131.030 76.720 131.090 ;
        RECT 81.200 131.230 81.520 131.290 ;
        RECT 81.200 131.090 81.720 131.230 ;
        RECT 81.200 131.030 81.520 131.090 ;
        RECT 33.680 129.380 34.000 129.440 ;
        RECT 34.650 129.380 34.940 129.430 ;
        RECT 36.560 129.380 36.880 129.440 ;
        RECT 33.680 129.240 34.940 129.380 ;
        RECT 36.360 129.240 36.880 129.380 ;
        RECT 33.680 129.180 34.000 129.240 ;
        RECT 34.650 129.200 34.940 129.240 ;
        RECT 36.560 129.180 36.880 129.240 ;
        RECT 83.130 129.380 83.420 129.430 ;
        RECT 87.920 129.380 88.240 129.440 ;
        RECT 83.130 129.240 88.240 129.380 ;
        RECT 83.130 129.200 83.420 129.240 ;
        RECT 87.920 129.180 88.240 129.240 ;
        RECT 97.530 129.380 97.820 129.430 ;
        RECT 101.360 129.380 101.680 129.440 ;
        RECT 97.530 129.240 101.680 129.380 ;
        RECT 97.530 129.200 97.820 129.240 ;
        RECT 101.360 129.180 101.680 129.240 ;
        RECT 110.960 129.380 111.280 129.440 ;
        RECT 112.410 129.380 112.700 129.430 ;
        RECT 110.960 129.240 112.700 129.380 ;
        RECT 110.960 129.180 111.280 129.240 ;
        RECT 112.410 129.200 112.700 129.240 ;
        RECT 36.560 128.640 36.880 128.700 ;
        RECT 42.800 128.640 43.120 128.700 ;
        RECT 100.880 128.640 101.200 128.700 ;
        RECT 36.560 128.500 46.870 128.640 ;
        RECT 36.560 128.440 36.880 128.500 ;
        RECT 42.800 128.440 43.120 128.500 ;
        RECT 46.730 128.320 46.870 128.500 ;
        RECT 100.010 128.500 101.200 128.640 ;
        RECT 43.850 128.130 45.430 128.270 ;
        RECT 16.880 127.900 17.200 127.960 ;
        RECT 16.680 127.760 17.200 127.900 ;
        RECT 16.880 127.700 17.200 127.760 ;
        RECT 39.440 127.900 39.760 127.960 ;
        RECT 43.850 127.900 43.990 128.130 ;
        RECT 45.290 127.950 45.430 128.130 ;
        RECT 45.690 128.090 45.980 128.320 ;
        RECT 46.650 128.090 46.940 128.320 ;
        RECT 47.610 128.270 47.900 128.320 ;
        RECT 79.280 128.270 79.600 128.330 ;
        RECT 82.170 128.270 82.460 128.320 ;
        RECT 47.610 128.130 68.950 128.270 ;
        RECT 47.610 128.090 47.900 128.130 ;
        RECT 39.440 127.760 43.990 127.900 ;
        RECT 39.440 127.700 39.760 127.760 ;
        RECT 44.250 127.720 44.540 127.950 ;
        RECT 45.210 127.720 45.500 127.950 ;
        RECT 45.770 127.900 45.910 128.090 ;
        RECT 52.410 127.900 52.700 127.950 ;
        RECT 45.770 127.760 52.700 127.900 ;
        RECT 52.410 127.720 52.700 127.760 ;
        RECT 26.000 127.530 26.320 127.590 ;
        RECT 44.330 127.530 44.470 127.720 ;
        RECT 26.000 127.390 44.470 127.530 ;
        RECT 45.290 127.530 45.430 127.720 ;
        RECT 47.600 127.530 47.920 127.590 ;
        RECT 68.810 127.580 68.950 128.130 ;
        RECT 78.410 128.130 82.460 128.270 ;
        RECT 75.440 127.900 75.760 127.960 ;
        RECT 78.410 127.950 78.550 128.130 ;
        RECT 79.280 128.070 79.600 128.130 ;
        RECT 82.170 128.090 82.460 128.130 ;
        RECT 82.650 128.270 82.940 128.320 ;
        RECT 83.600 128.270 83.920 128.330 ;
        RECT 82.650 128.130 83.920 128.270 ;
        RECT 82.650 128.090 82.940 128.130 ;
        RECT 75.240 127.760 75.760 127.900 ;
        RECT 75.440 127.700 75.760 127.760 ;
        RECT 78.330 127.720 78.620 127.950 ;
        RECT 80.730 127.720 81.020 127.950 ;
        RECT 82.250 127.900 82.390 128.090 ;
        RECT 83.600 128.070 83.920 128.130 ;
        RECT 95.120 128.270 95.440 128.330 ;
        RECT 100.010 128.320 100.150 128.500 ;
        RECT 100.880 128.440 101.200 128.500 ;
        RECT 98.970 128.270 99.260 128.320 ;
        RECT 95.120 128.130 99.260 128.270 ;
        RECT 95.120 128.070 95.440 128.130 ;
        RECT 98.970 128.090 99.260 128.130 ;
        RECT 99.930 128.090 100.220 128.320 ;
        RECT 100.400 128.270 100.720 128.330 ;
        RECT 103.280 128.270 103.600 128.330 ;
        RECT 100.400 128.130 103.600 128.270 ;
        RECT 100.400 128.070 100.720 128.130 ;
        RECT 103.280 128.070 103.600 128.130 ;
        RECT 83.120 127.900 83.440 127.960 ;
        RECT 82.250 127.760 83.440 127.900 ;
        RECT 45.290 127.390 47.920 127.530 ;
        RECT 26.000 127.330 26.320 127.390 ;
        RECT 47.600 127.330 47.920 127.390 ;
        RECT 68.730 127.530 69.020 127.580 ;
        RECT 80.810 127.530 80.950 127.720 ;
        RECT 83.120 127.700 83.440 127.760 ;
        RECT 100.880 127.900 101.200 127.960 ;
        RECT 118.160 127.900 118.480 127.960 ;
        RECT 120.090 127.900 120.380 127.950 ;
        RECT 100.880 127.760 101.400 127.900 ;
        RECT 118.160 127.760 120.380 127.900 ;
        RECT 100.880 127.700 101.200 127.760 ;
        RECT 118.160 127.700 118.480 127.760 ;
        RECT 120.090 127.720 120.380 127.760 ;
        RECT 68.730 127.390 80.950 127.530 ;
        RECT 68.730 127.350 69.020 127.390 ;
        RECT 15.440 127.160 15.760 127.220 ;
        RECT 15.240 127.020 15.760 127.160 ;
        RECT 15.440 126.960 15.760 127.020 ;
        RECT 31.760 127.160 32.080 127.220 ;
        RECT 37.530 127.160 37.820 127.210 ;
        RECT 58.160 127.160 58.480 127.220 ;
        RECT 31.760 127.020 37.820 127.160 ;
        RECT 57.960 127.020 58.480 127.160 ;
        RECT 31.760 126.960 32.080 127.020 ;
        RECT 37.530 126.980 37.820 127.020 ;
        RECT 58.160 126.960 58.480 127.020 ;
        RECT 74.490 127.160 74.780 127.210 ;
        RECT 80.240 127.160 80.560 127.220 ;
        RECT 74.490 127.020 80.560 127.160 ;
        RECT 74.490 126.980 74.780 127.020 ;
        RECT 80.240 126.960 80.560 127.020 ;
        RECT 110.970 127.160 111.260 127.210 ;
        RECT 111.920 127.160 112.240 127.220 ;
        RECT 118.640 127.160 118.960 127.220 ;
        RECT 110.970 127.020 112.240 127.160 ;
        RECT 118.440 127.020 118.960 127.160 ;
        RECT 110.970 126.980 111.260 127.020 ;
        RECT 111.920 126.960 112.240 127.020 ;
        RECT 118.640 126.960 118.960 127.020 ;
        RECT 5.760 126.430 142.080 126.800 ;
        RECT 11.130 125.310 11.420 125.360 ;
        RECT 15.440 125.310 15.760 125.370 ;
        RECT 44.240 125.310 44.560 125.370 ;
        RECT 58.160 125.310 58.480 125.370 ;
        RECT 77.360 125.310 77.680 125.370 ;
        RECT 94.160 125.310 94.480 125.370 ;
        RECT 11.130 125.170 15.760 125.310 ;
        RECT 44.040 125.170 44.560 125.310 ;
        RECT 57.960 125.170 58.480 125.310 ;
        RECT 77.160 125.170 77.680 125.310 ;
        RECT 93.960 125.170 94.480 125.310 ;
        RECT 11.130 125.130 11.420 125.170 ;
        RECT 15.440 125.110 15.760 125.170 ;
        RECT 44.240 125.110 44.560 125.170 ;
        RECT 58.160 125.110 58.480 125.170 ;
        RECT 77.360 125.110 77.680 125.170 ;
        RECT 94.160 125.110 94.480 125.170 ;
        RECT 114.330 125.310 114.620 125.360 ;
        RECT 118.640 125.310 118.960 125.370 ;
        RECT 114.330 125.170 118.960 125.310 ;
        RECT 114.330 125.130 114.620 125.170 ;
        RECT 118.640 125.110 118.960 125.170 ;
        RECT 38.000 124.940 38.320 125.000 ;
        RECT 107.600 124.940 107.920 125.000 ;
        RECT 111.920 124.940 112.240 125.000 ;
        RECT 126.330 124.940 126.620 124.990 ;
        RECT 37.800 124.800 38.320 124.940 ;
        RECT 38.000 124.740 38.320 124.800 ;
        RECT 102.410 124.800 107.920 124.940 ;
        RECT 111.720 124.800 112.240 124.940 ;
        RECT 11.610 124.570 11.900 124.620 ;
        RECT 20.240 124.570 20.560 124.630 ;
        RECT 29.840 124.570 30.160 124.630 ;
        RECT 11.610 124.430 20.560 124.570 ;
        RECT 29.640 124.430 30.160 124.570 ;
        RECT 11.610 124.390 11.900 124.430 ;
        RECT 20.240 124.370 20.560 124.430 ;
        RECT 29.840 124.370 30.160 124.430 ;
        RECT 41.360 124.570 41.680 124.630 ;
        RECT 47.130 124.570 47.420 124.620 ;
        RECT 41.360 124.430 47.420 124.570 ;
        RECT 41.360 124.370 41.680 124.430 ;
        RECT 47.130 124.390 47.420 124.430 ;
        RECT 47.600 124.570 47.920 124.630 ;
        RECT 81.200 124.570 81.520 124.630 ;
        RECT 47.600 124.430 48.120 124.570 ;
        RECT 76.010 124.430 81.520 124.570 ;
        RECT 47.600 124.370 47.920 124.430 ;
      LAYER met1 ;
        RECT 10.180 124.200 10.470 124.250 ;
        RECT 12.580 124.200 12.870 124.250 ;
        RECT 17.860 124.200 18.150 124.250 ;
        RECT 10.180 124.060 18.150 124.200 ;
        RECT 10.180 124.020 10.470 124.060 ;
        RECT 12.580 124.020 12.870 124.060 ;
        RECT 17.860 124.020 18.150 124.060 ;
        RECT 28.420 124.200 28.710 124.250 ;
        RECT 30.820 124.200 31.110 124.250 ;
        RECT 36.100 124.200 36.390 124.250 ;
        RECT 28.420 124.060 36.390 124.200 ;
        RECT 28.420 124.020 28.710 124.060 ;
        RECT 30.820 124.020 31.110 124.060 ;
        RECT 36.100 124.020 36.390 124.060 ;
      LAYER met1 ;
        RECT 42.800 124.200 43.120 124.260 ;
        RECT 46.170 124.200 46.460 124.250 ;
        RECT 42.800 124.060 46.460 124.200 ;
        RECT 42.800 124.000 43.120 124.060 ;
        RECT 46.170 124.020 46.460 124.060 ;
        RECT 74.970 124.200 75.260 124.250 ;
        RECT 75.440 124.200 75.760 124.260 ;
        RECT 76.010 124.250 76.150 124.430 ;
        RECT 81.200 124.370 81.520 124.430 ;
        RECT 89.840 124.570 90.160 124.630 ;
        RECT 90.810 124.570 91.100 124.620 ;
        RECT 98.000 124.570 98.320 124.630 ;
        RECT 101.360 124.570 101.680 124.630 ;
        RECT 89.840 124.430 91.100 124.570 ;
        RECT 97.800 124.430 98.320 124.570 ;
        RECT 101.160 124.430 101.680 124.570 ;
        RECT 89.840 124.370 90.160 124.430 ;
        RECT 90.810 124.390 91.100 124.430 ;
        RECT 98.000 124.370 98.320 124.430 ;
        RECT 101.360 124.370 101.680 124.430 ;
        RECT 101.840 124.570 102.160 124.630 ;
        RECT 102.410 124.620 102.550 124.800 ;
        RECT 107.600 124.740 107.920 124.800 ;
        RECT 111.920 124.740 112.240 124.800 ;
        RECT 112.490 124.800 126.620 124.940 ;
        RECT 102.330 124.570 102.620 124.620 ;
        RECT 101.840 124.430 102.620 124.570 ;
        RECT 101.840 124.370 102.160 124.430 ;
        RECT 102.330 124.390 102.620 124.430 ;
        RECT 107.130 124.570 107.420 124.620 ;
        RECT 112.490 124.570 112.630 124.800 ;
        RECT 126.330 124.760 126.620 124.800 ;
        RECT 114.800 124.570 115.120 124.630 ;
        RECT 107.130 124.430 112.630 124.570 ;
        RECT 114.600 124.430 115.120 124.570 ;
        RECT 107.130 124.390 107.420 124.430 ;
        RECT 74.970 124.060 75.760 124.200 ;
        RECT 74.970 124.020 75.260 124.060 ;
        RECT 75.440 124.000 75.760 124.060 ;
        RECT 75.930 124.020 76.220 124.250 ;
        RECT 76.400 124.200 76.720 124.260 ;
        RECT 76.890 124.200 77.180 124.250 ;
        RECT 95.120 124.200 95.440 124.260 ;
        RECT 95.610 124.200 95.900 124.250 ;
        RECT 76.400 124.060 77.180 124.200 ;
        RECT 76.400 124.000 76.720 124.060 ;
        RECT 76.890 124.020 77.180 124.060 ;
        RECT 91.850 124.060 95.900 124.200 ;
        RECT 75.530 123.830 75.670 124.000 ;
        RECT 91.850 123.880 91.990 124.060 ;
        RECT 95.120 124.000 95.440 124.060 ;
        RECT 95.610 124.020 95.900 124.060 ;
        RECT 96.570 124.020 96.860 124.250 ;
        RECT 97.050 124.200 97.340 124.250 ;
        RECT 97.520 124.200 97.840 124.260 ;
        RECT 100.400 124.200 100.720 124.260 ;
        RECT 103.760 124.200 104.080 124.260 ;
        RECT 104.720 124.200 105.040 124.260 ;
        RECT 97.050 124.060 100.720 124.200 ;
        RECT 103.560 124.060 104.080 124.200 ;
        RECT 104.520 124.060 105.040 124.200 ;
        RECT 97.050 124.020 97.340 124.060 ;
        RECT 91.770 123.830 92.060 123.880 ;
        RECT 75.530 123.690 92.060 123.830 ;
        RECT 96.650 123.830 96.790 124.020 ;
        RECT 97.520 124.000 97.840 124.060 ;
        RECT 100.400 124.000 100.720 124.060 ;
        RECT 103.760 124.000 104.080 124.060 ;
        RECT 104.720 124.000 105.040 124.060 ;
        RECT 107.210 123.830 107.350 124.390 ;
        RECT 114.800 124.370 115.120 124.430 ;
      LAYER met1 ;
        RECT 113.380 124.200 113.670 124.250 ;
        RECT 115.780 124.200 116.070 124.250 ;
        RECT 121.060 124.200 121.350 124.250 ;
        RECT 113.380 124.060 121.350 124.200 ;
        RECT 113.380 124.020 113.670 124.060 ;
        RECT 115.780 124.020 116.070 124.060 ;
        RECT 121.060 124.020 121.350 124.060 ;
      LAYER met1 ;
        RECT 96.650 123.690 107.350 123.830 ;
        RECT 91.770 123.650 92.060 123.690 ;
        RECT 102.810 123.460 103.100 123.510 ;
        RECT 112.880 123.460 113.200 123.520 ;
        RECT 102.810 123.320 113.200 123.460 ;
        RECT 102.810 123.280 103.100 123.320 ;
        RECT 112.880 123.260 113.200 123.320 ;
        RECT 23.130 123.090 23.420 123.140 ;
        RECT 25.040 123.090 25.360 123.150 ;
        RECT 41.360 123.090 41.680 123.150 ;
        RECT 23.130 122.950 25.360 123.090 ;
        RECT 41.160 122.950 41.680 123.090 ;
        RECT 23.130 122.910 23.420 122.950 ;
        RECT 25.040 122.890 25.360 122.950 ;
        RECT 41.360 122.890 41.680 122.950 ;
        RECT 57.680 123.090 58.000 123.150 ;
        RECT 59.610 123.090 59.900 123.140 ;
        RECT 108.080 123.090 108.400 123.150 ;
        RECT 57.680 122.950 59.900 123.090 ;
        RECT 107.880 122.950 108.400 123.090 ;
        RECT 57.680 122.890 58.000 122.950 ;
        RECT 59.610 122.910 59.900 122.950 ;
        RECT 108.080 122.890 108.400 122.950 ;
        RECT 20.240 121.240 20.560 121.300 ;
        RECT 20.040 121.100 20.560 121.240 ;
        RECT 20.240 121.040 20.560 121.100 ;
        RECT 28.890 121.240 29.180 121.290 ;
        RECT 29.840 121.240 30.160 121.300 ;
        RECT 28.890 121.100 30.160 121.240 ;
        RECT 28.890 121.060 29.180 121.100 ;
        RECT 29.840 121.040 30.160 121.100 ;
        RECT 36.090 121.240 36.380 121.290 ;
        RECT 38.000 121.240 38.320 121.300 ;
        RECT 36.090 121.100 38.320 121.240 ;
        RECT 36.090 121.060 36.380 121.100 ;
        RECT 38.000 121.040 38.320 121.100 ;
        RECT 43.770 121.240 44.060 121.290 ;
        RECT 49.520 121.240 49.840 121.300 ;
        RECT 88.400 121.240 88.720 121.300 ;
        RECT 43.770 121.100 88.720 121.240 ;
        RECT 43.770 121.060 44.060 121.100 ;
        RECT 49.520 121.040 49.840 121.100 ;
        RECT 88.400 121.040 88.720 121.100 ;
        RECT 95.610 121.240 95.900 121.290 ;
        RECT 103.760 121.240 104.080 121.300 ;
        RECT 95.610 121.100 104.080 121.240 ;
        RECT 95.610 121.060 95.900 121.100 ;
        RECT 103.760 121.040 104.080 121.100 ;
        RECT 105.690 121.240 105.980 121.290 ;
        RECT 114.800 121.240 115.120 121.300 ;
        RECT 105.690 121.100 115.120 121.240 ;
        RECT 105.690 121.060 105.980 121.100 ;
        RECT 114.800 121.040 115.120 121.100 ;
        RECT 33.680 120.870 34.000 120.930 ;
        RECT 45.210 120.870 45.500 120.920 ;
        RECT 57.680 120.870 58.000 120.930 ;
        RECT 16.490 120.730 58.000 120.870 ;
        RECT 12.090 120.500 12.380 120.550 ;
        RECT 16.490 120.500 16.630 120.730 ;
        RECT 33.680 120.670 34.000 120.730 ;
        RECT 45.210 120.690 45.500 120.730 ;
        RECT 57.680 120.670 58.000 120.730 ;
        RECT 74.960 120.870 75.280 120.930 ;
        RECT 75.450 120.870 75.740 120.920 ;
        RECT 74.960 120.730 75.740 120.870 ;
        RECT 74.960 120.670 75.280 120.730 ;
        RECT 75.450 120.690 75.740 120.730 ;
        RECT 86.000 120.870 86.320 120.930 ;
        RECT 101.840 120.870 102.160 120.930 ;
        RECT 86.000 120.730 96.310 120.870 ;
        RECT 101.640 120.730 102.160 120.870 ;
        RECT 86.000 120.670 86.320 120.730 ;
        RECT 12.090 120.360 16.630 120.500 ;
        RECT 16.880 120.500 17.200 120.560 ;
        RECT 37.530 120.500 37.820 120.550 ;
        RECT 40.880 120.500 41.200 120.560 ;
        RECT 68.720 120.500 69.040 120.560 ;
        RECT 16.880 120.360 41.200 120.500 ;
        RECT 68.280 120.360 90.550 120.500 ;
        RECT 12.090 120.320 12.380 120.360 ;
        RECT 16.880 120.300 17.200 120.360 ;
        RECT 37.530 120.320 37.820 120.360 ;
        RECT 40.880 120.300 41.200 120.360 ;
        RECT 68.720 120.300 69.040 120.360 ;
        RECT 22.170 120.130 22.460 120.180 ;
        RECT 26.960 120.130 27.280 120.190 ;
        RECT 30.810 120.130 31.100 120.180 ;
        RECT 41.360 120.130 41.680 120.190 ;
        RECT 78.320 120.130 78.640 120.190 ;
        RECT 79.760 120.130 80.080 120.190 ;
        RECT 90.410 120.180 90.550 120.360 ;
        RECT 94.640 120.300 94.960 120.560 ;
        RECT 22.170 119.990 31.100 120.130 ;
        RECT 22.170 119.950 22.460 119.990 ;
        RECT 26.960 119.930 27.280 119.990 ;
        RECT 30.810 119.950 31.100 119.990 ;
        RECT 33.290 119.990 41.680 120.130 ;
        RECT 78.120 119.990 78.640 120.130 ;
        RECT 79.560 119.990 80.080 120.130 ;
        RECT 24.570 119.580 24.860 119.810 ;
        RECT 25.040 119.760 25.360 119.820 ;
        RECT 31.760 119.760 32.080 119.820 ;
        RECT 33.290 119.810 33.430 119.990 ;
        RECT 41.360 119.930 41.680 119.990 ;
        RECT 78.320 119.930 78.640 119.990 ;
        RECT 79.760 119.930 80.080 119.990 ;
        RECT 90.330 119.950 90.620 120.180 ;
        RECT 91.770 120.130 92.060 120.180 ;
        RECT 94.730 120.130 94.870 120.300 ;
        RECT 91.770 119.990 94.870 120.130 ;
        RECT 91.770 119.950 92.060 119.990 ;
        RECT 25.040 119.620 32.080 119.760 ;
        RECT 24.650 119.390 24.790 119.580 ;
        RECT 25.040 119.560 25.360 119.620 ;
        RECT 31.760 119.560 32.080 119.620 ;
        RECT 33.210 119.580 33.500 119.810 ;
        RECT 33.690 119.580 33.980 119.810 ;
        RECT 52.890 119.760 53.180 119.810 ;
        RECT 62.480 119.760 62.800 119.820 ;
        RECT 52.890 119.620 62.800 119.760 ;
        RECT 52.890 119.580 53.180 119.620 ;
        RECT 25.520 119.390 25.840 119.450 ;
        RECT 33.770 119.390 33.910 119.580 ;
        RECT 62.480 119.560 62.800 119.620 ;
        RECT 78.800 119.760 79.120 119.820 ;
        RECT 80.250 119.760 80.540 119.810 ;
        RECT 78.800 119.620 80.540 119.760 ;
        RECT 78.800 119.560 79.120 119.620 ;
        RECT 80.250 119.580 80.540 119.620 ;
        RECT 83.130 119.760 83.420 119.810 ;
        RECT 85.520 119.760 85.840 119.820 ;
        RECT 83.130 119.620 85.840 119.760 ;
        RECT 83.130 119.580 83.420 119.620 ;
        RECT 85.520 119.560 85.840 119.620 ;
        RECT 86.490 119.580 86.780 119.810 ;
        RECT 92.250 119.760 92.540 119.810 ;
        RECT 94.160 119.760 94.480 119.820 ;
        RECT 95.120 119.760 95.440 119.820 ;
        RECT 96.170 119.810 96.310 120.730 ;
        RECT 101.840 120.670 102.160 120.730 ;
        RECT 101.930 120.130 102.070 120.670 ;
        RECT 102.320 120.500 102.640 120.560 ;
        RECT 102.320 120.360 107.350 120.500 ;
        RECT 102.320 120.300 102.640 120.360 ;
        RECT 107.210 120.190 107.350 120.360 ;
        RECT 106.640 120.130 106.960 120.190 ;
        RECT 101.930 119.990 105.430 120.130 ;
        RECT 106.440 119.990 106.960 120.130 ;
        RECT 92.250 119.620 94.480 119.760 ;
        RECT 94.920 119.620 95.440 119.760 ;
        RECT 92.250 119.580 92.540 119.620 ;
        RECT 24.650 119.250 33.910 119.390 ;
        RECT 86.570 119.390 86.710 119.580 ;
        RECT 94.160 119.560 94.480 119.620 ;
        RECT 95.120 119.560 95.440 119.620 ;
        RECT 96.090 119.580 96.380 119.810 ;
        RECT 96.570 119.580 96.860 119.810 ;
        RECT 97.520 119.760 97.840 119.820 ;
        RECT 105.290 119.810 105.430 119.990 ;
        RECT 106.640 119.930 106.960 119.990 ;
        RECT 107.120 120.130 107.440 120.190 ;
        RECT 107.120 119.990 107.880 120.130 ;
        RECT 107.120 119.930 107.440 119.990 ;
        RECT 97.320 119.620 97.840 119.760 ;
        RECT 89.840 119.390 90.160 119.450 ;
        RECT 86.570 119.250 90.160 119.390 ;
        RECT 25.520 119.190 25.840 119.250 ;
        RECT 89.840 119.190 90.160 119.250 ;
        RECT 93.680 119.390 94.000 119.450 ;
        RECT 96.650 119.390 96.790 119.580 ;
        RECT 97.520 119.560 97.840 119.620 ;
        RECT 101.370 119.580 101.660 119.810 ;
        RECT 104.250 119.580 104.540 119.810 ;
        RECT 105.210 119.580 105.500 119.810 ;
        RECT 93.680 119.250 96.790 119.390 ;
        RECT 93.680 119.190 94.000 119.250 ;
        RECT 23.120 119.020 23.440 119.080 ;
        RECT 60.560 119.020 60.880 119.080 ;
        RECT 22.920 118.880 23.440 119.020 ;
        RECT 60.360 118.880 60.880 119.020 ;
        RECT 23.120 118.820 23.440 118.880 ;
        RECT 60.560 118.820 60.880 118.880 ;
        RECT 71.600 119.020 71.920 119.080 ;
        RECT 74.010 119.020 74.300 119.070 ;
        RECT 71.600 118.880 74.300 119.020 ;
        RECT 71.600 118.820 71.920 118.880 ;
        RECT 74.010 118.840 74.300 118.880 ;
        RECT 81.680 119.020 82.000 119.080 ;
        RECT 83.610 119.020 83.900 119.070 ;
        RECT 81.680 118.880 83.900 119.020 ;
        RECT 81.680 118.820 82.000 118.880 ;
        RECT 83.610 118.840 83.900 118.880 ;
        RECT 87.930 119.020 88.220 119.070 ;
        RECT 95.120 119.020 95.440 119.080 ;
        RECT 87.930 118.880 95.440 119.020 ;
        RECT 101.450 119.020 101.590 119.580 ;
        RECT 104.330 119.390 104.470 119.580 ;
        RECT 108.080 119.390 108.400 119.450 ;
        RECT 104.330 119.250 108.400 119.390 ;
        RECT 108.080 119.190 108.400 119.250 ;
        RECT 108.560 119.020 108.880 119.080 ;
        RECT 101.450 118.880 108.880 119.020 ;
        RECT 87.930 118.840 88.220 118.880 ;
        RECT 95.120 118.820 95.440 118.880 ;
        RECT 108.560 118.820 108.880 118.880 ;
        RECT 5.760 118.290 142.080 118.660 ;
        RECT 60.560 117.170 60.880 117.230 ;
        RECT 86.000 117.170 86.320 117.230 ;
        RECT 60.360 117.030 60.880 117.170 ;
        RECT 85.800 117.030 86.320 117.170 ;
        RECT 60.560 116.970 60.880 117.030 ;
        RECT 86.000 116.970 86.320 117.030 ;
        RECT 93.210 117.170 93.500 117.220 ;
        RECT 106.640 117.170 106.960 117.230 ;
        RECT 93.210 117.030 106.960 117.170 ;
        RECT 93.210 116.990 93.500 117.030 ;
        RECT 106.640 116.970 106.960 117.030 ;
        RECT 47.600 116.800 47.920 116.860 ;
        RECT 43.850 116.660 47.920 116.800 ;
        RECT 43.850 116.490 43.990 116.660 ;
        RECT 47.600 116.600 47.920 116.660 ;
        RECT 50.010 116.800 50.300 116.850 ;
        RECT 52.400 116.800 52.720 116.860 ;
        RECT 71.600 116.800 71.920 116.860 ;
        RECT 50.010 116.660 52.720 116.800 ;
        RECT 71.400 116.660 71.920 116.800 ;
        RECT 50.010 116.620 50.300 116.660 ;
        RECT 52.400 116.600 52.720 116.660 ;
        RECT 71.600 116.600 71.920 116.660 ;
        RECT 88.400 116.800 88.720 116.860 ;
        RECT 111.920 116.800 112.240 116.860 ;
        RECT 88.400 116.660 112.240 116.800 ;
        RECT 88.400 116.600 88.720 116.660 ;
        RECT 111.920 116.600 112.240 116.660 ;
        RECT 15.450 116.430 15.740 116.480 ;
        RECT 16.880 116.430 17.200 116.490 ;
        RECT 15.450 116.290 17.200 116.430 ;
        RECT 15.450 116.250 15.740 116.290 ;
        RECT 16.880 116.230 17.200 116.290 ;
        RECT 23.120 116.430 23.440 116.490 ;
        RECT 25.040 116.430 25.360 116.490 ;
        RECT 23.120 116.290 25.360 116.430 ;
        RECT 23.120 116.230 23.440 116.290 ;
        RECT 25.040 116.230 25.360 116.290 ;
        RECT 26.010 116.430 26.300 116.480 ;
        RECT 29.360 116.430 29.680 116.490 ;
        RECT 42.810 116.430 43.100 116.480 ;
        RECT 43.760 116.430 44.080 116.490 ;
        RECT 61.520 116.430 61.840 116.490 ;
        RECT 26.010 116.290 43.100 116.430 ;
        RECT 43.320 116.290 44.080 116.430 ;
        RECT 26.010 116.250 26.300 116.290 ;
        RECT 29.360 116.230 29.680 116.290 ;
        RECT 42.810 116.250 43.100 116.290 ;
        RECT 43.760 116.230 44.080 116.290 ;
        RECT 46.250 116.290 61.840 116.430 ;
        RECT 46.250 116.110 46.390 116.290 ;
        RECT 61.520 116.230 61.840 116.290 ;
        RECT 74.490 116.430 74.780 116.480 ;
        RECT 82.640 116.430 82.960 116.490 ;
        RECT 74.490 116.290 82.960 116.430 ;
        RECT 74.490 116.250 74.780 116.290 ;
        RECT 82.640 116.230 82.960 116.290 ;
        RECT 89.840 116.430 90.160 116.490 ;
        RECT 90.330 116.430 90.620 116.480 ;
        RECT 96.570 116.430 96.860 116.480 ;
        RECT 89.840 116.290 96.860 116.430 ;
        RECT 89.840 116.230 90.160 116.290 ;
        RECT 90.330 116.250 90.620 116.290 ;
        RECT 96.570 116.250 96.860 116.290 ;
        RECT 97.530 116.430 97.820 116.480 ;
        RECT 101.840 116.430 102.160 116.490 ;
        RECT 104.720 116.430 105.040 116.490 ;
        RECT 97.530 116.290 101.110 116.430 ;
        RECT 101.640 116.290 102.160 116.430 ;
        RECT 104.520 116.290 105.040 116.430 ;
        RECT 97.530 116.250 97.820 116.290 ;
        RECT 45.210 116.060 45.500 116.110 ;
        RECT 42.890 115.920 45.500 116.060 ;
        RECT 42.890 115.750 43.030 115.920 ;
        RECT 45.210 115.880 45.500 115.920 ;
        RECT 46.170 115.880 46.460 116.110 ;
        RECT 52.410 116.060 52.700 116.110 ;
        RECT 56.720 116.060 57.040 116.120 ;
        RECT 57.680 116.060 58.000 116.120 ;
        RECT 62.010 116.060 62.300 116.110 ;
        RECT 52.410 115.920 57.040 116.060 ;
        RECT 57.480 115.920 62.300 116.060 ;
        RECT 52.410 115.880 52.700 115.920 ;
        RECT 56.720 115.860 57.040 115.920 ;
        RECT 57.680 115.860 58.000 115.920 ;
        RECT 62.010 115.880 62.300 115.920 ;
      LAYER met1 ;
        RECT 73.060 116.060 73.350 116.110 ;
        RECT 75.460 116.060 75.750 116.110 ;
        RECT 80.740 116.060 81.030 116.110 ;
        RECT 73.060 115.920 81.030 116.060 ;
        RECT 73.060 115.880 73.350 115.920 ;
        RECT 75.460 115.880 75.750 115.920 ;
        RECT 80.740 115.880 81.030 115.920 ;
      LAYER met1 ;
        RECT 95.120 116.060 95.440 116.120 ;
        RECT 95.610 116.060 95.900 116.110 ;
        RECT 95.120 115.920 95.900 116.060 ;
        RECT 95.120 115.860 95.440 115.920 ;
        RECT 95.610 115.880 95.900 115.920 ;
        RECT 96.080 116.060 96.400 116.120 ;
        RECT 100.410 116.060 100.700 116.110 ;
        RECT 100.970 116.060 101.110 116.290 ;
        RECT 101.840 116.230 102.160 116.290 ;
        RECT 104.720 116.230 105.040 116.290 ;
        RECT 110.960 116.430 111.280 116.490 ;
        RECT 112.890 116.430 113.180 116.480 ;
        RECT 110.960 116.290 113.180 116.430 ;
        RECT 110.960 116.230 111.280 116.290 ;
        RECT 112.890 116.250 113.180 116.290 ;
        RECT 122.010 116.430 122.300 116.480 ;
        RECT 124.400 116.430 124.720 116.490 ;
        RECT 122.010 116.290 124.720 116.430 ;
        RECT 122.010 116.250 122.300 116.290 ;
        RECT 124.400 116.230 124.720 116.290 ;
        RECT 101.360 116.060 101.680 116.120 ;
        RECT 108.560 116.060 108.880 116.120 ;
        RECT 96.080 115.920 96.600 116.060 ;
        RECT 97.130 115.920 100.700 116.060 ;
        RECT 100.920 115.920 103.510 116.060 ;
        RECT 108.360 115.920 108.880 116.060 ;
        RECT 96.080 115.860 96.400 115.920 ;
        RECT 37.520 115.690 37.840 115.750 ;
        RECT 42.800 115.690 43.120 115.750 ;
        RECT 37.520 115.550 43.120 115.690 ;
        RECT 37.520 115.490 37.840 115.550 ;
        RECT 42.800 115.490 43.120 115.550 ;
        RECT 56.250 115.690 56.540 115.740 ;
        RECT 61.040 115.690 61.360 115.750 ;
        RECT 56.250 115.550 61.360 115.690 ;
        RECT 56.250 115.510 56.540 115.550 ;
        RECT 61.040 115.490 61.360 115.550 ;
        RECT 72.080 115.690 72.400 115.750 ;
        RECT 74.010 115.690 74.300 115.740 ;
        RECT 72.080 115.550 74.300 115.690 ;
        RECT 72.080 115.490 72.400 115.550 ;
        RECT 74.010 115.510 74.300 115.550 ;
        RECT 85.040 115.690 85.360 115.750 ;
        RECT 97.130 115.690 97.270 115.920 ;
        RECT 100.410 115.880 100.700 115.920 ;
        RECT 101.360 115.860 101.680 115.920 ;
        RECT 85.040 115.550 97.270 115.690 ;
        RECT 85.040 115.490 85.360 115.550 ;
        RECT 44.250 115.320 44.540 115.370 ;
        RECT 52.880 115.320 53.200 115.380 ;
        RECT 44.250 115.180 53.200 115.320 ;
        RECT 44.250 115.140 44.540 115.180 ;
        RECT 52.880 115.120 53.200 115.180 ;
        RECT 64.880 115.320 65.200 115.380 ;
        RECT 66.810 115.320 67.100 115.370 ;
        RECT 64.880 115.180 67.100 115.320 ;
        RECT 64.880 115.120 65.200 115.180 ;
        RECT 66.810 115.140 67.100 115.180 ;
        RECT 68.250 115.320 68.540 115.370 ;
        RECT 71.600 115.320 71.920 115.380 ;
        RECT 97.520 115.320 97.840 115.380 ;
        RECT 68.250 115.180 71.920 115.320 ;
        RECT 68.250 115.140 68.540 115.180 ;
        RECT 71.600 115.120 71.920 115.180 ;
        RECT 93.290 115.180 97.840 115.320 ;
        RECT 103.370 115.320 103.510 115.920 ;
        RECT 108.560 115.860 108.880 115.920 ;
        RECT 103.370 115.180 113.590 115.320 ;
        RECT 14.000 114.950 14.320 115.010 ;
        RECT 13.800 114.810 14.320 114.950 ;
        RECT 14.000 114.750 14.320 114.810 ;
        RECT 87.920 114.950 88.240 115.010 ;
        RECT 88.890 114.950 89.180 115.000 ;
        RECT 93.290 114.950 93.430 115.180 ;
        RECT 97.520 115.120 97.840 115.180 ;
        RECT 87.920 114.810 93.430 114.950 ;
        RECT 110.000 114.950 110.320 115.010 ;
        RECT 111.450 114.950 111.740 115.000 ;
        RECT 110.000 114.810 111.740 114.950 ;
        RECT 113.450 114.950 113.590 115.180 ;
        RECT 116.330 115.180 119.350 115.320 ;
        RECT 116.330 114.950 116.470 115.180 ;
        RECT 117.200 114.950 117.520 115.010 ;
        RECT 113.450 114.810 116.470 114.950 ;
        RECT 117.000 114.810 117.520 114.950 ;
        RECT 87.920 114.750 88.240 114.810 ;
        RECT 88.890 114.770 89.180 114.810 ;
        RECT 110.000 114.750 110.320 114.810 ;
        RECT 111.450 114.770 111.740 114.810 ;
        RECT 117.200 114.750 117.520 114.810 ;
        RECT 118.160 114.950 118.480 115.010 ;
        RECT 118.650 114.950 118.940 115.000 ;
        RECT 118.160 114.810 118.940 114.950 ;
        RECT 119.210 114.950 119.350 115.180 ;
        RECT 122.490 114.950 122.780 115.000 ;
        RECT 119.210 114.810 122.780 114.950 ;
        RECT 118.160 114.750 118.480 114.810 ;
        RECT 118.650 114.770 118.940 114.810 ;
        RECT 122.490 114.770 122.780 114.810 ;
        RECT 20.730 113.100 21.020 113.150 ;
        RECT 25.040 113.100 25.360 113.160 ;
        RECT 72.080 113.100 72.400 113.160 ;
        RECT 82.640 113.100 82.960 113.160 ;
        RECT 20.730 112.960 25.360 113.100 ;
        RECT 71.880 112.960 72.400 113.100 ;
        RECT 82.440 112.960 82.960 113.100 ;
        RECT 20.730 112.920 21.020 112.960 ;
        RECT 25.040 112.900 25.360 112.960 ;
        RECT 72.080 112.900 72.400 112.960 ;
        RECT 82.640 112.900 82.960 112.960 ;
        RECT 89.850 113.100 90.140 113.150 ;
        RECT 93.680 113.100 94.000 113.160 ;
        RECT 124.400 113.100 124.720 113.160 ;
        RECT 89.850 112.960 94.000 113.100 ;
        RECT 124.200 112.960 124.720 113.100 ;
        RECT 89.850 112.920 90.140 112.960 ;
        RECT 93.680 112.900 94.000 112.960 ;
        RECT 124.400 112.900 124.720 112.960 ;
        RECT 8.730 112.360 9.020 112.410 ;
        RECT 14.000 112.360 14.320 112.420 ;
        RECT 8.730 112.220 14.320 112.360 ;
        RECT 8.730 112.180 9.020 112.220 ;
        RECT 14.000 112.160 14.320 112.220 ;
        RECT 86.000 112.160 86.320 112.420 ;
        RECT 107.120 112.360 107.440 112.420 ;
        RECT 87.050 112.220 107.440 112.360 ;
      LAYER met1 ;
        RECT 7.780 112.000 8.070 112.040 ;
        RECT 10.180 112.000 10.470 112.040 ;
        RECT 15.460 112.000 15.750 112.040 ;
        RECT 7.780 111.860 15.750 112.000 ;
      LAYER met1 ;
        RECT 26.480 111.990 26.800 112.050 ;
      LAYER met1 ;
        RECT 7.780 111.810 8.070 111.860 ;
        RECT 10.180 111.810 10.470 111.860 ;
        RECT 15.460 111.810 15.750 111.860 ;
      LAYER met1 ;
        RECT 24.650 111.850 26.800 111.990 ;
        RECT 24.650 111.670 24.790 111.850 ;
        RECT 26.480 111.790 26.800 111.850 ;
        RECT 26.960 111.990 27.280 112.050 ;
        RECT 27.930 111.990 28.220 112.040 ;
        RECT 29.360 111.990 29.680 112.050 ;
        RECT 26.960 111.850 27.480 111.990 ;
        RECT 27.930 111.850 29.680 111.990 ;
        RECT 26.960 111.790 27.280 111.850 ;
        RECT 27.930 111.810 28.220 111.850 ;
        RECT 29.360 111.790 29.680 111.850 ;
        RECT 45.690 111.810 45.980 112.040 ;
        RECT 52.400 111.990 52.720 112.050 ;
        RECT 52.200 111.850 52.720 111.990 ;
        RECT 24.570 111.440 24.860 111.670 ;
        RECT 25.040 111.620 25.360 111.680 ;
        RECT 25.530 111.620 25.820 111.670 ;
        RECT 25.040 111.480 25.820 111.620 ;
        RECT 25.040 111.420 25.360 111.480 ;
        RECT 25.530 111.440 25.820 111.480 ;
        RECT 38.970 111.440 39.260 111.670 ;
        RECT 45.770 111.620 45.910 111.810 ;
        RECT 52.400 111.790 52.720 111.850 ;
        RECT 59.130 111.810 59.420 112.040 ;
        RECT 66.320 111.990 66.640 112.050 ;
        RECT 66.810 111.990 67.100 112.040 ;
        RECT 66.320 111.850 67.100 111.990 ;
        RECT 55.290 111.620 55.580 111.670 ;
        RECT 45.770 111.480 55.580 111.620 ;
        RECT 59.210 111.620 59.350 111.810 ;
        RECT 66.320 111.790 66.640 111.850 ;
        RECT 66.810 111.810 67.100 111.850 ;
        RECT 74.960 111.990 75.280 112.050 ;
        RECT 79.770 111.990 80.060 112.040 ;
        RECT 74.960 111.850 80.060 111.990 ;
        RECT 74.960 111.790 75.280 111.850 ;
        RECT 79.770 111.810 80.060 111.850 ;
        RECT 85.050 111.990 85.340 112.040 ;
        RECT 86.090 111.990 86.230 112.160 ;
        RECT 85.050 111.850 86.230 111.990 ;
        RECT 85.050 111.810 85.340 111.850 ;
        RECT 64.400 111.620 64.720 111.680 ;
        RECT 73.530 111.620 73.820 111.670 ;
        RECT 59.210 111.480 73.820 111.620 ;
        RECT 55.290 111.440 55.580 111.480 ;
        RECT 9.210 111.250 9.500 111.300 ;
        RECT 9.210 111.110 25.750 111.250 ;
        RECT 9.210 111.070 9.500 111.110 ;
        RECT 25.610 110.930 25.750 111.110 ;
        RECT 25.530 110.700 25.820 110.930 ;
        RECT 37.520 110.880 37.840 110.940 ;
        RECT 37.320 110.740 37.840 110.880 ;
        RECT 39.050 110.880 39.190 111.440 ;
        RECT 64.400 111.420 64.720 111.480 ;
        RECT 73.530 111.440 73.820 111.480 ;
        RECT 78.810 111.620 79.100 111.670 ;
        RECT 82.160 111.620 82.480 111.680 ;
        RECT 78.810 111.480 82.480 111.620 ;
        RECT 78.810 111.440 79.100 111.480 ;
        RECT 82.160 111.420 82.480 111.480 ;
        RECT 85.530 111.440 85.820 111.670 ;
        RECT 86.480 111.620 86.800 111.680 ;
        RECT 87.050 111.670 87.190 112.220 ;
        RECT 107.120 112.160 107.440 112.220 ;
        RECT 99.930 111.810 100.220 112.040 ;
        RECT 100.400 111.990 100.720 112.050 ;
        RECT 106.650 111.990 106.940 112.040 ;
        RECT 110.000 111.990 110.320 112.050 ;
        RECT 100.400 111.850 106.940 111.990 ;
        RECT 109.800 111.850 110.320 111.990 ;
        RECT 86.280 111.480 86.800 111.620 ;
        RECT 44.250 111.250 44.540 111.300 ;
        RECT 44.720 111.250 45.040 111.310 ;
        RECT 44.250 111.110 45.040 111.250 ;
        RECT 44.250 111.070 44.540 111.110 ;
        RECT 44.720 111.050 45.040 111.110 ;
        RECT 50.970 111.250 51.260 111.300 ;
        RECT 62.000 111.250 62.320 111.310 ;
        RECT 65.360 111.250 65.680 111.310 ;
        RECT 50.970 111.110 62.320 111.250 ;
        RECT 65.160 111.110 65.680 111.250 ;
        RECT 50.970 111.070 51.260 111.110 ;
        RECT 62.000 111.050 62.320 111.110 ;
        RECT 65.360 111.050 65.680 111.110 ;
        RECT 80.720 111.250 81.040 111.310 ;
        RECT 85.040 111.250 85.360 111.310 ;
        RECT 85.610 111.250 85.750 111.440 ;
        RECT 86.480 111.420 86.800 111.480 ;
        RECT 86.970 111.440 87.260 111.670 ;
        RECT 91.760 111.620 92.080 111.680 ;
        RECT 91.560 111.480 92.080 111.620 ;
        RECT 91.760 111.420 92.080 111.480 ;
        RECT 93.690 111.440 93.980 111.670 ;
        RECT 96.080 111.620 96.400 111.680 ;
        RECT 95.880 111.480 96.400 111.620 ;
        RECT 100.010 111.620 100.150 111.810 ;
        RECT 100.400 111.790 100.720 111.850 ;
        RECT 106.650 111.810 106.940 111.850 ;
        RECT 110.000 111.790 110.320 111.850 ;
      LAYER met1 ;
        RECT 111.460 112.000 111.750 112.040 ;
        RECT 113.860 112.000 114.150 112.040 ;
        RECT 119.140 112.000 119.430 112.040 ;
        RECT 111.460 111.860 119.430 112.000 ;
        RECT 111.460 111.810 111.750 111.860 ;
        RECT 113.860 111.810 114.150 111.860 ;
        RECT 119.140 111.810 119.430 111.860 ;
      LAYER met1 ;
        RECT 102.810 111.620 103.100 111.670 ;
        RECT 112.880 111.620 113.200 111.680 ;
        RECT 100.010 111.480 103.100 111.620 ;
        RECT 112.680 111.480 113.200 111.620 ;
        RECT 80.720 111.110 85.750 111.250 ;
        RECT 93.770 111.250 93.910 111.440 ;
        RECT 96.080 111.420 96.400 111.480 ;
        RECT 102.810 111.440 103.100 111.480 ;
        RECT 112.880 111.420 113.200 111.480 ;
        RECT 105.680 111.250 106.000 111.310 ;
        RECT 93.770 111.110 106.000 111.250 ;
        RECT 80.720 111.050 81.040 111.110 ;
        RECT 85.040 111.050 85.360 111.110 ;
        RECT 105.680 111.050 106.000 111.110 ;
        RECT 117.200 111.250 117.520 111.310 ;
        RECT 121.050 111.250 121.340 111.300 ;
        RECT 117.200 111.110 121.340 111.250 ;
        RECT 117.200 111.050 117.520 111.110 ;
        RECT 121.050 111.070 121.340 111.110 ;
        RECT 52.400 110.880 52.720 110.940 ;
        RECT 39.050 110.740 52.720 110.880 ;
        RECT 37.520 110.680 37.840 110.740 ;
        RECT 52.400 110.680 52.720 110.740 ;
        RECT 79.280 110.880 79.600 110.940 ;
        RECT 79.770 110.880 80.060 110.930 ;
        RECT 79.280 110.740 80.060 110.880 ;
        RECT 79.280 110.680 79.600 110.740 ;
        RECT 79.770 110.700 80.060 110.740 ;
        RECT 5.760 110.150 142.080 110.520 ;
        RECT 52.880 109.030 53.200 109.090 ;
        RECT 52.680 108.890 53.200 109.030 ;
        RECT 52.880 108.830 53.200 108.890 ;
        RECT 83.600 109.030 83.920 109.090 ;
        RECT 85.040 109.030 85.360 109.090 ;
        RECT 107.120 109.030 107.440 109.090 ;
        RECT 112.410 109.030 112.700 109.080 ;
        RECT 113.840 109.030 114.160 109.090 ;
        RECT 83.600 108.890 88.630 109.030 ;
        RECT 83.600 108.830 83.920 108.890 ;
        RECT 85.040 108.830 85.360 108.890 ;
        RECT 61.040 108.660 61.360 108.720 ;
        RECT 69.200 108.660 69.520 108.720 ;
        RECT 60.840 108.520 61.360 108.660 ;
        RECT 69.000 108.520 69.520 108.660 ;
        RECT 61.040 108.460 61.360 108.520 ;
        RECT 69.200 108.460 69.520 108.520 ;
        RECT 76.010 108.520 87.190 108.660 ;
        RECT 23.120 108.290 23.440 108.350 ;
        RECT 24.080 108.290 24.400 108.350 ;
        RECT 26.960 108.290 27.280 108.350 ;
        RECT 31.760 108.290 32.080 108.350 ;
        RECT 22.920 108.150 23.440 108.290 ;
        RECT 23.880 108.150 24.400 108.290 ;
        RECT 23.120 108.090 23.440 108.150 ;
        RECT 24.080 108.090 24.400 108.150 ;
        RECT 25.610 108.150 27.280 108.290 ;
        RECT 31.560 108.150 32.080 108.290 ;
        RECT 25.610 107.970 25.750 108.150 ;
        RECT 26.960 108.090 27.280 108.150 ;
        RECT 31.760 108.090 32.080 108.150 ;
        RECT 32.240 108.290 32.560 108.350 ;
        RECT 76.010 108.340 76.150 108.520 ;
        RECT 32.240 108.150 32.760 108.290 ;
        RECT 32.240 108.090 32.560 108.150 ;
        RECT 75.930 108.110 76.220 108.340 ;
        RECT 78.330 108.110 78.620 108.340 ;
        RECT 79.280 108.290 79.600 108.350 ;
        RECT 82.640 108.290 82.960 108.350 ;
        RECT 87.050 108.340 87.190 108.520 ;
        RECT 79.080 108.150 79.600 108.290 ;
        RECT 25.530 107.740 25.820 107.970 ;
        RECT 26.480 107.920 26.800 107.980 ;
        RECT 26.280 107.780 26.800 107.920 ;
        RECT 26.480 107.720 26.800 107.780 ;
      LAYER met1 ;
        RECT 30.820 107.920 31.110 107.970 ;
        RECT 33.220 107.920 33.510 107.970 ;
        RECT 38.500 107.920 38.790 107.970 ;
        RECT 30.820 107.780 38.790 107.920 ;
        RECT 30.820 107.740 31.110 107.780 ;
        RECT 33.220 107.740 33.510 107.780 ;
        RECT 38.500 107.740 38.790 107.780 ;
        RECT 51.460 107.920 51.750 107.970 ;
        RECT 53.860 107.920 54.150 107.970 ;
        RECT 59.140 107.920 59.430 107.970 ;
        RECT 51.460 107.780 59.430 107.920 ;
        RECT 51.460 107.740 51.750 107.780 ;
        RECT 53.860 107.740 54.150 107.780 ;
        RECT 59.140 107.740 59.430 107.780 ;
      LAYER met1 ;
        RECT 65.360 107.920 65.680 107.980 ;
        RECT 70.650 107.920 70.940 107.970 ;
        RECT 65.360 107.780 70.940 107.920 ;
        RECT 65.360 107.720 65.680 107.780 ;
        RECT 70.650 107.740 70.940 107.780 ;
        RECT 74.010 107.740 74.300 107.970 ;
        RECT 75.450 107.740 75.740 107.970 ;
        RECT 78.410 107.920 78.550 108.110 ;
        RECT 79.280 108.090 79.600 108.150 ;
        RECT 79.850 108.150 82.960 108.290 ;
        RECT 79.850 107.920 79.990 108.150 ;
        RECT 82.640 108.090 82.960 108.150 ;
        RECT 86.970 108.110 87.260 108.340 ;
        RECT 87.920 108.290 88.240 108.350 ;
        RECT 87.720 108.150 88.240 108.290 ;
        RECT 88.490 108.290 88.630 108.890 ;
        RECT 107.120 108.890 114.160 109.030 ;
        RECT 107.120 108.830 107.440 108.890 ;
        RECT 112.410 108.850 112.700 108.890 ;
        RECT 113.840 108.830 114.160 108.890 ;
        RECT 117.210 109.030 117.500 109.080 ;
        RECT 118.160 109.030 118.480 109.090 ;
        RECT 117.210 108.890 118.480 109.030 ;
        RECT 117.210 108.850 117.500 108.890 ;
        RECT 118.160 108.830 118.480 108.890 ;
        RECT 91.760 108.660 92.080 108.720 ;
        RECT 107.610 108.660 107.900 108.710 ;
        RECT 108.560 108.660 108.880 108.720 ;
        RECT 123.920 108.660 124.240 108.720 ;
        RECT 91.760 108.520 99.190 108.660 ;
        RECT 91.760 108.460 92.080 108.520 ;
        RECT 99.050 108.340 99.190 108.520 ;
        RECT 107.610 108.520 108.880 108.660 ;
        RECT 123.720 108.520 124.240 108.660 ;
        RECT 107.610 108.480 107.900 108.520 ;
        RECT 108.560 108.460 108.880 108.520 ;
        RECT 123.920 108.460 124.240 108.520 ;
        RECT 92.250 108.290 92.540 108.340 ;
        RECT 88.490 108.150 92.540 108.290 ;
        RECT 87.920 108.090 88.240 108.150 ;
        RECT 92.250 108.110 92.540 108.150 ;
        RECT 98.970 108.110 99.260 108.340 ;
        RECT 109.040 108.290 109.360 108.350 ;
        RECT 113.850 108.290 114.140 108.340 ;
        RECT 109.040 108.150 114.140 108.290 ;
        RECT 109.040 108.090 109.360 108.150 ;
        RECT 113.850 108.110 114.140 108.150 ;
        RECT 80.720 107.920 81.040 107.980 ;
        RECT 81.680 107.920 82.000 107.980 ;
        RECT 85.520 107.920 85.840 107.980 ;
        RECT 78.410 107.780 79.990 107.920 ;
        RECT 80.520 107.780 81.040 107.920 ;
        RECT 81.480 107.780 82.000 107.920 ;
        RECT 85.320 107.780 85.840 107.920 ;
        RECT 61.520 107.180 61.840 107.240 ;
        RECT 74.090 107.180 74.230 107.740 ;
        RECT 75.530 107.550 75.670 107.740 ;
        RECT 80.720 107.720 81.040 107.780 ;
        RECT 81.680 107.720 82.000 107.780 ;
        RECT 85.520 107.720 85.840 107.780 ;
        RECT 86.000 107.920 86.320 107.980 ;
        RECT 86.490 107.920 86.780 107.970 ;
        RECT 86.000 107.780 86.780 107.920 ;
        RECT 86.000 107.720 86.320 107.780 ;
        RECT 86.490 107.740 86.780 107.780 ;
        RECT 94.640 107.920 94.960 107.980 ;
        RECT 96.090 107.920 96.380 107.970 ;
        RECT 100.400 107.920 100.720 107.980 ;
        RECT 94.640 107.780 100.720 107.920 ;
        RECT 94.640 107.720 94.960 107.780 ;
        RECT 96.090 107.740 96.380 107.780 ;
        RECT 100.400 107.720 100.720 107.780 ;
        RECT 102.320 107.920 102.640 107.980 ;
        RECT 102.810 107.920 103.100 107.970 ;
        RECT 102.320 107.780 103.100 107.920 ;
        RECT 102.320 107.720 102.640 107.780 ;
        RECT 102.810 107.740 103.100 107.780 ;
        RECT 103.280 107.920 103.600 107.980 ;
        RECT 109.530 107.920 109.820 107.970 ;
        RECT 125.370 107.920 125.660 107.970 ;
        RECT 103.280 107.780 109.820 107.920 ;
        RECT 103.280 107.720 103.600 107.780 ;
        RECT 109.530 107.740 109.820 107.780 ;
        RECT 118.730 107.780 125.660 107.920 ;
        RECT 85.040 107.550 85.360 107.610 ;
        RECT 75.530 107.410 85.360 107.550 ;
        RECT 85.040 107.350 85.360 107.410 ;
        RECT 84.090 107.180 84.380 107.230 ;
        RECT 86.480 107.180 86.800 107.240 ;
        RECT 61.520 107.040 74.230 107.180 ;
        RECT 78.890 107.040 83.830 107.180 ;
        RECT 61.520 106.980 61.840 107.040 ;
        RECT 13.040 106.810 13.360 106.870 ;
        RECT 24.570 106.810 24.860 106.860 ;
        RECT 13.040 106.670 24.860 106.810 ;
        RECT 13.040 106.610 13.360 106.670 ;
        RECT 24.570 106.630 24.860 106.670 ;
        RECT 47.130 106.810 47.420 106.860 ;
        RECT 55.280 106.810 55.600 106.870 ;
        RECT 47.130 106.670 55.600 106.810 ;
        RECT 47.130 106.630 47.420 106.670 ;
        RECT 55.280 106.610 55.600 106.670 ;
        RECT 72.080 106.810 72.400 106.870 ;
        RECT 78.890 106.810 79.030 107.040 ;
        RECT 79.760 106.810 80.080 106.870 ;
        RECT 72.080 106.670 79.030 106.810 ;
        RECT 79.560 106.670 80.080 106.810 ;
        RECT 83.690 106.810 83.830 107.040 ;
        RECT 84.090 107.040 86.800 107.180 ;
        RECT 84.090 107.000 84.380 107.040 ;
        RECT 86.480 106.980 86.800 107.040 ;
        RECT 109.040 106.810 109.360 106.870 ;
        RECT 83.690 106.670 109.360 106.810 ;
        RECT 72.080 106.610 72.400 106.670 ;
        RECT 79.760 106.610 80.080 106.670 ;
        RECT 109.040 106.610 109.360 106.670 ;
        RECT 117.680 106.810 118.000 106.870 ;
        RECT 118.730 106.860 118.870 107.780 ;
        RECT 125.370 107.740 125.660 107.780 ;
        RECT 118.650 106.810 118.940 106.860 ;
        RECT 117.680 106.670 118.940 106.810 ;
        RECT 117.680 106.610 118.000 106.670 ;
        RECT 118.650 106.630 118.940 106.670 ;
        RECT 26.480 104.960 26.800 105.020 ;
        RECT 27.930 104.960 28.220 105.010 ;
        RECT 26.480 104.820 28.220 104.960 ;
        RECT 26.480 104.760 26.800 104.820 ;
        RECT 27.930 104.780 28.220 104.820 ;
        RECT 31.290 104.960 31.580 105.010 ;
        RECT 32.240 104.960 32.560 105.020 ;
        RECT 31.290 104.820 32.560 104.960 ;
        RECT 31.290 104.780 31.580 104.820 ;
        RECT 32.240 104.760 32.560 104.820 ;
        RECT 33.210 104.960 33.500 105.010 ;
        RECT 37.520 104.960 37.840 105.020 ;
        RECT 33.210 104.820 37.840 104.960 ;
        RECT 33.210 104.780 33.500 104.820 ;
        RECT 37.520 104.760 37.840 104.820 ;
        RECT 61.520 104.960 61.840 105.020 ;
        RECT 62.490 104.960 62.780 105.010 ;
        RECT 61.520 104.820 62.780 104.960 ;
        RECT 61.520 104.760 61.840 104.820 ;
        RECT 62.490 104.780 62.780 104.820 ;
        RECT 79.770 104.960 80.060 105.010 ;
        RECT 85.520 104.960 85.840 105.020 ;
        RECT 79.770 104.820 85.840 104.960 ;
        RECT 79.770 104.780 80.060 104.820 ;
        RECT 85.520 104.760 85.840 104.820 ;
        RECT 98.000 104.960 98.320 105.020 ;
        RECT 98.490 104.960 98.780 105.010 ;
        RECT 98.000 104.820 98.780 104.960 ;
        RECT 98.000 104.760 98.320 104.820 ;
        RECT 98.490 104.780 98.780 104.820 ;
        RECT 117.680 104.220 118.000 104.280 ;
        RECT 135.930 104.220 136.220 104.270 ;
        RECT 66.410 104.080 136.220 104.220 ;
      LAYER met1 ;
        RECT 11.620 103.860 11.910 103.900 ;
        RECT 14.020 103.860 14.310 103.900 ;
        RECT 19.300 103.860 19.590 103.900 ;
        RECT 11.620 103.720 19.590 103.860 ;
      LAYER met1 ;
        RECT 43.760 103.850 44.080 103.910 ;
        RECT 44.720 103.850 45.040 103.910 ;
      LAYER met1 ;
        RECT 11.620 103.670 11.910 103.720 ;
        RECT 14.020 103.670 14.310 103.720 ;
        RECT 19.300 103.670 19.590 103.720 ;
      LAYER met1 ;
        RECT 36.170 103.710 44.080 103.850 ;
        RECT 44.520 103.710 45.040 103.850 ;
        RECT 13.040 103.480 13.360 103.540 ;
        RECT 36.170 103.530 36.310 103.710 ;
        RECT 43.760 103.650 44.080 103.710 ;
        RECT 44.720 103.650 45.040 103.710 ;
        RECT 51.450 103.850 51.740 103.900 ;
        RECT 52.400 103.850 52.720 103.910 ;
        RECT 58.170 103.850 58.460 103.900 ;
        RECT 51.450 103.710 52.720 103.850 ;
        RECT 51.450 103.670 51.740 103.710 ;
        RECT 52.400 103.650 52.720 103.710 ;
        RECT 57.770 103.710 58.460 103.850 ;
        RECT 12.840 103.340 13.360 103.480 ;
        RECT 13.040 103.280 13.360 103.340 ;
        RECT 24.570 103.480 24.860 103.530 ;
        RECT 27.450 103.480 27.740 103.530 ;
        RECT 34.170 103.480 34.460 103.530 ;
        RECT 24.570 103.340 34.460 103.480 ;
        RECT 24.570 103.300 24.860 103.340 ;
        RECT 27.450 103.300 27.740 103.340 ;
        RECT 34.170 103.300 34.460 103.340 ;
        RECT 36.090 103.300 36.380 103.530 ;
        RECT 40.880 103.480 41.200 103.540 ;
        RECT 54.320 103.480 54.640 103.540 ;
        RECT 40.680 103.340 41.200 103.480 ;
        RECT 54.120 103.340 54.640 103.480 ;
        RECT 40.880 103.280 41.200 103.340 ;
        RECT 54.320 103.280 54.640 103.340 ;
        RECT 21.200 103.110 21.520 103.170 ;
        RECT 21.000 102.970 21.520 103.110 ;
        RECT 21.200 102.910 21.520 102.970 ;
        RECT 50.010 103.110 50.300 103.160 ;
        RECT 57.200 103.110 57.520 103.170 ;
        RECT 57.770 103.110 57.910 103.710 ;
        RECT 58.170 103.670 58.460 103.710 ;
        RECT 66.410 103.480 66.550 104.080 ;
        RECT 117.680 104.020 118.000 104.080 ;
        RECT 135.930 104.040 136.220 104.080 ;
      LAYER met1 ;
        RECT 66.820 103.860 67.110 103.900 ;
        RECT 69.220 103.860 69.510 103.900 ;
        RECT 74.500 103.860 74.790 103.900 ;
        RECT 66.820 103.720 74.790 103.860 ;
        RECT 66.820 103.670 67.110 103.720 ;
        RECT 69.220 103.670 69.510 103.720 ;
        RECT 74.500 103.670 74.790 103.720 ;
      LAYER met1 ;
        RECT 85.040 103.850 85.360 103.910 ;
        RECT 86.010 103.850 86.300 103.900 ;
        RECT 92.720 103.850 93.040 103.910 ;
        RECT 85.040 103.710 86.300 103.850 ;
        RECT 92.520 103.710 93.040 103.850 ;
        RECT 85.040 103.650 85.360 103.710 ;
        RECT 86.010 103.670 86.300 103.710 ;
        RECT 92.720 103.650 93.040 103.710 ;
        RECT 94.160 103.850 94.480 103.910 ;
        RECT 99.930 103.850 100.220 103.900 ;
        RECT 109.520 103.850 109.840 103.910 ;
        RECT 94.160 103.710 100.220 103.850 ;
        RECT 109.320 103.710 109.840 103.850 ;
        RECT 94.160 103.650 94.480 103.710 ;
        RECT 99.930 103.670 100.220 103.710 ;
        RECT 109.520 103.650 109.840 103.710 ;
        RECT 116.250 103.850 116.540 103.900 ;
        RECT 117.200 103.850 117.520 103.910 ;
        RECT 125.360 103.850 125.680 103.910 ;
        RECT 116.250 103.710 117.520 103.850 ;
        RECT 125.160 103.710 125.680 103.850 ;
        RECT 116.250 103.670 116.540 103.710 ;
        RECT 117.200 103.650 117.520 103.710 ;
        RECT 125.360 103.650 125.680 103.710 ;
        RECT 63.530 103.340 66.550 103.480 ;
        RECT 68.250 103.480 68.540 103.530 ;
        RECT 79.760 103.480 80.080 103.540 ;
        RECT 82.160 103.480 82.480 103.540 ;
        RECT 68.250 103.340 80.080 103.480 ;
        RECT 81.960 103.340 82.480 103.480 ;
        RECT 58.160 103.110 58.480 103.170 ;
        RECT 63.530 103.110 63.670 103.340 ;
        RECT 68.250 103.300 68.540 103.340 ;
        RECT 79.760 103.280 80.080 103.340 ;
        RECT 82.160 103.280 82.480 103.340 ;
        RECT 85.520 103.480 85.840 103.540 ;
        RECT 88.890 103.480 89.180 103.530 ;
        RECT 85.520 103.340 89.180 103.480 ;
        RECT 85.520 103.280 85.840 103.340 ;
        RECT 88.890 103.300 89.180 103.340 ;
        RECT 101.360 103.480 101.680 103.540 ;
        RECT 102.320 103.480 102.640 103.540 ;
        RECT 105.680 103.480 106.000 103.540 ;
        RECT 101.360 103.340 101.880 103.480 ;
        RECT 102.120 103.340 102.640 103.480 ;
        RECT 105.480 103.340 106.000 103.480 ;
        RECT 101.360 103.280 101.680 103.340 ;
        RECT 102.320 103.280 102.640 103.340 ;
        RECT 105.680 103.280 106.000 103.340 ;
        RECT 111.440 103.480 111.760 103.540 ;
        RECT 112.410 103.480 112.700 103.530 ;
        RECT 111.440 103.340 112.700 103.480 ;
        RECT 111.440 103.280 111.760 103.340 ;
        RECT 112.410 103.300 112.700 103.340 ;
        RECT 65.360 103.110 65.680 103.170 ;
        RECT 76.400 103.110 76.720 103.170 ;
        RECT 50.010 102.970 57.520 103.110 ;
        RECT 57.720 102.970 63.670 103.110 ;
        RECT 65.160 102.970 65.680 103.110 ;
        RECT 76.200 102.970 76.720 103.110 ;
        RECT 50.010 102.930 50.300 102.970 ;
        RECT 57.200 102.910 57.520 102.970 ;
        RECT 58.160 102.910 58.480 102.970 ;
        RECT 65.360 102.910 65.680 102.970 ;
        RECT 76.400 102.910 76.720 102.970 ;
        RECT 123.930 103.110 124.220 103.160 ;
        RECT 124.880 103.110 125.200 103.170 ;
        RECT 123.930 102.970 125.200 103.110 ;
        RECT 123.930 102.930 124.220 102.970 ;
        RECT 124.880 102.910 125.200 102.970 ;
        RECT 5.760 102.010 142.080 102.380 ;
        RECT 16.410 100.890 16.700 100.940 ;
        RECT 21.200 100.890 21.520 100.950 ;
        RECT 16.410 100.750 21.520 100.890 ;
        RECT 16.410 100.710 16.700 100.750 ;
        RECT 21.200 100.690 21.520 100.750 ;
        RECT 65.360 100.890 65.680 100.950 ;
        RECT 66.810 100.890 67.100 100.940 ;
        RECT 65.360 100.750 67.100 100.890 ;
        RECT 65.360 100.690 65.680 100.750 ;
        RECT 66.810 100.710 67.100 100.750 ;
        RECT 78.320 100.890 78.640 100.950 ;
        RECT 81.200 100.890 81.520 100.950 ;
        RECT 78.320 100.750 81.520 100.890 ;
        RECT 78.320 100.690 78.640 100.750 ;
        RECT 81.200 100.690 81.520 100.750 ;
        RECT 83.120 100.890 83.440 100.950 ;
        RECT 83.120 100.750 85.270 100.890 ;
        RECT 83.120 100.690 83.440 100.750 ;
        RECT 31.760 100.520 32.080 100.580 ;
        RECT 32.250 100.520 32.540 100.570 ;
        RECT 43.280 100.520 43.600 100.580 ;
        RECT 31.760 100.380 32.540 100.520 ;
        RECT 43.080 100.380 43.600 100.520 ;
        RECT 31.760 100.320 32.080 100.380 ;
        RECT 32.250 100.340 32.540 100.380 ;
        RECT 43.280 100.320 43.600 100.380 ;
        RECT 50.010 100.520 50.300 100.570 ;
        RECT 53.840 100.520 54.160 100.580 ;
        RECT 74.960 100.520 75.280 100.580 ;
        RECT 85.130 100.520 85.270 100.750 ;
        RECT 99.930 100.520 100.220 100.570 ;
        RECT 100.880 100.520 101.200 100.580 ;
        RECT 50.010 100.380 54.160 100.520 ;
        RECT 74.760 100.380 75.280 100.520 ;
        RECT 50.010 100.340 50.300 100.380 ;
        RECT 53.840 100.320 54.160 100.380 ;
        RECT 74.960 100.320 75.280 100.380 ;
        RECT 78.410 100.380 84.790 100.520 ;
        RECT 85.130 100.380 93.430 100.520 ;
        RECT 22.160 100.150 22.480 100.210 ;
        RECT 21.960 100.010 22.480 100.150 ;
        RECT 22.160 99.950 22.480 100.010 ;
        RECT 29.370 99.970 29.660 100.200 ;
        RECT 33.680 100.150 34.000 100.210 ;
        RECT 52.400 100.150 52.720 100.210 ;
        RECT 54.330 100.150 54.620 100.200 ;
        RECT 33.480 100.010 34.000 100.150 ;
        RECT 29.450 99.780 29.590 99.970 ;
        RECT 33.680 99.950 34.000 100.010 ;
        RECT 44.330 100.010 51.670 100.150 ;
        RECT 44.330 99.780 44.470 100.010 ;
        RECT 51.530 99.830 51.670 100.010 ;
        RECT 52.400 100.010 54.620 100.150 ;
        RECT 52.400 99.950 52.720 100.010 ;
        RECT 54.330 99.970 54.620 100.010 ;
        RECT 56.720 100.150 57.040 100.210 ;
        RECT 61.040 100.150 61.360 100.210 ;
        RECT 62.000 100.150 62.320 100.210 ;
        RECT 75.440 100.150 75.760 100.210 ;
        RECT 56.720 100.010 58.390 100.150 ;
        RECT 60.840 100.010 61.360 100.150 ;
        RECT 61.800 100.010 62.320 100.150 ;
        RECT 56.720 99.950 57.040 100.010 ;
        RECT 29.450 99.640 44.470 99.780 ;
        RECT 44.730 99.600 45.020 99.830 ;
        RECT 51.450 99.780 51.740 99.830 ;
        RECT 57.680 99.780 58.000 99.840 ;
        RECT 58.250 99.830 58.390 100.010 ;
        RECT 61.040 99.950 61.360 100.010 ;
        RECT 62.000 99.950 62.320 100.010 ;
        RECT 74.090 100.010 75.760 100.150 ;
        RECT 51.450 99.640 58.000 99.780 ;
        RECT 51.450 99.600 51.740 99.640 ;
        RECT 44.810 99.410 44.950 99.600 ;
        RECT 57.680 99.580 58.000 99.640 ;
        RECT 58.170 99.600 58.460 99.830 ;
        RECT 62.480 99.780 62.800 99.840 ;
        RECT 62.280 99.640 62.800 99.780 ;
        RECT 62.480 99.580 62.800 99.640 ;
        RECT 63.450 99.600 63.740 99.830 ;
        RECT 64.410 99.780 64.700 99.830 ;
        RECT 68.720 99.780 69.040 99.840 ;
        RECT 72.560 99.780 72.880 99.840 ;
        RECT 74.090 99.830 74.230 100.010 ;
        RECT 75.440 99.950 75.760 100.010 ;
        RECT 64.410 99.640 69.040 99.780 ;
        RECT 72.360 99.640 72.880 99.780 ;
        RECT 64.410 99.600 64.700 99.640 ;
        RECT 54.320 99.410 54.640 99.470 ;
        RECT 44.810 99.270 54.640 99.410 ;
        RECT 54.320 99.210 54.640 99.270 ;
        RECT 57.200 99.410 57.520 99.470 ;
        RECT 63.530 99.410 63.670 99.600 ;
        RECT 68.720 99.580 69.040 99.640 ;
        RECT 72.560 99.580 72.880 99.640 ;
        RECT 74.010 99.600 74.300 99.830 ;
        RECT 74.490 99.780 74.780 99.830 ;
        RECT 78.410 99.780 78.550 100.380 ;
        RECT 84.650 100.200 84.790 100.380 ;
        RECT 93.290 100.200 93.430 100.380 ;
        RECT 99.930 100.380 101.200 100.520 ;
        RECT 99.930 100.340 100.220 100.380 ;
        RECT 100.880 100.320 101.200 100.380 ;
        RECT 102.320 100.520 102.640 100.580 ;
        RECT 110.960 100.520 111.280 100.580 ;
        RECT 102.320 100.380 111.280 100.520 ;
        RECT 102.320 100.320 102.640 100.380 ;
        RECT 78.810 100.150 79.100 100.200 ;
        RECT 78.810 100.010 83.350 100.150 ;
        RECT 78.810 99.970 79.100 100.010 ;
        RECT 74.490 99.640 78.550 99.780 ;
        RECT 74.490 99.600 74.780 99.640 ;
        RECT 81.690 99.600 81.980 99.830 ;
        RECT 83.210 99.780 83.350 100.010 ;
        RECT 84.570 99.970 84.860 100.200 ;
        RECT 93.210 99.970 93.500 100.200 ;
        RECT 101.360 100.150 101.680 100.210 ;
        RECT 103.370 100.200 103.510 100.380 ;
        RECT 110.960 100.320 111.280 100.380 ;
        RECT 102.810 100.150 103.100 100.200 ;
        RECT 101.360 100.010 103.100 100.150 ;
        RECT 101.360 99.950 101.680 100.010 ;
        RECT 102.810 99.970 103.100 100.010 ;
        RECT 103.290 99.970 103.580 100.200 ;
        RECT 104.240 100.150 104.560 100.210 ;
        RECT 104.040 100.010 104.560 100.150 ;
        RECT 104.240 99.950 104.560 100.010 ;
        RECT 107.600 100.150 107.920 100.210 ;
        RECT 108.570 100.150 108.860 100.200 ;
        RECT 113.840 100.150 114.160 100.210 ;
        RECT 107.600 100.010 108.860 100.150 ;
        RECT 113.640 100.010 114.160 100.150 ;
        RECT 107.600 99.950 107.920 100.010 ;
        RECT 108.570 99.970 108.860 100.010 ;
        RECT 113.840 99.950 114.160 100.010 ;
        RECT 118.160 100.150 118.480 100.210 ;
        RECT 118.650 100.150 118.940 100.200 ;
        RECT 118.160 100.010 118.940 100.150 ;
        RECT 118.160 99.950 118.480 100.010 ;
        RECT 118.650 99.970 118.940 100.010 ;
        RECT 125.360 100.150 125.680 100.210 ;
        RECT 128.250 100.150 128.540 100.200 ;
        RECT 125.360 100.010 128.540 100.150 ;
        RECT 125.360 99.950 125.680 100.010 ;
        RECT 128.250 99.970 128.540 100.010 ;
        RECT 88.410 99.780 88.700 99.830 ;
        RECT 83.210 99.640 88.700 99.780 ;
        RECT 88.410 99.600 88.700 99.640 ;
        RECT 97.050 99.780 97.340 99.830 ;
        RECT 101.840 99.780 102.160 99.840 ;
        RECT 97.050 99.640 102.160 99.780 ;
        RECT 97.050 99.600 97.340 99.640 ;
        RECT 57.200 99.270 63.670 99.410 ;
        RECT 67.280 99.410 67.600 99.470 ;
        RECT 81.770 99.410 81.910 99.600 ;
        RECT 101.840 99.580 102.160 99.640 ;
        RECT 123.920 99.780 124.240 99.840 ;
        RECT 132.090 99.780 132.380 99.830 ;
        RECT 123.920 99.640 132.380 99.780 ;
        RECT 123.920 99.580 124.240 99.640 ;
        RECT 132.090 99.600 132.380 99.640 ;
        RECT 93.200 99.410 93.520 99.470 ;
        RECT 67.280 99.270 93.520 99.410 ;
        RECT 57.200 99.210 57.520 99.270 ;
        RECT 67.280 99.210 67.600 99.270 ;
        RECT 93.200 99.210 93.520 99.270 ;
        RECT 111.930 99.410 112.220 99.460 ;
        RECT 116.720 99.410 117.040 99.470 ;
        RECT 111.930 99.270 117.040 99.410 ;
        RECT 111.930 99.230 112.220 99.270 ;
        RECT 116.720 99.210 117.040 99.270 ;
        RECT 38.010 99.040 38.300 99.090 ;
        RECT 58.160 99.040 58.480 99.100 ;
        RECT 38.010 98.900 58.480 99.040 ;
        RECT 38.010 98.860 38.300 98.900 ;
        RECT 58.160 98.840 58.480 98.900 ;
        RECT 100.400 99.040 100.720 99.100 ;
        RECT 107.130 99.040 107.420 99.090 ;
        RECT 117.200 99.040 117.520 99.100 ;
        RECT 100.400 98.900 107.420 99.040 ;
        RECT 100.400 98.840 100.720 98.900 ;
        RECT 107.130 98.860 107.420 98.900 ;
        RECT 107.690 98.900 117.520 99.040 ;
        RECT 14.480 98.670 14.800 98.730 ;
        RECT 17.850 98.670 18.140 98.720 ;
        RECT 23.120 98.670 23.440 98.730 ;
        RECT 14.480 98.530 18.140 98.670 ;
        RECT 22.920 98.530 23.440 98.670 ;
        RECT 14.480 98.470 14.800 98.530 ;
        RECT 17.850 98.490 18.140 98.530 ;
        RECT 23.120 98.470 23.440 98.530 ;
        RECT 29.850 98.670 30.140 98.720 ;
        RECT 30.320 98.670 30.640 98.730 ;
        RECT 29.850 98.530 30.640 98.670 ;
        RECT 29.850 98.490 30.140 98.530 ;
        RECT 30.320 98.470 30.640 98.530 ;
        RECT 36.570 98.670 36.860 98.720 ;
        RECT 54.800 98.670 55.120 98.730 ;
        RECT 36.570 98.530 55.120 98.670 ;
        RECT 36.570 98.490 36.860 98.530 ;
        RECT 54.800 98.470 55.120 98.530 ;
        RECT 68.250 98.670 68.540 98.720 ;
        RECT 69.200 98.670 69.520 98.730 ;
        RECT 107.690 98.670 107.830 98.900 ;
        RECT 117.200 98.840 117.520 98.900 ;
        RECT 68.250 98.530 107.830 98.670 ;
        RECT 68.250 98.490 68.540 98.530 ;
        RECT 69.200 98.470 69.520 98.530 ;
        RECT 20.730 96.820 21.020 96.870 ;
        RECT 22.160 96.820 22.480 96.880 ;
        RECT 20.730 96.680 22.480 96.820 ;
        RECT 20.730 96.640 21.020 96.680 ;
        RECT 22.160 96.620 22.480 96.680 ;
        RECT 33.680 96.820 34.000 96.880 ;
        RECT 34.650 96.820 34.940 96.870 ;
        RECT 33.680 96.680 34.940 96.820 ;
        RECT 33.680 96.620 34.000 96.680 ;
        RECT 34.650 96.640 34.940 96.680 ;
        RECT 37.530 96.820 37.820 96.870 ;
        RECT 43.760 96.820 44.080 96.880 ;
        RECT 37.530 96.680 44.080 96.820 ;
        RECT 37.530 96.640 37.820 96.680 ;
        RECT 43.760 96.620 44.080 96.680 ;
        RECT 54.800 96.820 55.120 96.880 ;
        RECT 63.450 96.820 63.740 96.870 ;
        RECT 66.320 96.820 66.640 96.880 ;
        RECT 67.280 96.820 67.600 96.880 ;
        RECT 54.800 96.680 57.910 96.820 ;
        RECT 54.800 96.620 55.120 96.680 ;
        RECT 30.320 96.450 30.640 96.510 ;
        RECT 38.970 96.450 39.260 96.500 ;
        RECT 56.720 96.450 57.040 96.510 ;
        RECT 30.320 96.310 57.040 96.450 ;
        RECT 57.770 96.450 57.910 96.680 ;
        RECT 63.450 96.680 66.640 96.820 ;
        RECT 67.080 96.680 67.600 96.820 ;
        RECT 63.450 96.640 63.740 96.680 ;
        RECT 66.320 96.620 66.640 96.680 ;
        RECT 67.280 96.620 67.600 96.680 ;
        RECT 69.690 96.820 69.980 96.870 ;
        RECT 76.400 96.820 76.720 96.880 ;
        RECT 69.690 96.680 76.720 96.820 ;
        RECT 69.690 96.640 69.980 96.680 ;
        RECT 76.400 96.620 76.720 96.680 ;
        RECT 95.610 96.820 95.900 96.870 ;
        RECT 101.360 96.820 101.680 96.880 ;
        RECT 103.280 96.820 103.600 96.880 ;
        RECT 95.610 96.680 103.600 96.820 ;
        RECT 95.610 96.640 95.900 96.680 ;
        RECT 101.360 96.620 101.680 96.680 ;
        RECT 103.280 96.620 103.600 96.680 ;
        RECT 104.240 96.820 104.560 96.880 ;
        RECT 114.330 96.820 114.620 96.870 ;
        RECT 116.720 96.820 117.040 96.880 ;
        RECT 104.240 96.680 114.620 96.820 ;
        RECT 116.520 96.680 117.040 96.820 ;
        RECT 104.240 96.620 104.560 96.680 ;
        RECT 114.330 96.640 114.620 96.680 ;
        RECT 116.720 96.620 117.040 96.680 ;
        RECT 117.200 96.820 117.520 96.880 ;
        RECT 118.170 96.820 118.460 96.870 ;
        RECT 117.200 96.680 118.460 96.820 ;
        RECT 117.200 96.620 117.520 96.680 ;
        RECT 118.170 96.640 118.460 96.680 ;
        RECT 64.400 96.450 64.720 96.510 ;
        RECT 71.130 96.450 71.420 96.500 ;
        RECT 57.770 96.310 71.420 96.450 ;
        RECT 30.320 96.250 30.640 96.310 ;
        RECT 38.970 96.270 39.260 96.310 ;
        RECT 56.720 96.250 57.040 96.310 ;
        RECT 64.400 96.250 64.720 96.310 ;
        RECT 71.130 96.270 71.420 96.310 ;
        RECT 75.930 96.450 76.220 96.500 ;
        RECT 86.000 96.450 86.320 96.510 ;
        RECT 89.840 96.450 90.160 96.510 ;
        RECT 75.930 96.310 86.320 96.450 ;
        RECT 75.930 96.270 76.220 96.310 ;
        RECT 86.000 96.250 86.320 96.310 ;
        RECT 86.570 96.310 90.160 96.450 ;
        RECT 23.120 96.080 23.440 96.140 ;
        RECT 61.040 96.080 61.360 96.140 ;
        RECT 23.120 95.940 61.360 96.080 ;
        RECT 23.120 95.880 23.440 95.940 ;
      LAYER met1 ;
        RECT 7.780 95.720 8.070 95.760 ;
        RECT 10.180 95.720 10.470 95.760 ;
        RECT 15.460 95.720 15.750 95.760 ;
        RECT 7.780 95.580 15.750 95.720 ;
        RECT 7.780 95.530 8.070 95.580 ;
        RECT 10.180 95.530 10.470 95.580 ;
        RECT 15.460 95.530 15.750 95.580 ;
      LAYER met1 ;
        RECT 24.080 95.710 24.400 95.770 ;
        RECT 26.960 95.710 27.280 95.770 ;
        RECT 28.010 95.760 28.150 95.940 ;
        RECT 61.040 95.880 61.360 95.940 ;
        RECT 74.010 96.080 74.300 96.130 ;
        RECT 86.570 96.080 86.710 96.310 ;
        RECT 89.840 96.250 90.160 96.310 ;
        RECT 74.010 95.940 86.710 96.080 ;
        RECT 86.960 96.080 87.280 96.140 ;
        RECT 86.960 95.940 112.630 96.080 ;
        RECT 74.010 95.900 74.300 95.940 ;
        RECT 27.450 95.710 27.740 95.760 ;
        RECT 24.080 95.570 26.230 95.710 ;
        RECT 24.080 95.510 24.400 95.570 ;
        RECT 25.050 95.340 25.340 95.390 ;
        RECT 25.520 95.340 25.840 95.400 ;
        RECT 26.090 95.390 26.230 95.570 ;
        RECT 26.960 95.570 27.740 95.710 ;
        RECT 26.960 95.510 27.280 95.570 ;
        RECT 27.450 95.530 27.740 95.570 ;
        RECT 27.930 95.530 28.220 95.760 ;
        RECT 43.280 95.710 43.600 95.770 ;
        RECT 45.690 95.710 45.980 95.760 ;
        RECT 52.400 95.710 52.720 95.770 ;
        RECT 43.280 95.570 45.980 95.710 ;
        RECT 52.200 95.570 52.720 95.710 ;
        RECT 43.280 95.510 43.600 95.570 ;
        RECT 45.690 95.530 45.980 95.570 ;
        RECT 52.400 95.510 52.720 95.570 ;
        RECT 52.880 95.710 53.200 95.770 ;
        RECT 57.680 95.710 58.000 95.770 ;
        RECT 77.450 95.760 77.590 95.940 ;
        RECT 86.960 95.880 87.280 95.940 ;
        RECT 59.130 95.710 59.420 95.760 ;
        RECT 52.880 95.570 55.510 95.710 ;
        RECT 52.880 95.510 53.200 95.570 ;
        RECT 25.050 95.200 25.840 95.340 ;
        RECT 25.050 95.160 25.340 95.200 ;
        RECT 25.520 95.140 25.840 95.200 ;
        RECT 26.010 95.340 26.300 95.390 ;
        RECT 28.400 95.340 28.720 95.400 ;
        RECT 26.010 95.200 28.720 95.340 ;
        RECT 26.010 95.160 26.300 95.200 ;
        RECT 28.400 95.140 28.720 95.200 ;
        RECT 36.560 95.340 36.880 95.400 ;
        RECT 55.370 95.390 55.510 95.570 ;
        RECT 57.680 95.570 75.670 95.710 ;
        RECT 57.680 95.510 58.000 95.570 ;
        RECT 59.130 95.530 59.420 95.570 ;
        RECT 41.850 95.340 42.140 95.390 ;
        RECT 36.560 95.200 42.140 95.340 ;
        RECT 36.560 95.140 36.880 95.200 ;
        RECT 41.850 95.160 42.140 95.200 ;
        RECT 55.290 95.160 55.580 95.390 ;
        RECT 66.810 95.340 67.100 95.390 ;
        RECT 72.080 95.340 72.400 95.400 ;
        RECT 66.810 95.200 72.400 95.340 ;
        RECT 66.810 95.160 67.100 95.200 ;
        RECT 72.080 95.140 72.400 95.200 ;
        RECT 74.970 95.160 75.260 95.390 ;
        RECT 50.970 94.970 51.260 95.020 ;
        RECT 52.880 94.970 53.200 95.030 ;
        RECT 50.970 94.830 53.200 94.970 ;
        RECT 50.970 94.790 51.260 94.830 ;
        RECT 52.880 94.770 53.200 94.830 ;
        RECT 57.200 94.970 57.520 95.030 ;
        RECT 74.010 94.970 74.300 95.020 ;
        RECT 57.200 94.830 74.300 94.970 ;
        RECT 57.200 94.770 57.520 94.830 ;
        RECT 74.010 94.790 74.300 94.830 ;
        RECT 8.720 94.600 9.040 94.660 ;
        RECT 8.520 94.460 9.040 94.600 ;
        RECT 8.720 94.400 9.040 94.460 ;
        RECT 9.210 94.600 9.500 94.650 ;
        RECT 26.010 94.600 26.300 94.650 ;
        RECT 9.210 94.460 26.300 94.600 ;
        RECT 9.210 94.420 9.500 94.460 ;
        RECT 26.010 94.420 26.300 94.460 ;
        RECT 33.210 94.600 33.500 94.650 ;
        RECT 36.080 94.600 36.400 94.660 ;
        RECT 62.000 94.600 62.320 94.660 ;
        RECT 33.210 94.460 36.400 94.600 ;
        RECT 61.800 94.460 62.320 94.600 ;
        RECT 75.050 94.600 75.190 95.160 ;
        RECT 75.530 94.970 75.670 95.570 ;
        RECT 77.370 95.530 77.660 95.760 ;
        RECT 83.610 95.710 83.900 95.760 ;
        RECT 90.320 95.710 90.640 95.770 ;
        RECT 93.200 95.710 93.520 95.770 ;
        RECT 83.610 95.570 86.230 95.710 ;
        RECT 90.120 95.570 90.640 95.710 ;
        RECT 93.000 95.570 93.520 95.710 ;
        RECT 83.610 95.530 83.900 95.570 ;
        RECT 75.930 95.340 76.220 95.390 ;
        RECT 79.280 95.340 79.600 95.400 ;
        RECT 75.930 95.200 79.600 95.340 ;
        RECT 75.930 95.160 76.220 95.200 ;
        RECT 79.280 95.140 79.600 95.200 ;
        RECT 78.800 94.970 79.120 95.030 ;
        RECT 81.200 94.970 81.520 95.030 ;
        RECT 75.530 94.830 79.120 94.970 ;
        RECT 81.000 94.830 81.520 94.970 ;
        RECT 78.800 94.770 79.120 94.830 ;
        RECT 81.200 94.770 81.520 94.830 ;
        RECT 84.080 94.600 84.400 94.660 ;
        RECT 75.050 94.460 84.400 94.600 ;
        RECT 86.090 94.600 86.230 95.570 ;
        RECT 90.320 95.510 90.640 95.570 ;
        RECT 93.200 95.510 93.520 95.570 ;
        RECT 93.690 95.530 93.980 95.760 ;
        RECT 95.130 95.530 95.420 95.760 ;
        RECT 102.810 95.710 103.100 95.760 ;
        RECT 108.080 95.710 108.400 95.770 ;
        RECT 102.810 95.570 108.400 95.710 ;
        RECT 102.810 95.530 103.100 95.570 ;
        RECT 86.480 95.340 86.800 95.400 ;
        RECT 93.770 95.340 93.910 95.530 ;
        RECT 86.480 95.200 93.910 95.340 ;
        RECT 86.480 95.140 86.800 95.200 ;
        RECT 87.920 94.970 88.240 95.030 ;
        RECT 87.720 94.830 88.240 94.970 ;
        RECT 87.920 94.770 88.240 94.830 ;
        RECT 93.200 94.970 93.520 95.030 ;
        RECT 95.210 94.970 95.350 95.530 ;
        RECT 108.080 95.510 108.400 95.570 ;
        RECT 108.560 95.710 108.880 95.770 ;
        RECT 112.490 95.760 112.630 95.940 ;
        RECT 109.530 95.710 109.820 95.760 ;
        RECT 108.560 95.570 109.820 95.710 ;
        RECT 108.560 95.510 108.880 95.570 ;
        RECT 109.530 95.530 109.820 95.570 ;
        RECT 112.410 95.530 112.700 95.760 ;
        RECT 113.850 95.530 114.140 95.760 ;
        RECT 123.920 95.710 124.240 95.770 ;
        RECT 125.370 95.710 125.660 95.760 ;
        RECT 123.920 95.570 125.660 95.710 ;
        RECT 107.600 95.340 107.920 95.400 ;
        RECT 113.930 95.340 114.070 95.530 ;
        RECT 123.920 95.510 124.240 95.570 ;
        RECT 125.370 95.530 125.660 95.570 ;
        RECT 107.600 95.200 114.070 95.340 ;
        RECT 107.600 95.140 107.920 95.200 ;
        RECT 100.880 94.970 101.200 95.030 ;
        RECT 93.200 94.830 95.350 94.970 ;
        RECT 100.680 94.830 101.200 94.970 ;
        RECT 93.200 94.770 93.520 94.830 ;
        RECT 100.880 94.770 101.200 94.830 ;
        RECT 108.090 94.970 108.380 95.020 ;
        RECT 109.520 94.970 109.840 95.030 ;
        RECT 108.090 94.830 109.840 94.970 ;
        RECT 108.090 94.790 108.380 94.830 ;
        RECT 109.520 94.770 109.840 94.830 ;
        RECT 123.930 94.970 124.220 95.020 ;
        RECT 132.080 94.970 132.400 95.030 ;
        RECT 123.930 94.830 132.400 94.970 ;
        RECT 123.930 94.790 124.220 94.830 ;
        RECT 132.080 94.770 132.400 94.830 ;
        RECT 93.290 94.600 93.430 94.770 ;
        RECT 86.090 94.460 93.430 94.600 ;
        RECT 33.210 94.420 33.500 94.460 ;
        RECT 36.080 94.400 36.400 94.460 ;
        RECT 62.000 94.400 62.320 94.460 ;
        RECT 84.080 94.400 84.400 94.460 ;
        RECT 5.760 93.870 142.080 94.240 ;
        RECT 8.720 92.750 9.040 92.810 ;
        RECT 13.050 92.750 13.340 92.800 ;
        RECT 8.720 92.610 13.340 92.750 ;
        RECT 8.720 92.550 9.040 92.610 ;
        RECT 13.050 92.570 13.340 92.610 ;
        RECT 21.680 92.750 22.000 92.810 ;
        RECT 28.410 92.750 28.700 92.800 ;
        RECT 21.680 92.610 28.700 92.750 ;
        RECT 21.680 92.550 22.000 92.610 ;
        RECT 28.410 92.570 28.700 92.610 ;
        RECT 36.080 92.750 36.400 92.810 ;
        RECT 45.690 92.750 45.980 92.800 ;
        RECT 92.720 92.750 93.040 92.810 ;
        RECT 36.080 92.610 45.980 92.750 ;
        RECT 36.080 92.550 36.400 92.610 ;
        RECT 45.690 92.570 45.980 92.610 ;
        RECT 77.450 92.610 93.040 92.750 ;
        RECT 25.050 92.380 25.340 92.430 ;
        RECT 25.520 92.380 25.840 92.440 ;
        RECT 57.210 92.380 57.500 92.430 ;
        RECT 62.000 92.380 62.320 92.440 ;
        RECT 77.450 92.430 77.590 92.610 ;
        RECT 92.720 92.550 93.040 92.610 ;
        RECT 101.840 92.750 102.160 92.810 ;
        RECT 107.120 92.750 107.440 92.810 ;
        RECT 110.960 92.750 111.280 92.810 ;
        RECT 101.840 92.610 110.230 92.750 ;
        RECT 110.760 92.610 111.280 92.750 ;
        RECT 101.840 92.550 102.160 92.610 ;
        RECT 107.120 92.550 107.440 92.610 ;
        RECT 25.050 92.240 30.550 92.380 ;
        RECT 25.050 92.200 25.340 92.240 ;
        RECT 25.520 92.180 25.840 92.240 ;
        RECT 24.080 92.010 24.400 92.070 ;
        RECT 27.450 92.010 27.740 92.060 ;
        RECT 28.400 92.010 28.720 92.070 ;
        RECT 23.880 91.870 24.400 92.010 ;
        RECT 24.080 91.810 24.400 91.870 ;
        RECT 26.570 91.870 27.740 92.010 ;
        RECT 28.200 91.870 28.720 92.010 ;
        RECT 26.570 91.270 26.710 91.870 ;
        RECT 27.450 91.830 27.740 91.870 ;
        RECT 28.400 91.810 28.720 91.870 ;
        RECT 26.960 91.640 27.280 91.700 ;
        RECT 30.410 91.690 30.550 92.240 ;
        RECT 57.210 92.240 62.320 92.380 ;
        RECT 57.210 92.200 57.500 92.240 ;
        RECT 62.000 92.180 62.320 92.240 ;
        RECT 77.370 92.200 77.660 92.430 ;
        RECT 84.090 92.380 84.380 92.430 ;
        RECT 90.320 92.380 90.640 92.440 ;
        RECT 84.090 92.240 90.640 92.380 ;
        RECT 84.090 92.200 84.380 92.240 ;
        RECT 90.320 92.180 90.640 92.240 ;
        RECT 97.050 92.380 97.340 92.430 ;
        RECT 97.050 92.240 109.750 92.380 ;
        RECT 97.050 92.200 97.340 92.240 ;
        RECT 39.930 92.010 40.220 92.060 ;
        RECT 53.360 92.010 53.680 92.070 ;
        RECT 39.930 91.870 53.680 92.010 ;
        RECT 39.930 91.830 40.220 91.870 ;
        RECT 53.360 91.810 53.680 91.870 ;
        RECT 57.680 92.010 58.000 92.070 ;
        RECT 60.090 92.010 60.380 92.060 ;
        RECT 57.680 91.870 60.380 92.010 ;
        RECT 57.680 91.810 58.000 91.870 ;
        RECT 60.090 91.830 60.380 91.870 ;
        RECT 79.280 92.010 79.600 92.070 ;
        RECT 88.410 92.010 88.700 92.060 ;
        RECT 79.280 91.870 88.700 92.010 ;
        RECT 79.280 91.810 79.600 91.870 ;
        RECT 88.410 91.830 88.700 91.870 ;
        RECT 97.520 92.010 97.840 92.070 ;
        RECT 101.850 92.010 102.140 92.060 ;
        RECT 97.520 91.870 102.140 92.010 ;
        RECT 97.520 91.810 97.840 91.870 ;
        RECT 101.850 91.830 102.140 91.870 ;
        RECT 102.320 92.010 102.640 92.070 ;
        RECT 109.610 92.060 109.750 92.240 ;
        RECT 108.570 92.010 108.860 92.060 ;
        RECT 102.320 91.870 108.860 92.010 ;
        RECT 102.320 91.810 102.640 91.870 ;
        RECT 108.570 91.830 108.860 91.870 ;
        RECT 109.530 91.830 109.820 92.060 ;
        RECT 110.090 92.010 110.230 92.610 ;
        RECT 110.960 92.550 111.280 92.610 ;
        RECT 123.920 92.380 124.240 92.440 ;
        RECT 123.720 92.240 124.240 92.380 ;
        RECT 123.920 92.180 124.240 92.240 ;
        RECT 113.850 92.010 114.140 92.060 ;
        RECT 110.090 91.870 114.140 92.010 ;
        RECT 113.850 91.830 114.140 91.870 ;
        RECT 117.680 92.010 118.000 92.070 ;
        RECT 118.650 92.010 118.940 92.060 ;
        RECT 117.680 91.870 118.940 92.010 ;
        RECT 117.680 91.810 118.000 91.870 ;
        RECT 118.650 91.830 118.940 91.870 ;
        RECT 29.850 91.640 30.140 91.690 ;
        RECT 26.960 91.500 30.140 91.640 ;
        RECT 26.960 91.440 27.280 91.500 ;
        RECT 29.850 91.460 30.140 91.500 ;
        RECT 30.330 91.460 30.620 91.690 ;
      LAYER met1 ;
        RECT 58.660 91.640 58.950 91.690 ;
        RECT 61.060 91.640 61.350 91.690 ;
        RECT 66.340 91.640 66.630 91.690 ;
        RECT 58.660 91.500 66.630 91.640 ;
        RECT 58.660 91.460 58.950 91.500 ;
        RECT 61.060 91.460 61.350 91.500 ;
        RECT 66.340 91.460 66.630 91.500 ;
      LAYER met1 ;
        RECT 72.080 91.640 72.400 91.700 ;
        RECT 78.810 91.640 79.100 91.690 ;
        RECT 79.760 91.640 80.080 91.700 ;
        RECT 85.520 91.640 85.840 91.700 ;
        RECT 92.240 91.640 92.560 91.700 ;
        RECT 72.080 91.500 80.080 91.640 ;
        RECT 85.320 91.500 85.840 91.640 ;
        RECT 92.040 91.500 92.560 91.640 ;
        RECT 72.080 91.440 72.400 91.500 ;
        RECT 78.810 91.460 79.100 91.500 ;
        RECT 79.760 91.440 80.080 91.500 ;
        RECT 85.520 91.440 85.840 91.500 ;
        RECT 92.240 91.440 92.560 91.500 ;
        RECT 92.720 91.640 93.040 91.700 ;
        RECT 98.970 91.640 99.260 91.690 ;
        RECT 105.690 91.640 105.980 91.690 ;
        RECT 92.720 91.500 105.980 91.640 ;
        RECT 92.720 91.440 93.040 91.500 ;
        RECT 98.970 91.460 99.260 91.500 ;
        RECT 105.690 91.460 105.980 91.500 ;
        RECT 108.080 91.640 108.400 91.700 ;
        RECT 110.970 91.640 111.260 91.690 ;
        RECT 114.810 91.640 115.100 91.690 ;
        RECT 108.080 91.500 115.100 91.640 ;
        RECT 29.360 91.270 29.680 91.330 ;
        RECT 35.120 91.270 35.440 91.330 ;
        RECT 26.570 91.130 35.440 91.270 ;
        RECT 29.360 91.070 29.680 91.130 ;
        RECT 35.120 91.070 35.440 91.130 ;
        RECT 59.610 91.270 59.900 91.320 ;
        RECT 63.920 91.270 64.240 91.330 ;
        RECT 59.610 91.130 64.240 91.270 ;
        RECT 105.770 91.270 105.910 91.460 ;
        RECT 108.080 91.440 108.400 91.500 ;
        RECT 110.970 91.460 111.260 91.500 ;
        RECT 114.810 91.460 115.100 91.500 ;
        RECT 124.880 91.640 125.200 91.700 ;
        RECT 125.370 91.640 125.660 91.690 ;
        RECT 124.880 91.500 125.660 91.640 ;
        RECT 124.880 91.440 125.200 91.500 ;
        RECT 125.370 91.460 125.660 91.500 ;
        RECT 110.480 91.270 110.800 91.330 ;
        RECT 105.770 91.130 110.800 91.270 ;
        RECT 59.610 91.090 59.900 91.130 ;
        RECT 63.920 91.070 64.240 91.130 ;
        RECT 110.480 91.070 110.800 91.130 ;
        RECT 28.400 90.900 28.720 90.960 ;
        RECT 33.210 90.900 33.500 90.950 ;
        RECT 28.400 90.760 33.500 90.900 ;
        RECT 28.400 90.700 28.720 90.760 ;
        RECT 33.210 90.720 33.500 90.760 ;
        RECT 117.210 90.900 117.500 90.950 ;
        RECT 120.560 90.900 120.880 90.960 ;
        RECT 117.210 90.760 120.880 90.900 ;
        RECT 117.210 90.720 117.500 90.760 ;
        RECT 120.560 90.700 120.880 90.760 ;
        RECT 14.480 90.530 14.800 90.590 ;
        RECT 34.640 90.530 34.960 90.590 ;
        RECT 14.280 90.390 14.800 90.530 ;
        RECT 34.440 90.390 34.960 90.530 ;
        RECT 14.480 90.330 14.800 90.390 ;
        RECT 34.640 90.330 34.960 90.390 ;
        RECT 71.120 90.530 71.440 90.590 ;
        RECT 71.610 90.530 71.900 90.580 ;
        RECT 71.120 90.390 71.900 90.530 ;
        RECT 71.120 90.330 71.440 90.390 ;
        RECT 71.610 90.350 71.900 90.390 ;
        RECT 26.960 88.680 27.280 88.740 ;
        RECT 27.450 88.680 27.740 88.730 ;
        RECT 53.360 88.680 53.680 88.740 ;
        RECT 57.680 88.680 58.000 88.740 ;
        RECT 63.920 88.680 64.240 88.740 ;
        RECT 26.960 88.540 27.740 88.680 ;
        RECT 53.160 88.540 53.680 88.680 ;
        RECT 57.480 88.540 58.000 88.680 ;
        RECT 63.720 88.540 64.240 88.680 ;
        RECT 26.960 88.480 27.280 88.540 ;
        RECT 27.450 88.500 27.740 88.540 ;
        RECT 53.360 88.480 53.680 88.540 ;
        RECT 57.680 88.480 58.000 88.540 ;
        RECT 63.920 88.480 64.240 88.540 ;
        RECT 64.400 88.680 64.720 88.740 ;
        RECT 65.370 88.680 65.660 88.730 ;
        RECT 64.400 88.540 65.660 88.680 ;
        RECT 64.400 88.480 64.720 88.540 ;
        RECT 65.370 88.500 65.660 88.540 ;
        RECT 69.690 88.680 69.980 88.730 ;
        RECT 86.480 88.680 86.800 88.740 ;
        RECT 69.690 88.540 86.800 88.680 ;
        RECT 69.690 88.500 69.980 88.540 ;
        RECT 86.480 88.480 86.800 88.540 ;
        RECT 107.120 88.680 107.440 88.740 ;
        RECT 110.970 88.680 111.260 88.730 ;
        RECT 118.160 88.680 118.480 88.740 ;
        RECT 107.120 88.540 111.260 88.680 ;
        RECT 117.960 88.540 118.480 88.680 ;
        RECT 107.120 88.480 107.440 88.540 ;
        RECT 110.970 88.500 111.260 88.540 ;
        RECT 118.160 88.480 118.480 88.540 ;
        RECT 21.690 88.310 21.980 88.360 ;
        RECT 29.360 88.310 29.680 88.370 ;
        RECT 21.690 88.170 29.680 88.310 ;
        RECT 21.690 88.130 21.980 88.170 ;
        RECT 29.360 88.110 29.680 88.170 ;
        RECT 28.890 87.940 29.180 87.990 ;
        RECT 33.680 87.940 34.000 88.000 ;
        RECT 98.960 87.940 99.280 88.000 ;
        RECT 28.890 87.800 42.550 87.940 ;
        RECT 28.890 87.760 29.180 87.800 ;
        RECT 29.360 87.570 29.680 87.630 ;
        RECT 21.290 87.430 29.680 87.570 ;
        RECT 21.290 87.250 21.430 87.430 ;
        RECT 29.360 87.370 29.680 87.430 ;
        RECT 21.210 87.020 21.500 87.250 ;
        RECT 24.570 87.200 24.860 87.250 ;
        RECT 29.930 87.200 30.070 87.800 ;
        RECT 33.680 87.740 34.000 87.800 ;
        RECT 42.410 87.620 42.550 87.800 ;
        RECT 74.090 87.800 99.280 87.940 ;
        RECT 35.610 87.570 35.900 87.620 ;
        RECT 35.610 87.430 38.710 87.570 ;
        RECT 35.610 87.390 35.900 87.430 ;
        RECT 31.760 87.200 32.080 87.260 ;
        RECT 38.570 87.250 38.710 87.430 ;
        RECT 42.330 87.390 42.620 87.620 ;
        RECT 49.040 87.570 49.360 87.630 ;
        RECT 48.840 87.430 49.360 87.570 ;
        RECT 49.040 87.370 49.360 87.430 ;
        RECT 53.840 87.570 54.160 87.630 ;
        RECT 54.330 87.570 54.620 87.620 ;
        RECT 55.280 87.570 55.600 87.630 ;
        RECT 59.120 87.570 59.440 87.630 ;
        RECT 53.840 87.430 54.620 87.570 ;
        RECT 55.080 87.430 55.600 87.570 ;
        RECT 58.920 87.430 59.440 87.570 ;
        RECT 53.840 87.370 54.160 87.430 ;
        RECT 54.330 87.390 54.620 87.430 ;
        RECT 55.280 87.370 55.600 87.430 ;
        RECT 59.120 87.370 59.440 87.430 ;
        RECT 24.570 87.060 30.070 87.200 ;
        RECT 31.560 87.060 32.080 87.200 ;
        RECT 24.570 87.020 24.860 87.060 ;
        RECT 31.760 87.000 32.080 87.060 ;
        RECT 38.490 87.020 38.780 87.250 ;
        RECT 51.930 87.200 52.220 87.250 ;
        RECT 52.880 87.200 53.200 87.260 ;
        RECT 60.080 87.200 60.400 87.260 ;
        RECT 39.050 87.060 52.220 87.200 ;
        RECT 52.680 87.060 53.200 87.200 ;
        RECT 59.880 87.060 60.400 87.200 ;
        RECT 25.050 86.830 25.340 86.880 ;
        RECT 34.640 86.830 34.960 86.890 ;
        RECT 25.050 86.690 34.960 86.830 ;
        RECT 25.050 86.650 25.340 86.690 ;
        RECT 34.640 86.630 34.960 86.690 ;
        RECT 35.120 86.830 35.440 86.890 ;
        RECT 39.050 86.830 39.190 87.060 ;
        RECT 51.930 87.020 52.220 87.060 ;
        RECT 52.880 87.000 53.200 87.060 ;
        RECT 60.080 87.000 60.400 87.060 ;
        RECT 61.530 87.020 61.820 87.250 ;
        RECT 69.210 87.200 69.500 87.250 ;
        RECT 72.570 87.200 72.860 87.250 ;
        RECT 74.090 87.200 74.230 87.800 ;
        RECT 98.960 87.740 99.280 87.800 ;
        RECT 101.850 87.940 102.140 87.990 ;
        RECT 114.810 87.940 115.100 87.990 ;
        RECT 101.850 87.800 115.100 87.940 ;
        RECT 101.850 87.760 102.140 87.800 ;
        RECT 114.810 87.760 115.100 87.800 ;
        RECT 81.210 87.570 81.500 87.620 ;
        RECT 86.480 87.570 86.800 87.630 ;
        RECT 87.920 87.570 88.240 87.630 ;
        RECT 97.520 87.570 97.840 87.630 ;
        RECT 103.280 87.570 103.600 87.630 ;
        RECT 109.050 87.570 109.340 87.620 ;
        RECT 110.480 87.570 110.800 87.630 ;
        RECT 81.210 87.430 86.800 87.570 ;
        RECT 87.720 87.430 88.240 87.570 ;
        RECT 97.320 87.430 97.840 87.570 ;
        RECT 103.080 87.430 103.600 87.570 ;
        RECT 81.210 87.390 81.500 87.430 ;
        RECT 86.480 87.370 86.800 87.430 ;
        RECT 87.920 87.370 88.240 87.430 ;
        RECT 97.520 87.370 97.840 87.430 ;
        RECT 103.280 87.370 103.600 87.430 ;
        RECT 103.850 87.430 109.340 87.570 ;
        RECT 110.280 87.430 110.800 87.570 ;
        RECT 84.090 87.200 84.380 87.250 ;
        RECT 69.210 87.060 74.230 87.200 ;
        RECT 74.570 87.060 84.380 87.200 ;
        RECT 69.210 87.020 69.500 87.060 ;
        RECT 72.570 87.020 72.860 87.060 ;
        RECT 35.120 86.690 39.190 86.830 ;
        RECT 35.120 86.630 35.440 86.690 ;
        RECT 46.650 86.650 46.940 86.880 ;
        RECT 61.610 86.830 61.750 87.020 ;
        RECT 71.120 86.830 71.440 86.890 ;
        RECT 74.570 86.880 74.710 87.060 ;
        RECT 84.090 87.020 84.380 87.060 ;
        RECT 92.240 87.200 92.560 87.260 ;
        RECT 93.690 87.200 93.980 87.250 ;
        RECT 92.240 87.060 93.980 87.200 ;
        RECT 92.240 87.000 92.560 87.060 ;
        RECT 93.690 87.020 93.980 87.060 ;
        RECT 100.400 87.200 100.720 87.260 ;
        RECT 103.850 87.200 103.990 87.430 ;
        RECT 109.050 87.390 109.340 87.430 ;
        RECT 110.480 87.370 110.800 87.430 ;
        RECT 100.400 87.060 103.990 87.200 ;
        RECT 119.610 87.200 119.900 87.250 ;
        RECT 120.560 87.200 120.880 87.260 ;
        RECT 119.610 87.060 120.880 87.200 ;
        RECT 100.400 87.000 100.720 87.060 ;
        RECT 119.610 87.020 119.900 87.060 ;
        RECT 120.560 87.000 120.880 87.060 ;
        RECT 74.010 86.830 74.300 86.880 ;
        RECT 61.610 86.690 74.300 86.830 ;
        RECT 26.000 86.460 26.320 86.520 ;
        RECT 46.730 86.460 46.870 86.650 ;
        RECT 71.120 86.630 71.440 86.690 ;
        RECT 74.010 86.650 74.300 86.690 ;
        RECT 74.490 86.650 74.780 86.880 ;
        RECT 79.770 86.830 80.060 86.880 ;
        RECT 80.240 86.830 80.560 86.890 ;
        RECT 79.770 86.690 80.560 86.830 ;
        RECT 79.770 86.650 80.060 86.690 ;
        RECT 80.240 86.630 80.560 86.690 ;
        RECT 104.730 86.650 105.020 86.880 ;
        RECT 74.960 86.460 75.280 86.520 ;
        RECT 26.000 86.320 46.870 86.460 ;
        RECT 74.760 86.320 75.280 86.460 ;
        RECT 26.000 86.260 26.320 86.320 ;
        RECT 74.960 86.260 75.280 86.320 ;
        RECT 104.240 86.460 104.560 86.520 ;
        RECT 104.810 86.460 104.950 86.650 ;
        RECT 113.360 86.460 113.680 86.520 ;
        RECT 104.240 86.320 104.950 86.460 ;
        RECT 113.160 86.320 113.680 86.460 ;
        RECT 104.240 86.260 104.560 86.320 ;
        RECT 113.360 86.260 113.680 86.320 ;
        RECT 5.760 85.730 142.080 86.100 ;
        RECT 11.130 84.610 11.420 84.660 ;
        RECT 21.680 84.610 22.000 84.670 ;
        RECT 11.130 84.470 22.000 84.610 ;
        RECT 11.130 84.430 11.420 84.470 ;
        RECT 21.680 84.410 22.000 84.470 ;
        RECT 22.650 84.610 22.940 84.660 ;
        RECT 24.080 84.610 24.400 84.670 ;
        RECT 49.520 84.610 49.840 84.670 ;
        RECT 102.330 84.610 102.620 84.660 ;
        RECT 107.600 84.610 107.920 84.670 ;
        RECT 22.650 84.470 24.400 84.610 ;
        RECT 22.650 84.430 22.940 84.470 ;
        RECT 24.080 84.410 24.400 84.470 ;
        RECT 26.570 84.470 49.840 84.610 ;
        RECT 19.280 84.240 19.600 84.300 ;
        RECT 19.080 84.100 19.600 84.240 ;
        RECT 19.280 84.040 19.600 84.100 ;
        RECT 19.760 84.240 20.080 84.300 ;
        RECT 26.570 84.240 26.710 84.470 ;
        RECT 49.520 84.410 49.840 84.470 ;
        RECT 74.090 84.470 82.870 84.610 ;
        RECT 32.240 84.240 32.560 84.300 ;
        RECT 19.760 84.100 26.710 84.240 ;
        RECT 19.760 84.040 20.080 84.100 ;
        RECT 26.570 83.920 26.710 84.100 ;
        RECT 29.930 84.100 32.560 84.240 ;
        RECT 29.930 83.930 30.070 84.100 ;
        RECT 32.240 84.040 32.560 84.100 ;
        RECT 72.080 84.240 72.400 84.300 ;
        RECT 73.530 84.240 73.820 84.290 ;
        RECT 72.080 84.100 73.820 84.240 ;
        RECT 72.080 84.040 72.400 84.100 ;
        RECT 73.530 84.060 73.820 84.100 ;
        RECT 26.490 83.690 26.780 83.920 ;
        RECT 29.370 83.870 29.660 83.920 ;
        RECT 29.840 83.870 30.160 83.930 ;
        RECT 29.370 83.730 30.160 83.870 ;
        RECT 29.370 83.690 29.660 83.730 ;
        RECT 29.840 83.670 30.160 83.730 ;
        RECT 30.330 83.870 30.620 83.920 ;
        RECT 34.640 83.870 34.960 83.930 ;
        RECT 30.330 83.730 34.960 83.870 ;
        RECT 30.330 83.690 30.620 83.730 ;
        RECT 34.640 83.670 34.960 83.730 ;
        RECT 36.560 83.870 36.880 83.930 ;
        RECT 39.450 83.870 39.740 83.920 ;
        RECT 36.560 83.730 39.740 83.870 ;
        RECT 36.560 83.670 36.880 83.730 ;
        RECT 39.450 83.690 39.740 83.730 ;
        RECT 45.200 83.870 45.520 83.930 ;
        RECT 74.090 83.920 74.230 84.470 ;
        RECT 74.960 84.240 75.280 84.300 ;
        RECT 77.370 84.240 77.660 84.290 ;
        RECT 78.330 84.240 78.620 84.290 ;
        RECT 79.280 84.240 79.600 84.300 ;
        RECT 74.960 84.100 78.070 84.240 ;
        RECT 74.960 84.040 75.280 84.100 ;
        RECT 77.370 84.060 77.660 84.100 ;
        RECT 49.050 83.870 49.340 83.920 ;
        RECT 45.200 83.730 49.340 83.870 ;
        RECT 45.200 83.670 45.520 83.730 ;
        RECT 49.050 83.690 49.340 83.730 ;
        RECT 55.770 83.690 56.060 83.920 ;
        RECT 72.570 83.690 72.860 83.920 ;
        RECT 74.010 83.690 74.300 83.920 ;
      LAYER met1 ;
        RECT 9.700 83.500 9.990 83.550 ;
        RECT 12.100 83.500 12.390 83.550 ;
        RECT 17.380 83.500 17.670 83.550 ;
      LAYER met1 ;
        RECT 31.760 83.500 32.080 83.560 ;
      LAYER met1 ;
        RECT 9.700 83.360 17.670 83.500 ;
      LAYER met1 ;
        RECT 31.560 83.360 32.080 83.500 ;
      LAYER met1 ;
        RECT 9.700 83.320 9.990 83.360 ;
        RECT 12.100 83.320 12.390 83.360 ;
        RECT 17.380 83.320 17.670 83.360 ;
      LAYER met1 ;
        RECT 31.760 83.300 32.080 83.360 ;
        RECT 32.730 83.500 33.020 83.550 ;
        RECT 35.120 83.500 35.440 83.560 ;
        RECT 32.730 83.360 35.440 83.500 ;
        RECT 32.730 83.320 33.020 83.360 ;
        RECT 35.120 83.300 35.440 83.360 ;
        RECT 43.290 83.500 43.580 83.550 ;
        RECT 44.240 83.500 44.560 83.560 ;
        RECT 43.290 83.360 44.560 83.500 ;
        RECT 43.290 83.320 43.580 83.360 ;
        RECT 44.240 83.300 44.560 83.360 ;
        RECT 52.890 83.500 53.180 83.550 ;
        RECT 55.850 83.500 55.990 83.690 ;
        RECT 59.600 83.500 59.920 83.560 ;
        RECT 52.890 83.360 55.990 83.500 ;
        RECT 59.400 83.360 59.920 83.500 ;
        RECT 72.650 83.500 72.790 83.690 ;
        RECT 76.890 83.500 77.180 83.550 ;
        RECT 72.650 83.360 77.180 83.500 ;
        RECT 77.930 83.500 78.070 84.100 ;
        RECT 78.330 84.100 79.600 84.240 ;
        RECT 78.330 84.060 78.620 84.100 ;
        RECT 79.280 84.040 79.600 84.100 ;
        RECT 82.730 84.240 82.870 84.470 ;
        RECT 102.330 84.470 107.920 84.610 ;
        RECT 102.330 84.430 102.620 84.470 ;
        RECT 107.600 84.410 107.920 84.470 ;
        RECT 108.570 84.610 108.860 84.660 ;
        RECT 113.360 84.610 113.680 84.670 ;
        RECT 108.570 84.470 113.680 84.610 ;
        RECT 108.570 84.430 108.860 84.470 ;
        RECT 113.360 84.410 113.680 84.470 ;
        RECT 86.480 84.240 86.800 84.300 ;
        RECT 111.920 84.240 112.240 84.300 ;
        RECT 114.800 84.240 115.120 84.300 ;
        RECT 116.730 84.240 117.020 84.290 ;
        RECT 82.730 84.100 84.790 84.240 ;
        RECT 82.730 83.920 82.870 84.100 ;
        RECT 84.650 83.930 84.790 84.100 ;
        RECT 86.480 84.100 94.870 84.240 ;
        RECT 86.480 84.040 86.800 84.100 ;
        RECT 82.650 83.690 82.940 83.920 ;
        RECT 84.560 83.870 84.880 83.930 ;
        RECT 94.730 83.920 94.870 84.100 ;
        RECT 111.920 84.100 117.020 84.240 ;
        RECT 111.920 84.040 112.240 84.100 ;
        RECT 114.800 84.040 115.120 84.100 ;
        RECT 116.730 84.060 117.020 84.100 ;
        RECT 84.360 83.730 84.880 83.870 ;
        RECT 84.560 83.670 84.880 83.730 ;
        RECT 85.530 83.870 85.820 83.920 ;
        RECT 87.930 83.870 88.220 83.920 ;
        RECT 85.530 83.730 88.220 83.870 ;
        RECT 85.530 83.690 85.820 83.730 ;
        RECT 87.930 83.690 88.220 83.730 ;
        RECT 94.650 83.690 94.940 83.920 ;
        RECT 101.360 83.870 101.680 83.930 ;
        RECT 101.160 83.730 101.680 83.870 ;
        RECT 101.360 83.670 101.680 83.730 ;
        RECT 91.760 83.500 92.080 83.560 ;
        RECT 77.930 83.360 82.870 83.500 ;
        RECT 91.560 83.360 92.080 83.500 ;
        RECT 52.890 83.320 53.180 83.360 ;
        RECT 59.600 83.300 59.920 83.360 ;
        RECT 76.890 83.320 77.180 83.360 ;
        RECT 25.050 82.760 25.340 82.810 ;
        RECT 31.280 82.760 31.600 82.820 ;
        RECT 25.050 82.620 31.600 82.760 ;
        RECT 25.050 82.580 25.340 82.620 ;
        RECT 31.280 82.560 31.600 82.620 ;
        RECT 50.480 82.760 50.800 82.820 ;
        RECT 66.330 82.760 66.620 82.810 ;
        RECT 50.480 82.620 66.620 82.760 ;
        RECT 76.970 82.760 77.110 83.320 ;
        RECT 82.730 83.130 82.870 83.360 ;
        RECT 91.760 83.300 92.080 83.360 ;
        RECT 98.490 83.320 98.780 83.550 ;
      LAYER met1 ;
        RECT 107.140 83.500 107.430 83.550 ;
        RECT 109.540 83.500 109.830 83.550 ;
        RECT 114.820 83.500 115.110 83.550 ;
        RECT 107.140 83.360 115.110 83.500 ;
        RECT 107.140 83.320 107.430 83.360 ;
        RECT 109.540 83.320 109.830 83.360 ;
        RECT 114.820 83.320 115.110 83.360 ;
      LAYER met1 ;
        RECT 85.040 83.130 85.360 83.190 ;
        RECT 98.570 83.130 98.710 83.320 ;
        RECT 82.730 82.990 98.710 83.130 ;
        RECT 85.040 82.930 85.360 82.990 ;
        RECT 91.760 82.760 92.080 82.820 ;
        RECT 76.970 82.620 92.080 82.760 ;
        RECT 50.480 82.560 50.800 82.620 ;
        RECT 66.330 82.580 66.620 82.620 ;
        RECT 91.760 82.560 92.080 82.620 ;
        RECT 30.800 82.390 31.120 82.450 ;
        RECT 35.120 82.390 35.440 82.450 ;
        RECT 30.600 82.250 31.120 82.390 ;
        RECT 34.920 82.250 35.440 82.390 ;
        RECT 30.800 82.190 31.120 82.250 ;
        RECT 35.120 82.190 35.440 82.250 ;
        RECT 36.080 82.390 36.400 82.450 ;
        RECT 36.570 82.390 36.860 82.440 ;
        RECT 36.080 82.250 36.860 82.390 ;
        RECT 36.080 82.190 36.400 82.250 ;
        RECT 36.570 82.210 36.860 82.250 ;
        RECT 64.880 82.390 65.200 82.450 ;
        RECT 79.760 82.390 80.080 82.450 ;
        RECT 64.880 82.250 65.400 82.390 ;
        RECT 79.560 82.250 80.080 82.390 ;
        RECT 64.880 82.190 65.200 82.250 ;
        RECT 79.760 82.190 80.080 82.250 ;
        RECT 83.130 82.390 83.420 82.440 ;
        RECT 90.800 82.390 91.120 82.450 ;
        RECT 83.130 82.250 91.120 82.390 ;
        RECT 83.130 82.210 83.420 82.250 ;
        RECT 90.800 82.190 91.120 82.250 ;
        RECT 14.970 80.540 15.260 80.590 ;
        RECT 19.280 80.540 19.600 80.600 ;
        RECT 14.970 80.400 19.600 80.540 ;
        RECT 14.970 80.360 15.260 80.400 ;
        RECT 19.280 80.340 19.600 80.400 ;
        RECT 29.360 80.540 29.680 80.600 ;
        RECT 38.010 80.540 38.300 80.590 ;
        RECT 29.360 80.400 38.300 80.540 ;
        RECT 29.360 80.340 29.680 80.400 ;
        RECT 38.010 80.360 38.300 80.400 ;
        RECT 57.210 80.540 57.500 80.590 ;
        RECT 60.080 80.540 60.400 80.600 ;
        RECT 57.210 80.400 60.400 80.540 ;
        RECT 57.210 80.360 57.500 80.400 ;
        RECT 60.080 80.340 60.400 80.400 ;
        RECT 74.490 80.540 74.780 80.590 ;
        RECT 79.760 80.540 80.080 80.600 ;
        RECT 74.490 80.400 80.080 80.540 ;
        RECT 74.490 80.360 74.780 80.400 ;
        RECT 79.760 80.340 80.080 80.400 ;
        RECT 102.810 80.540 103.100 80.590 ;
        RECT 103.280 80.540 103.600 80.600 ;
        RECT 102.810 80.400 103.600 80.540 ;
        RECT 102.810 80.360 103.100 80.400 ;
        RECT 103.280 80.340 103.600 80.400 ;
        RECT 114.800 80.540 115.120 80.600 ;
        RECT 116.240 80.540 116.560 80.600 ;
        RECT 114.800 80.400 116.560 80.540 ;
        RECT 114.800 80.340 115.120 80.400 ;
        RECT 116.240 80.340 116.560 80.400 ;
        RECT 72.080 80.170 72.400 80.230 ;
        RECT 95.120 80.170 95.440 80.230 ;
        RECT 72.080 80.030 95.440 80.170 ;
        RECT 72.080 79.970 72.400 80.030 ;
        RECT 95.120 79.970 95.440 80.030 ;
        RECT 101.360 80.170 101.680 80.230 ;
        RECT 124.890 80.170 125.180 80.220 ;
        RECT 101.360 80.030 125.180 80.170 ;
        RECT 101.360 79.970 101.680 80.030 ;
        RECT 124.890 79.990 125.180 80.030 ;
        RECT 35.120 79.800 35.440 79.860 ;
        RECT 104.240 79.800 104.560 79.860 ;
        RECT 130.640 79.800 130.960 79.860 ;
        RECT 22.730 79.660 35.440 79.800 ;
        RECT 22.730 79.120 22.870 79.660 ;
        RECT 35.120 79.600 35.440 79.660 ;
        RECT 83.690 79.660 104.560 79.800 ;
      LAYER met1 ;
        RECT 25.060 79.440 25.350 79.480 ;
        RECT 27.460 79.440 27.750 79.480 ;
        RECT 32.740 79.440 33.030 79.480 ;
        RECT 25.060 79.300 33.030 79.440 ;
        RECT 25.060 79.250 25.350 79.300 ;
        RECT 27.460 79.250 27.750 79.300 ;
        RECT 32.740 79.250 33.030 79.300 ;
        RECT 44.260 79.440 44.550 79.480 ;
        RECT 46.660 79.440 46.950 79.480 ;
        RECT 51.940 79.440 52.230 79.480 ;
        RECT 44.260 79.300 52.230 79.440 ;
        RECT 44.260 79.250 44.550 79.300 ;
        RECT 46.660 79.250 46.950 79.300 ;
        RECT 51.940 79.250 52.230 79.300 ;
      LAYER met1 ;
        RECT 65.370 79.430 65.660 79.480 ;
        RECT 70.640 79.430 70.960 79.490 ;
        RECT 83.690 79.430 83.830 79.660 ;
        RECT 104.240 79.600 104.560 79.660 ;
        RECT 115.370 79.660 130.960 79.800 ;
        RECT 85.040 79.430 85.360 79.490 ;
        RECT 91.760 79.430 92.080 79.490 ;
        RECT 65.370 79.290 70.960 79.430 ;
        RECT 65.370 79.250 65.660 79.290 ;
        RECT 70.640 79.230 70.960 79.290 ;
        RECT 78.890 79.290 83.830 79.430 ;
        RECT 84.840 79.290 85.360 79.430 ;
        RECT 91.560 79.290 92.080 79.430 ;
        RECT 14.480 79.060 14.800 79.120 ;
        RECT 16.410 79.060 16.700 79.110 ;
        RECT 22.640 79.060 22.960 79.120 ;
        RECT 14.480 78.920 22.960 79.060 ;
        RECT 14.480 78.860 14.800 78.920 ;
        RECT 16.410 78.880 16.700 78.920 ;
        RECT 22.640 78.860 22.960 78.920 ;
        RECT 26.490 79.060 26.780 79.110 ;
        RECT 30.800 79.060 31.120 79.120 ;
        RECT 26.490 78.920 31.120 79.060 ;
        RECT 26.490 78.880 26.780 78.920 ;
        RECT 30.800 78.860 31.120 78.920 ;
        RECT 31.280 79.060 31.600 79.120 ;
        RECT 45.210 79.060 45.500 79.110 ;
        RECT 31.280 78.920 45.500 79.060 ;
        RECT 31.280 78.860 31.600 78.920 ;
        RECT 45.210 78.880 45.500 78.920 ;
        RECT 62.490 79.060 62.780 79.110 ;
        RECT 70.160 79.060 70.480 79.120 ;
        RECT 71.600 79.060 71.920 79.120 ;
        RECT 62.490 78.920 70.480 79.060 ;
        RECT 71.400 78.920 71.920 79.060 ;
        RECT 62.490 78.880 62.780 78.920 ;
        RECT 70.160 78.860 70.480 78.920 ;
        RECT 71.600 78.860 71.920 78.920 ;
        RECT 72.560 78.690 72.880 78.750 ;
        RECT 74.970 78.690 75.260 78.740 ;
        RECT 78.890 78.690 79.030 79.290 ;
        RECT 85.040 79.230 85.360 79.290 ;
        RECT 91.760 79.230 92.080 79.290 ;
        RECT 95.120 79.430 95.440 79.490 ;
        RECT 100.400 79.430 100.720 79.490 ;
        RECT 111.930 79.430 112.220 79.480 ;
        RECT 115.370 79.430 115.510 79.660 ;
        RECT 130.640 79.600 130.960 79.660 ;
        RECT 116.240 79.430 116.560 79.490 ;
        RECT 120.570 79.430 120.860 79.480 ;
        RECT 95.120 79.290 106.390 79.430 ;
        RECT 95.120 79.230 95.440 79.290 ;
        RECT 100.400 79.230 100.720 79.290 ;
        RECT 83.690 78.920 105.910 79.060 ;
        RECT 83.690 78.740 83.830 78.920 ;
        RECT 72.560 78.550 79.030 78.690 ;
        RECT 72.560 78.490 72.880 78.550 ;
        RECT 74.970 78.510 75.260 78.550 ;
        RECT 83.610 78.510 83.900 78.740 ;
        RECT 84.080 78.690 84.400 78.750 ;
        RECT 89.370 78.690 89.660 78.740 ;
        RECT 84.080 78.550 89.660 78.690 ;
        RECT 84.080 78.490 84.400 78.550 ;
        RECT 89.370 78.510 89.660 78.550 ;
        RECT 91.760 78.690 92.080 78.750 ;
        RECT 100.490 78.740 100.630 78.920 ;
        RECT 95.130 78.690 95.420 78.740 ;
        RECT 91.760 78.550 95.420 78.690 ;
        RECT 91.760 78.490 92.080 78.550 ;
        RECT 95.130 78.510 95.420 78.550 ;
        RECT 96.090 78.510 96.380 78.740 ;
        RECT 100.410 78.510 100.700 78.740 ;
        RECT 101.370 78.690 101.660 78.740 ;
        RECT 102.320 78.690 102.640 78.750 ;
        RECT 105.770 78.740 105.910 78.920 ;
        RECT 101.370 78.550 102.640 78.690 ;
        RECT 101.370 78.510 101.660 78.550 ;
        RECT 21.680 78.320 22.000 78.380 ;
        RECT 26.010 78.320 26.300 78.370 ;
        RECT 45.680 78.320 46.000 78.380 ;
        RECT 21.680 78.180 26.300 78.320 ;
        RECT 45.480 78.180 46.000 78.320 ;
        RECT 21.680 78.120 22.000 78.180 ;
        RECT 26.010 78.140 26.300 78.180 ;
        RECT 45.680 78.120 46.000 78.180 ;
        RECT 84.560 78.320 84.880 78.380 ;
        RECT 96.170 78.320 96.310 78.510 ;
        RECT 84.560 78.180 96.310 78.320 ;
        RECT 97.530 78.320 97.820 78.370 ;
        RECT 101.450 78.320 101.590 78.510 ;
        RECT 102.320 78.490 102.640 78.550 ;
        RECT 105.690 78.510 105.980 78.740 ;
        RECT 106.250 78.690 106.390 79.290 ;
        RECT 111.930 79.290 115.510 79.430 ;
        RECT 115.800 79.290 120.860 79.430 ;
        RECT 111.930 79.250 112.220 79.290 ;
        RECT 116.240 79.230 116.560 79.290 ;
        RECT 120.570 79.250 120.860 79.290 ;
        RECT 106.650 78.690 106.940 78.740 ;
        RECT 106.250 78.550 106.940 78.690 ;
        RECT 106.650 78.510 106.940 78.550 ;
        RECT 107.120 78.690 107.440 78.750 ;
        RECT 110.490 78.690 110.780 78.740 ;
        RECT 107.120 78.550 110.780 78.690 ;
        RECT 107.120 78.490 107.440 78.550 ;
        RECT 110.490 78.510 110.780 78.550 ;
        RECT 108.080 78.320 108.400 78.380 ;
        RECT 114.800 78.320 115.120 78.380 ;
        RECT 119.120 78.320 119.440 78.380 ;
        RECT 123.440 78.320 123.760 78.380 ;
        RECT 97.530 78.180 101.590 78.320 ;
        RECT 107.880 78.180 108.400 78.320 ;
        RECT 114.600 78.180 115.120 78.320 ;
        RECT 118.920 78.180 119.440 78.320 ;
        RECT 123.240 78.180 123.760 78.320 ;
        RECT 84.560 78.120 84.880 78.180 ;
        RECT 97.530 78.140 97.820 78.180 ;
        RECT 108.080 78.120 108.400 78.180 ;
        RECT 114.800 78.120 115.120 78.180 ;
        RECT 119.120 78.120 119.440 78.180 ;
        RECT 123.440 78.120 123.760 78.180 ;
        RECT 5.760 77.590 142.080 77.960 ;
        RECT 21.680 76.470 22.000 76.530 ;
        RECT 45.680 76.470 46.000 76.530 ;
        RECT 21.480 76.330 22.000 76.470 ;
        RECT 21.680 76.270 22.000 76.330 ;
        RECT 28.010 76.330 46.000 76.470 ;
        RECT 17.370 76.100 17.660 76.150 ;
        RECT 28.010 76.100 28.150 76.330 ;
        RECT 45.680 76.270 46.000 76.330 ;
        RECT 64.890 76.470 65.180 76.520 ;
        RECT 65.360 76.470 65.680 76.530 ;
        RECT 114.800 76.470 115.120 76.530 ;
        RECT 64.890 76.330 65.680 76.470 ;
        RECT 64.890 76.290 65.180 76.330 ;
        RECT 65.360 76.270 65.680 76.330 ;
        RECT 73.130 76.330 115.120 76.470 ;
        RECT 17.370 75.960 28.150 76.100 ;
        RECT 28.410 76.100 28.700 76.150 ;
        RECT 31.760 76.100 32.080 76.160 ;
        RECT 28.410 75.960 32.080 76.100 ;
        RECT 17.370 75.920 17.660 75.960 ;
        RECT 28.410 75.920 28.700 75.960 ;
        RECT 31.760 75.900 32.080 75.960 ;
        RECT 35.130 75.920 35.420 76.150 ;
        RECT 41.850 76.100 42.140 76.150 ;
        RECT 43.760 76.100 44.080 76.160 ;
        RECT 41.850 75.960 44.080 76.100 ;
        RECT 41.850 75.920 42.140 75.960 ;
        RECT 35.210 75.730 35.350 75.920 ;
        RECT 43.760 75.900 44.080 75.960 ;
        RECT 57.690 76.100 57.980 76.150 ;
        RECT 71.120 76.100 71.440 76.160 ;
        RECT 72.560 76.100 72.880 76.160 ;
        RECT 73.130 76.150 73.270 76.330 ;
        RECT 114.800 76.270 115.120 76.330 ;
        RECT 116.730 76.470 117.020 76.520 ;
        RECT 119.120 76.470 119.440 76.530 ;
        RECT 116.730 76.330 119.440 76.470 ;
        RECT 116.730 76.290 117.020 76.330 ;
        RECT 119.120 76.270 119.440 76.330 ;
        RECT 57.690 75.960 72.880 76.100 ;
        RECT 57.690 75.920 57.980 75.960 ;
        RECT 71.120 75.900 71.440 75.960 ;
        RECT 72.560 75.900 72.880 75.960 ;
        RECT 73.050 75.920 73.340 76.150 ;
        RECT 82.640 76.100 82.960 76.160 ;
        RECT 98.490 76.100 98.780 76.150 ;
        RECT 101.360 76.100 101.680 76.160 ;
        RECT 104.240 76.100 104.560 76.160 ;
        RECT 82.440 75.960 82.960 76.100 ;
        RECT 82.640 75.900 82.960 75.960 ;
        RECT 86.570 75.960 98.780 76.100 ;
        RECT 101.160 75.960 101.680 76.100 ;
        RECT 104.040 75.960 104.560 76.100 ;
        RECT 44.720 75.730 45.040 75.790 ;
        RECT 47.600 75.730 47.920 75.790 ;
        RECT 35.210 75.590 45.040 75.730 ;
        RECT 47.400 75.590 47.920 75.730 ;
        RECT 44.720 75.530 45.040 75.590 ;
        RECT 47.600 75.530 47.920 75.590 ;
        RECT 57.690 75.730 57.980 75.780 ;
        RECT 60.080 75.730 60.400 75.790 ;
        RECT 79.280 75.730 79.600 75.790 ;
        RECT 57.690 75.590 60.400 75.730 ;
        RECT 79.080 75.590 79.600 75.730 ;
        RECT 57.690 75.550 57.980 75.590 ;
        RECT 60.080 75.530 60.400 75.590 ;
        RECT 79.280 75.530 79.600 75.590 ;
        RECT 80.250 75.730 80.540 75.780 ;
        RECT 84.560 75.730 84.880 75.790 ;
        RECT 86.570 75.780 86.710 75.960 ;
        RECT 98.490 75.920 98.780 75.960 ;
        RECT 101.360 75.900 101.680 75.960 ;
        RECT 104.240 75.900 104.560 75.960 ;
        RECT 110.970 76.100 111.260 76.150 ;
        RECT 117.210 76.100 117.500 76.150 ;
        RECT 123.440 76.100 123.760 76.160 ;
        RECT 110.970 75.960 116.950 76.100 ;
        RECT 110.970 75.920 111.260 75.960 ;
        RECT 116.810 75.790 116.950 75.960 ;
        RECT 117.210 75.960 123.760 76.100 ;
        RECT 117.210 75.920 117.500 75.960 ;
        RECT 123.440 75.900 123.760 75.960 ;
        RECT 80.250 75.590 84.880 75.730 ;
        RECT 80.250 75.550 80.540 75.590 ;
        RECT 84.560 75.530 84.880 75.590 ;
        RECT 86.490 75.550 86.780 75.780 ;
        RECT 86.970 75.730 87.260 75.780 ;
        RECT 89.850 75.730 90.140 75.780 ;
        RECT 93.680 75.730 94.000 75.790 ;
        RECT 86.970 75.590 90.140 75.730 ;
        RECT 93.480 75.590 94.000 75.730 ;
        RECT 86.970 75.550 87.260 75.590 ;
        RECT 89.850 75.550 90.140 75.590 ;
        RECT 93.680 75.530 94.000 75.590 ;
        RECT 96.560 75.730 96.880 75.790 ;
        RECT 97.050 75.730 97.340 75.780 ;
        RECT 96.560 75.590 97.340 75.730 ;
        RECT 96.560 75.530 96.880 75.590 ;
        RECT 97.050 75.550 97.340 75.590 ;
        RECT 105.690 75.730 105.980 75.780 ;
        RECT 108.080 75.730 108.400 75.790 ;
        RECT 110.000 75.730 110.320 75.790 ;
        RECT 105.690 75.590 108.400 75.730 ;
        RECT 109.800 75.590 110.320 75.730 ;
        RECT 105.690 75.550 105.980 75.590 ;
        RECT 108.080 75.530 108.400 75.590 ;
        RECT 110.000 75.530 110.320 75.590 ;
        RECT 111.450 75.730 111.740 75.780 ;
        RECT 113.370 75.730 113.660 75.780 ;
        RECT 111.450 75.590 113.660 75.730 ;
        RECT 111.450 75.550 111.740 75.590 ;
        RECT 113.370 75.550 113.660 75.590 ;
        RECT 116.720 75.530 117.040 75.790 ;
        RECT 29.360 75.360 29.680 75.420 ;
        RECT 29.850 75.360 30.140 75.410 ;
        RECT 36.560 75.360 36.880 75.420 ;
        RECT 43.280 75.360 43.600 75.420 ;
        RECT 29.360 75.220 30.140 75.360 ;
        RECT 36.360 75.220 36.880 75.360 ;
        RECT 43.080 75.220 43.600 75.360 ;
        RECT 29.360 75.160 29.680 75.220 ;
        RECT 29.850 75.180 30.140 75.220 ;
        RECT 36.560 75.160 36.880 75.220 ;
        RECT 43.280 75.160 43.600 75.220 ;
        RECT 51.450 75.360 51.740 75.410 ;
        RECT 58.160 75.360 58.480 75.420 ;
        RECT 51.450 75.220 58.480 75.360 ;
        RECT 51.450 75.180 51.740 75.220 ;
        RECT 58.160 75.160 58.480 75.220 ;
      LAYER met1 ;
        RECT 63.460 75.360 63.750 75.410 ;
        RECT 65.860 75.360 66.150 75.410 ;
        RECT 71.140 75.360 71.430 75.410 ;
      LAYER met1 ;
        RECT 85.040 75.360 85.360 75.420 ;
      LAYER met1 ;
        RECT 63.460 75.220 71.430 75.360 ;
      LAYER met1 ;
        RECT 84.840 75.220 85.360 75.360 ;
      LAYER met1 ;
        RECT 63.460 75.180 63.750 75.220 ;
        RECT 65.860 75.180 66.150 75.220 ;
        RECT 71.140 75.180 71.430 75.220 ;
      LAYER met1 ;
        RECT 85.040 75.160 85.360 75.220 ;
        RECT 85.520 75.360 85.840 75.420 ;
        RECT 90.800 75.360 91.120 75.420 ;
        RECT 98.960 75.360 99.280 75.420 ;
        RECT 100.400 75.360 100.720 75.420 ;
        RECT 85.520 75.220 86.040 75.360 ;
        RECT 90.600 75.220 91.120 75.360 ;
        RECT 98.520 75.220 100.720 75.360 ;
        RECT 85.520 75.160 85.840 75.220 ;
        RECT 90.800 75.160 91.120 75.220 ;
        RECT 98.960 75.160 99.280 75.220 ;
        RECT 100.400 75.160 100.720 75.220 ;
      LAYER met1 ;
        RECT 115.780 75.360 116.070 75.410 ;
        RECT 118.180 75.360 118.470 75.410 ;
        RECT 123.460 75.360 123.750 75.410 ;
        RECT 115.780 75.220 123.750 75.360 ;
        RECT 115.780 75.180 116.070 75.220 ;
        RECT 118.180 75.180 118.470 75.220 ;
        RECT 123.460 75.180 123.750 75.220 ;
      LAYER met1 ;
        RECT 92.250 74.990 92.540 75.040 ;
        RECT 102.320 74.990 102.640 75.050 ;
        RECT 92.250 74.850 102.640 74.990 ;
        RECT 92.250 74.810 92.540 74.850 ;
        RECT 102.320 74.790 102.640 74.850 ;
        RECT 113.370 74.990 113.660 75.040 ;
        RECT 116.240 74.990 116.560 75.050 ;
        RECT 113.370 74.850 116.560 74.990 ;
        RECT 113.370 74.810 113.660 74.850 ;
        RECT 116.240 74.790 116.560 74.850 ;
        RECT 116.720 74.990 117.040 75.050 ;
        RECT 137.360 74.990 137.680 75.050 ;
        RECT 116.720 74.850 137.680 74.990 ;
        RECT 116.720 74.790 117.040 74.850 ;
        RECT 137.360 74.790 137.680 74.850 ;
        RECT 18.810 74.620 19.100 74.670 ;
        RECT 54.330 74.620 54.620 74.670 ;
        RECT 18.810 74.480 54.620 74.620 ;
        RECT 18.810 74.440 19.100 74.480 ;
        RECT 54.330 74.440 54.620 74.480 ;
        RECT 22.640 74.250 22.960 74.310 ;
        RECT 23.130 74.250 23.420 74.300 ;
        RECT 55.760 74.250 56.080 74.310 ;
        RECT 22.640 74.110 23.420 74.250 ;
        RECT 55.560 74.110 56.080 74.250 ;
        RECT 22.640 74.050 22.960 74.110 ;
        RECT 23.130 74.070 23.420 74.110 ;
        RECT 55.760 74.050 56.080 74.110 ;
        RECT 79.280 74.250 79.600 74.310 ;
        RECT 90.800 74.250 91.120 74.310 ;
        RECT 79.280 74.110 91.120 74.250 ;
        RECT 79.280 74.050 79.600 74.110 ;
        RECT 90.800 74.050 91.120 74.110 ;
        RECT 10.640 72.400 10.960 72.460 ;
        RECT 14.010 72.400 14.300 72.450 ;
        RECT 16.890 72.400 17.180 72.450 ;
        RECT 19.760 72.400 20.080 72.460 ;
        RECT 36.080 72.400 36.400 72.460 ;
        RECT 10.640 72.260 20.080 72.400 ;
        RECT 10.640 72.200 10.960 72.260 ;
        RECT 14.010 72.220 14.300 72.260 ;
        RECT 16.890 72.220 17.180 72.260 ;
        RECT 19.760 72.200 20.080 72.260 ;
        RECT 22.250 72.260 36.400 72.400 ;
        RECT 18.330 72.030 18.620 72.080 ;
        RECT 22.250 72.030 22.390 72.260 ;
        RECT 36.080 72.200 36.400 72.260 ;
        RECT 79.770 72.400 80.060 72.450 ;
        RECT 85.040 72.400 85.360 72.460 ;
        RECT 79.770 72.260 85.360 72.400 ;
        RECT 79.770 72.220 80.060 72.260 ;
        RECT 85.040 72.200 85.360 72.260 ;
        RECT 93.680 72.400 94.000 72.460 ;
        RECT 96.570 72.400 96.860 72.450 ;
        RECT 93.680 72.260 96.860 72.400 ;
        RECT 93.680 72.200 94.000 72.260 ;
        RECT 96.570 72.220 96.860 72.260 ;
        RECT 102.320 72.400 102.640 72.460 ;
        RECT 113.850 72.400 114.140 72.450 ;
        RECT 102.320 72.260 114.140 72.400 ;
        RECT 102.320 72.200 102.640 72.260 ;
        RECT 113.850 72.220 114.140 72.260 ;
        RECT 47.600 72.030 47.920 72.090 ;
        RECT 18.330 71.890 22.390 72.030 ;
        RECT 22.730 71.890 47.920 72.030 ;
        RECT 18.330 71.850 18.620 71.890 ;
        RECT 22.730 70.970 22.870 71.890 ;
        RECT 47.600 71.830 47.920 71.890 ;
        RECT 56.730 72.030 57.020 72.080 ;
        RECT 57.200 72.030 57.520 72.090 ;
        RECT 106.640 72.030 106.960 72.090 ;
        RECT 110.490 72.030 110.780 72.080 ;
        RECT 130.640 72.030 130.960 72.090 ;
        RECT 56.730 71.890 57.520 72.030 ;
        RECT 56.730 71.850 57.020 71.890 ;
        RECT 57.200 71.830 57.520 71.890 ;
        RECT 92.810 71.890 106.390 72.030 ;
        RECT 24.090 71.660 24.380 71.710 ;
        RECT 29.840 71.660 30.160 71.720 ;
        RECT 45.200 71.660 45.520 71.720 ;
        RECT 24.090 71.520 30.160 71.660 ;
        RECT 24.090 71.480 24.380 71.520 ;
        RECT 29.840 71.460 30.160 71.520 ;
        RECT 30.890 71.520 45.520 71.660 ;
        RECT 23.610 71.290 23.900 71.340 ;
        RECT 30.320 71.290 30.640 71.350 ;
        RECT 23.610 71.150 29.590 71.290 ;
        RECT 30.120 71.150 30.640 71.290 ;
        RECT 23.610 71.110 23.900 71.150 ;
        RECT 22.170 70.740 22.460 70.970 ;
        RECT 22.650 70.740 22.940 70.970 ;
        RECT 26.480 70.920 26.800 70.980 ;
        RECT 26.280 70.780 26.800 70.920 ;
        RECT 29.450 70.920 29.590 71.150 ;
        RECT 30.320 71.090 30.640 71.150 ;
        RECT 30.890 70.920 31.030 71.520 ;
        RECT 45.200 71.460 45.520 71.520 ;
        RECT 46.640 71.660 46.960 71.720 ;
        RECT 49.040 71.660 49.360 71.720 ;
        RECT 46.640 71.520 55.030 71.660 ;
        RECT 46.640 71.460 46.960 71.520 ;
        RECT 49.040 71.460 49.360 71.520 ;
        RECT 37.050 71.290 37.340 71.340 ;
        RECT 43.760 71.290 44.080 71.350 ;
        RECT 37.050 71.150 40.150 71.290 ;
        RECT 43.560 71.150 44.080 71.290 ;
        RECT 37.050 71.110 37.340 71.150 ;
        RECT 29.450 70.780 31.030 70.920 ;
        RECT 32.720 70.920 33.040 70.980 ;
        RECT 40.010 70.970 40.150 71.150 ;
        RECT 43.760 71.090 44.080 71.150 ;
        RECT 51.930 71.290 52.220 71.340 ;
        RECT 54.320 71.290 54.640 71.350 ;
        RECT 54.890 71.340 55.030 71.520 ;
        RECT 51.930 71.150 54.640 71.290 ;
        RECT 51.930 71.110 52.220 71.150 ;
        RECT 54.320 71.090 54.640 71.150 ;
        RECT 54.810 71.110 55.100 71.340 ;
        RECT 56.250 71.110 56.540 71.340 ;
        RECT 63.450 71.110 63.740 71.340 ;
        RECT 64.400 71.290 64.720 71.350 ;
        RECT 70.170 71.290 70.460 71.340 ;
        RECT 74.010 71.290 74.300 71.340 ;
        RECT 74.960 71.290 75.280 71.350 ;
        RECT 79.280 71.290 79.600 71.350 ;
        RECT 64.400 71.150 75.280 71.290 ;
        RECT 79.080 71.150 79.600 71.290 ;
        RECT 33.210 70.920 33.500 70.970 ;
        RECT 32.720 70.780 33.500 70.920 ;
        RECT 12.570 70.550 12.860 70.600 ;
        RECT 21.680 70.550 22.000 70.610 ;
        RECT 12.570 70.410 22.000 70.550 ;
        RECT 22.250 70.550 22.390 70.740 ;
        RECT 26.480 70.720 26.800 70.780 ;
        RECT 32.720 70.720 33.040 70.780 ;
        RECT 33.210 70.740 33.500 70.780 ;
        RECT 39.930 70.740 40.220 70.970 ;
        RECT 48.080 70.920 48.400 70.980 ;
        RECT 56.330 70.920 56.470 71.110 ;
        RECT 48.080 70.780 56.470 70.920 ;
        RECT 63.530 70.920 63.670 71.110 ;
        RECT 64.400 71.090 64.720 71.150 ;
        RECT 70.170 71.110 70.460 71.150 ;
        RECT 74.010 71.110 74.300 71.150 ;
        RECT 74.960 71.090 75.280 71.150 ;
        RECT 79.280 71.090 79.600 71.150 ;
        RECT 86.010 71.110 86.300 71.340 ;
        RECT 86.960 71.290 87.280 71.350 ;
        RECT 92.810 71.340 92.950 71.890 ;
        RECT 103.280 71.660 103.600 71.720 ;
        RECT 105.680 71.660 106.000 71.720 ;
        RECT 99.050 71.520 106.000 71.660 ;
        RECT 92.730 71.290 93.020 71.340 ;
        RECT 86.960 71.150 93.020 71.290 ;
        RECT 66.330 70.920 66.620 70.970 ;
        RECT 63.530 70.780 66.620 70.920 ;
        RECT 48.080 70.720 48.400 70.780 ;
        RECT 66.330 70.740 66.620 70.780 ;
        RECT 68.240 70.920 68.560 70.980 ;
        RECT 70.640 70.920 70.960 70.980 ;
        RECT 73.050 70.920 73.340 70.970 ;
        RECT 76.880 70.920 77.200 70.980 ;
        RECT 68.240 70.780 73.340 70.920 ;
        RECT 76.680 70.780 77.200 70.920 ;
        RECT 68.240 70.720 68.560 70.780 ;
        RECT 70.640 70.720 70.960 70.780 ;
        RECT 73.050 70.740 73.340 70.780 ;
        RECT 76.880 70.720 77.200 70.780 ;
        RECT 30.800 70.550 31.120 70.610 ;
        RECT 22.250 70.410 31.120 70.550 ;
        RECT 12.570 70.370 12.860 70.410 ;
        RECT 21.680 70.350 22.000 70.410 ;
        RECT 30.800 70.350 31.120 70.410 ;
        RECT 31.280 70.550 31.600 70.610 ;
        RECT 49.520 70.550 49.840 70.610 ;
        RECT 61.520 70.550 61.840 70.610 ;
        RECT 84.080 70.550 84.400 70.610 ;
        RECT 31.280 70.410 48.310 70.550 ;
        RECT 49.320 70.410 49.840 70.550 ;
        RECT 61.320 70.410 61.840 70.550 ;
        RECT 83.880 70.410 84.400 70.550 ;
        RECT 31.280 70.350 31.600 70.410 ;
        RECT 19.280 70.180 19.600 70.240 ;
        RECT 47.600 70.180 47.920 70.240 ;
        RECT 19.280 70.040 47.920 70.180 ;
        RECT 48.170 70.180 48.310 70.410 ;
        RECT 49.520 70.350 49.840 70.410 ;
        RECT 61.520 70.350 61.840 70.410 ;
        RECT 84.080 70.350 84.400 70.410 ;
        RECT 59.600 70.180 59.920 70.240 ;
        RECT 48.170 70.040 59.920 70.180 ;
        RECT 86.090 70.180 86.230 71.110 ;
        RECT 86.960 71.090 87.280 71.150 ;
        RECT 92.730 71.110 93.020 71.150 ;
        RECT 99.050 70.970 99.190 71.520 ;
        RECT 103.280 71.460 103.600 71.520 ;
        RECT 105.680 71.460 106.000 71.520 ;
        RECT 101.360 71.290 101.680 71.350 ;
        RECT 101.160 71.150 101.680 71.290 ;
        RECT 101.360 71.090 101.680 71.150 ;
        RECT 98.970 70.740 99.260 70.970 ;
        RECT 99.920 70.920 100.240 70.980 ;
        RECT 100.410 70.920 100.700 70.970 ;
        RECT 101.840 70.920 102.160 70.980 ;
        RECT 99.920 70.780 100.700 70.920 ;
        RECT 101.640 70.780 102.160 70.920 ;
        RECT 99.920 70.720 100.240 70.780 ;
        RECT 100.410 70.740 100.700 70.780 ;
        RECT 101.840 70.720 102.160 70.780 ;
        RECT 102.800 70.920 103.120 70.980 ;
        RECT 106.250 70.970 106.390 71.890 ;
        RECT 106.640 71.890 110.780 72.030 ;
        RECT 130.440 71.890 130.960 72.030 ;
        RECT 106.640 71.830 106.960 71.890 ;
        RECT 110.490 71.850 110.780 71.890 ;
        RECT 130.640 71.830 130.960 71.890 ;
        RECT 108.560 71.290 108.880 71.350 ;
        RECT 108.360 71.150 108.880 71.290 ;
        RECT 108.560 71.090 108.880 71.150 ;
        RECT 110.010 71.110 110.300 71.340 ;
        RECT 113.360 71.290 113.680 71.350 ;
        RECT 120.090 71.290 120.380 71.340 ;
        RECT 113.360 71.150 120.380 71.290 ;
        RECT 104.250 70.920 104.540 70.970 ;
        RECT 102.800 70.780 104.540 70.920 ;
        RECT 102.800 70.720 103.120 70.780 ;
        RECT 104.250 70.740 104.540 70.780 ;
        RECT 106.170 70.740 106.460 70.970 ;
        RECT 91.290 70.550 91.580 70.600 ;
        RECT 91.760 70.550 92.080 70.610 ;
        RECT 91.290 70.410 92.080 70.550 ;
        RECT 91.290 70.370 91.580 70.410 ;
        RECT 91.760 70.350 92.080 70.410 ;
        RECT 98.480 70.550 98.800 70.610 ;
        RECT 110.090 70.550 110.230 71.110 ;
        RECT 113.360 71.090 113.680 71.150 ;
        RECT 120.090 71.110 120.380 71.150 ;
        RECT 112.880 70.920 113.200 70.980 ;
        RECT 112.680 70.780 113.200 70.920 ;
        RECT 112.880 70.720 113.200 70.780 ;
        RECT 115.760 70.920 116.080 70.980 ;
        RECT 120.560 70.920 120.880 70.980 ;
        RECT 124.410 70.920 124.700 70.970 ;
        RECT 115.760 70.780 124.700 70.920 ;
        RECT 115.760 70.720 116.080 70.780 ;
        RECT 120.560 70.720 120.880 70.780 ;
        RECT 124.410 70.740 124.700 70.780 ;
        RECT 98.480 70.410 110.230 70.550 ;
        RECT 118.650 70.550 118.940 70.600 ;
        RECT 133.040 70.550 133.360 70.610 ;
        RECT 118.650 70.410 133.360 70.550 ;
        RECT 98.480 70.350 98.800 70.410 ;
        RECT 118.650 70.370 118.940 70.410 ;
        RECT 133.040 70.350 133.360 70.410 ;
        RECT 93.200 70.180 93.520 70.240 ;
        RECT 106.170 70.180 106.460 70.230 ;
        RECT 86.090 70.040 106.460 70.180 ;
        RECT 19.280 69.980 19.600 70.040 ;
        RECT 47.600 69.980 47.920 70.040 ;
        RECT 59.600 69.980 59.920 70.040 ;
        RECT 93.200 69.980 93.520 70.040 ;
        RECT 106.170 70.000 106.460 70.040 ;
        RECT 106.640 70.180 106.960 70.240 ;
        RECT 117.200 70.180 117.520 70.240 ;
        RECT 106.640 70.040 117.520 70.180 ;
        RECT 106.640 69.980 106.960 70.040 ;
        RECT 117.200 69.980 117.520 70.040 ;
        RECT 118.160 70.180 118.480 70.240 ;
        RECT 122.970 70.180 123.260 70.230 ;
        RECT 118.160 70.040 123.260 70.180 ;
        RECT 118.160 69.980 118.480 70.040 ;
        RECT 122.970 70.000 123.260 70.040 ;
        RECT 129.210 70.180 129.500 70.230 ;
        RECT 134.960 70.180 135.280 70.240 ;
        RECT 129.210 70.040 135.280 70.180 ;
        RECT 129.210 70.000 129.500 70.040 ;
        RECT 134.960 69.980 135.280 70.040 ;
        RECT 5.760 69.450 142.080 69.820 ;
        RECT 19.280 68.330 19.600 68.390 ;
        RECT 14.090 68.190 19.600 68.330 ;
        RECT 10.640 67.590 10.960 67.650 ;
        RECT 10.440 67.450 10.960 67.590 ;
        RECT 10.640 67.390 10.960 67.450 ;
        RECT 14.090 67.270 14.230 68.190 ;
        RECT 19.280 68.130 19.600 68.190 ;
        RECT 19.770 68.330 20.060 68.380 ;
        RECT 69.680 68.330 70.000 68.390 ;
        RECT 19.770 68.190 70.000 68.330 ;
        RECT 19.770 68.150 20.060 68.190 ;
        RECT 69.680 68.130 70.000 68.190 ;
        RECT 79.280 68.330 79.600 68.390 ;
        RECT 79.770 68.330 80.060 68.380 ;
        RECT 82.640 68.330 82.960 68.390 ;
        RECT 79.280 68.190 82.960 68.330 ;
        RECT 79.280 68.130 79.600 68.190 ;
        RECT 79.770 68.150 80.060 68.190 ;
        RECT 82.640 68.130 82.960 68.190 ;
        RECT 83.130 68.330 83.420 68.380 ;
        RECT 85.520 68.330 85.840 68.390 ;
        RECT 97.520 68.330 97.840 68.390 ;
        RECT 108.560 68.330 108.880 68.390 ;
        RECT 83.130 68.190 85.840 68.330 ;
        RECT 83.130 68.150 83.420 68.190 ;
        RECT 85.520 68.130 85.840 68.190 ;
        RECT 87.530 68.190 108.880 68.330 ;
        RECT 21.200 67.960 21.520 68.020 ;
        RECT 15.530 67.820 21.520 67.960 ;
        RECT 15.530 67.650 15.670 67.820 ;
        RECT 21.200 67.760 21.520 67.820 ;
        RECT 24.570 67.960 24.860 68.010 ;
        RECT 42.800 67.960 43.120 68.020 ;
        RECT 24.570 67.820 43.120 67.960 ;
        RECT 24.570 67.780 24.860 67.820 ;
        RECT 42.800 67.760 43.120 67.820 ;
        RECT 50.010 67.960 50.300 68.010 ;
        RECT 53.840 67.960 54.160 68.020 ;
        RECT 50.010 67.820 54.160 67.960 ;
        RECT 50.010 67.780 50.300 67.820 ;
        RECT 53.840 67.760 54.160 67.820 ;
        RECT 58.160 67.960 58.480 68.020 ;
        RECT 80.240 67.960 80.560 68.020 ;
        RECT 58.160 67.820 71.350 67.960 ;
        RECT 80.040 67.820 80.560 67.960 ;
        RECT 82.730 67.960 82.870 68.130 ;
        RECT 82.730 67.820 87.190 67.960 ;
        RECT 58.160 67.760 58.480 67.820 ;
        RECT 15.440 67.590 15.760 67.650 ;
        RECT 15.000 67.450 15.760 67.590 ;
        RECT 15.440 67.390 15.760 67.450 ;
        RECT 18.330 67.590 18.620 67.640 ;
        RECT 18.800 67.590 19.120 67.650 ;
        RECT 18.330 67.450 19.120 67.590 ;
        RECT 18.330 67.410 18.620 67.450 ;
        RECT 18.800 67.390 19.120 67.450 ;
        RECT 19.770 67.590 20.060 67.640 ;
        RECT 26.960 67.590 27.280 67.650 ;
        RECT 28.890 67.590 29.180 67.640 ;
        RECT 35.600 67.590 35.920 67.650 ;
        RECT 36.560 67.590 36.880 67.650 ;
        RECT 38.960 67.590 39.280 67.650 ;
        RECT 57.680 67.590 58.000 67.650 ;
        RECT 71.210 67.640 71.350 67.820 ;
        RECT 80.240 67.760 80.560 67.820 ;
        RECT 19.770 67.450 26.710 67.590 ;
        RECT 19.770 67.410 20.060 67.450 ;
        RECT 14.010 67.040 14.300 67.270 ;
        RECT 14.970 67.040 15.260 67.270 ;
        RECT 26.000 67.220 26.320 67.280 ;
        RECT 25.800 67.080 26.320 67.220 ;
        RECT 15.050 66.850 15.190 67.040 ;
        RECT 26.000 67.020 26.320 67.080 ;
        RECT 26.570 66.850 26.710 67.450 ;
        RECT 26.960 67.450 29.180 67.590 ;
        RECT 35.400 67.450 35.920 67.590 ;
        RECT 36.360 67.450 36.880 67.590 ;
        RECT 38.760 67.450 39.280 67.590 ;
        RECT 57.480 67.450 58.000 67.590 ;
        RECT 26.960 67.390 27.280 67.450 ;
        RECT 28.890 67.410 29.180 67.450 ;
        RECT 35.600 67.390 35.920 67.450 ;
        RECT 36.560 67.390 36.880 67.450 ;
        RECT 38.960 67.390 39.280 67.450 ;
        RECT 57.680 67.390 58.000 67.450 ;
        RECT 64.410 67.410 64.700 67.640 ;
        RECT 71.130 67.410 71.420 67.640 ;
        RECT 76.880 67.590 77.200 67.650 ;
        RECT 78.330 67.590 78.620 67.640 ;
        RECT 84.080 67.590 84.400 67.650 ;
        RECT 87.050 67.640 87.190 67.820 ;
        RECT 76.880 67.450 78.620 67.590 ;
        RECT 83.880 67.450 84.400 67.590 ;
        RECT 32.720 67.220 33.040 67.280 ;
        RECT 42.800 67.220 43.120 67.280 ;
        RECT 32.520 67.080 33.040 67.220 ;
        RECT 42.600 67.080 43.120 67.220 ;
        RECT 32.720 67.020 33.040 67.080 ;
        RECT 42.800 67.020 43.120 67.080 ;
        RECT 50.000 67.220 50.320 67.280 ;
        RECT 51.930 67.220 52.220 67.270 ;
        RECT 61.520 67.220 61.840 67.280 ;
        RECT 50.000 67.080 52.220 67.220 ;
        RECT 61.320 67.080 61.840 67.220 ;
        RECT 50.000 67.020 50.320 67.080 ;
        RECT 51.930 67.040 52.220 67.080 ;
        RECT 61.520 67.020 61.840 67.080 ;
        RECT 64.490 66.850 64.630 67.410 ;
        RECT 76.880 67.390 77.200 67.450 ;
        RECT 78.330 67.410 78.620 67.450 ;
        RECT 68.250 67.040 68.540 67.270 ;
        RECT 74.960 67.220 75.280 67.280 ;
        RECT 74.760 67.080 75.280 67.220 ;
        RECT 78.410 67.220 78.550 67.410 ;
        RECT 84.080 67.390 84.400 67.450 ;
        RECT 86.010 67.410 86.300 67.640 ;
        RECT 86.970 67.410 87.260 67.640 ;
        RECT 86.090 67.220 86.230 67.410 ;
        RECT 87.530 67.220 87.670 68.190 ;
        RECT 97.520 68.130 97.840 68.190 ;
        RECT 108.560 68.130 108.880 68.190 ;
        RECT 110.960 68.330 111.280 68.390 ;
        RECT 113.360 68.330 113.680 68.390 ;
        RECT 130.640 68.330 130.960 68.390 ;
        RECT 110.960 68.190 113.680 68.330 ;
        RECT 130.440 68.190 130.960 68.330 ;
        RECT 110.960 68.130 111.280 68.190 ;
        RECT 113.360 68.130 113.680 68.190 ;
        RECT 130.640 68.130 130.960 68.190 ;
        RECT 90.800 67.960 91.120 68.020 ;
        RECT 102.800 67.960 103.120 68.020 ;
        RECT 90.800 67.820 103.120 67.960 ;
        RECT 90.800 67.760 91.120 67.820 ;
        RECT 102.800 67.760 103.120 67.820 ;
        RECT 103.290 67.960 103.580 68.010 ;
        RECT 107.120 67.960 107.440 68.020 ;
        RECT 135.920 67.960 136.240 68.020 ;
        RECT 103.290 67.820 107.440 67.960 ;
        RECT 103.290 67.780 103.580 67.820 ;
        RECT 107.120 67.760 107.440 67.820 ;
        RECT 111.530 67.820 136.240 67.960 ;
        RECT 94.640 67.590 94.960 67.650 ;
        RECT 111.530 67.640 111.670 67.820 ;
        RECT 135.920 67.760 136.240 67.820 ;
        RECT 95.130 67.590 95.420 67.640 ;
        RECT 94.640 67.450 95.420 67.590 ;
        RECT 94.640 67.390 94.960 67.450 ;
        RECT 95.130 67.410 95.420 67.450 ;
        RECT 111.450 67.410 111.740 67.640 ;
        RECT 111.930 67.410 112.220 67.640 ;
        RECT 115.280 67.590 115.600 67.650 ;
        RECT 116.250 67.590 116.540 67.640 ;
        RECT 115.280 67.450 116.540 67.590 ;
        RECT 78.410 67.080 87.670 67.220 ;
      LAYER met1 ;
        RECT 93.700 67.220 93.990 67.270 ;
        RECT 96.100 67.220 96.390 67.270 ;
        RECT 101.380 67.220 101.670 67.270 ;
        RECT 93.700 67.080 101.670 67.220 ;
      LAYER met1 ;
        RECT 15.050 66.710 19.990 66.850 ;
        RECT 26.570 66.710 64.630 66.850 ;
        RECT 68.330 66.850 68.470 67.040 ;
        RECT 74.960 67.020 75.280 67.080 ;
      LAYER met1 ;
        RECT 93.700 67.040 93.990 67.080 ;
        RECT 96.100 67.040 96.390 67.080 ;
        RECT 101.380 67.040 101.670 67.080 ;
      LAYER met1 ;
        RECT 75.440 66.850 75.760 66.910 ;
        RECT 68.330 66.710 75.760 66.850 ;
        RECT 9.210 66.480 9.500 66.530 ;
        RECT 19.280 66.480 19.600 66.540 ;
        RECT 9.210 66.340 19.600 66.480 ;
        RECT 19.850 66.480 19.990 66.710 ;
        RECT 75.440 66.650 75.760 66.710 ;
        RECT 80.730 66.850 81.020 66.900 ;
        RECT 92.720 66.850 93.040 66.910 ;
        RECT 80.730 66.710 93.040 66.850 ;
        RECT 80.730 66.670 81.020 66.710 ;
        RECT 92.720 66.650 93.040 66.710 ;
        RECT 95.120 66.850 95.440 66.910 ;
        RECT 112.010 66.850 112.150 67.410 ;
        RECT 115.280 67.390 115.600 67.450 ;
        RECT 116.250 67.410 116.540 67.450 ;
        RECT 117.200 67.590 117.520 67.650 ;
        RECT 122.970 67.590 123.260 67.640 ;
        RECT 132.080 67.590 132.400 67.650 ;
        RECT 117.200 67.450 123.260 67.590 ;
        RECT 131.880 67.450 132.400 67.590 ;
        RECT 117.200 67.390 117.520 67.450 ;
        RECT 122.970 67.410 123.260 67.450 ;
        RECT 132.080 67.390 132.400 67.450 ;
        RECT 135.450 67.590 135.740 67.640 ;
        RECT 138.320 67.590 138.640 67.650 ;
        RECT 135.450 67.450 138.640 67.590 ;
        RECT 135.450 67.410 135.740 67.450 ;
        RECT 138.320 67.390 138.640 67.450 ;
        RECT 113.850 67.220 114.140 67.270 ;
        RECT 116.720 67.220 117.040 67.280 ;
        RECT 120.090 67.220 120.380 67.270 ;
        RECT 113.850 67.080 115.510 67.220 ;
        RECT 113.850 67.040 114.140 67.080 ;
        RECT 95.120 66.710 112.150 66.850 ;
        RECT 95.120 66.650 95.440 66.710 ;
        RECT 53.360 66.480 53.680 66.540 ;
        RECT 19.850 66.340 53.680 66.480 ;
        RECT 9.210 66.300 9.500 66.340 ;
        RECT 19.280 66.280 19.600 66.340 ;
        RECT 53.360 66.280 53.680 66.340 ;
        RECT 80.240 66.480 80.560 66.540 ;
        RECT 111.920 66.480 112.240 66.540 ;
        RECT 80.240 66.340 112.240 66.480 ;
        RECT 115.370 66.480 115.510 67.080 ;
        RECT 116.720 67.080 120.380 67.220 ;
        RECT 116.720 67.020 117.040 67.080 ;
        RECT 120.090 67.040 120.380 67.080 ;
        RECT 124.410 67.220 124.700 67.270 ;
        RECT 139.280 67.220 139.600 67.280 ;
        RECT 124.410 67.080 139.600 67.220 ;
        RECT 124.410 67.040 124.700 67.080 ;
        RECT 139.280 67.020 139.600 67.080 ;
        RECT 129.680 66.480 130.000 66.540 ;
        RECT 115.370 66.340 130.000 66.480 ;
        RECT 80.240 66.280 80.560 66.340 ;
        RECT 111.920 66.280 112.240 66.340 ;
        RECT 129.680 66.280 130.000 66.340 ;
        RECT 21.680 66.110 22.000 66.170 ;
        RECT 50.480 66.110 50.800 66.170 ;
        RECT 21.680 65.970 50.800 66.110 ;
        RECT 21.680 65.910 22.000 65.970 ;
        RECT 50.480 65.910 50.800 65.970 ;
        RECT 100.880 66.110 101.200 66.170 ;
        RECT 106.650 66.110 106.940 66.160 ;
        RECT 124.880 66.110 125.200 66.170 ;
        RECT 100.880 65.970 106.940 66.110 ;
        RECT 124.680 65.970 125.200 66.110 ;
        RECT 100.880 65.910 101.200 65.970 ;
        RECT 106.650 65.930 106.940 65.970 ;
        RECT 124.880 65.910 125.200 65.970 ;
        RECT 125.370 66.110 125.660 66.160 ;
        RECT 129.200 66.110 129.520 66.170 ;
        RECT 125.370 65.970 129.520 66.110 ;
        RECT 125.370 65.930 125.660 65.970 ;
        RECT 129.200 65.910 129.520 65.970 ;
        RECT 55.760 64.260 56.080 64.320 ;
        RECT 13.610 64.120 56.080 64.260 ;
        RECT 6.320 63.520 6.640 63.580 ;
        RECT 9.690 63.520 9.980 63.570 ;
        RECT 13.040 63.520 13.360 63.580 ;
        RECT 6.320 63.380 13.360 63.520 ;
        RECT 6.320 63.320 6.640 63.380 ;
        RECT 9.690 63.340 9.980 63.380 ;
        RECT 13.040 63.320 13.360 63.380 ;
        RECT 8.720 63.150 9.040 63.210 ;
        RECT 8.520 63.010 9.040 63.150 ;
        RECT 8.720 62.950 9.040 63.010 ;
        RECT 9.200 63.150 9.520 63.210 ;
        RECT 9.200 63.010 9.720 63.150 ;
        RECT 9.200 62.950 9.520 63.010 ;
        RECT 12.570 62.600 12.860 62.830 ;
        RECT 12.650 62.040 12.790 62.600 ;
        RECT 13.610 62.460 13.750 64.120 ;
        RECT 55.760 64.060 56.080 64.120 ;
        RECT 61.530 64.260 61.820 64.310 ;
        RECT 68.240 64.260 68.560 64.320 ;
        RECT 69.680 64.260 70.000 64.320 ;
        RECT 61.530 64.120 68.560 64.260 ;
        RECT 69.480 64.120 70.000 64.260 ;
        RECT 61.530 64.080 61.820 64.120 ;
        RECT 68.240 64.060 68.560 64.120 ;
        RECT 69.680 64.060 70.000 64.120 ;
        RECT 70.160 64.260 70.480 64.320 ;
        RECT 82.640 64.260 82.960 64.320 ;
        RECT 83.130 64.260 83.420 64.310 ;
        RECT 86.960 64.260 87.280 64.320 ;
        RECT 100.880 64.260 101.200 64.320 ;
        RECT 138.320 64.260 138.640 64.320 ;
        RECT 70.160 64.120 79.030 64.260 ;
        RECT 70.160 64.060 70.480 64.120 ;
        RECT 26.480 63.890 26.800 63.950 ;
        RECT 71.600 63.890 71.920 63.950 ;
        RECT 17.930 63.750 26.800 63.890 ;
        RECT 14.000 62.780 14.320 62.840 ;
        RECT 17.360 62.780 17.680 62.840 ;
        RECT 17.930 62.830 18.070 63.750 ;
        RECT 26.480 63.690 26.800 63.750 ;
        RECT 64.490 63.750 71.920 63.890 ;
        RECT 19.280 63.520 19.600 63.580 ;
        RECT 24.570 63.520 24.860 63.570 ;
        RECT 19.280 63.380 24.860 63.520 ;
        RECT 19.280 63.320 19.600 63.380 ;
        RECT 24.570 63.340 24.860 63.380 ;
        RECT 49.530 63.520 49.820 63.570 ;
        RECT 50.480 63.520 50.800 63.580 ;
        RECT 49.530 63.380 50.800 63.520 ;
        RECT 49.530 63.340 49.820 63.380 ;
        RECT 50.480 63.320 50.800 63.380 ;
        RECT 18.810 63.150 19.100 63.200 ;
        RECT 23.120 63.150 23.440 63.210 ;
        RECT 18.810 63.010 23.440 63.150 ;
        RECT 18.810 62.970 19.100 63.010 ;
        RECT 14.000 62.640 14.520 62.780 ;
        RECT 17.160 62.640 17.680 62.780 ;
        RECT 14.000 62.580 14.320 62.640 ;
        RECT 17.360 62.580 17.680 62.640 ;
        RECT 17.850 62.600 18.140 62.830 ;
        RECT 13.530 62.230 13.820 62.460 ;
        RECT 14.480 62.410 14.800 62.470 ;
        RECT 18.890 62.410 19.030 62.970 ;
        RECT 23.120 62.950 23.440 63.010 ;
      LAYER met1 ;
        RECT 23.620 63.160 23.910 63.200 ;
        RECT 26.020 63.160 26.310 63.200 ;
        RECT 31.300 63.160 31.590 63.200 ;
        RECT 23.620 63.020 31.590 63.160 ;
        RECT 23.620 62.970 23.910 63.020 ;
        RECT 26.020 62.970 26.310 63.020 ;
        RECT 31.300 62.970 31.590 63.020 ;
      LAYER met1 ;
        RECT 38.000 63.150 38.320 63.210 ;
        RECT 42.810 63.150 43.100 63.200 ;
        RECT 38.000 63.010 43.100 63.150 ;
        RECT 38.000 62.950 38.320 63.010 ;
        RECT 42.810 62.970 43.100 63.010 ;
      LAYER met1 ;
        RECT 48.580 63.160 48.870 63.200 ;
        RECT 50.980 63.160 51.270 63.200 ;
        RECT 56.260 63.160 56.550 63.200 ;
        RECT 48.580 63.020 56.550 63.160 ;
      LAYER met1 ;
        RECT 64.490 63.150 64.630 63.750 ;
        RECT 71.600 63.690 71.920 63.750 ;
        RECT 72.080 63.150 72.400 63.210 ;
      LAYER met1 ;
        RECT 48.580 62.970 48.870 63.020 ;
        RECT 50.980 62.970 51.270 63.020 ;
        RECT 56.260 62.970 56.550 63.020 ;
      LAYER met1 ;
        RECT 64.010 63.010 64.630 63.150 ;
        RECT 67.850 63.010 72.400 63.150 ;
        RECT 78.890 63.150 79.030 64.120 ;
        RECT 82.640 64.120 83.420 64.260 ;
        RECT 86.760 64.120 87.280 64.260 ;
        RECT 100.680 64.120 101.200 64.260 ;
        RECT 138.120 64.120 138.640 64.260 ;
        RECT 82.640 64.060 82.960 64.120 ;
        RECT 83.130 64.080 83.420 64.120 ;
        RECT 86.960 64.060 87.280 64.120 ;
        RECT 100.880 64.060 101.200 64.120 ;
        RECT 138.320 64.060 138.640 64.120 ;
        RECT 121.050 63.520 121.340 63.570 ;
        RECT 88.970 63.380 121.340 63.520 ;
        RECT 79.290 63.150 79.580 63.200 ;
        RECT 87.920 63.150 88.240 63.210 ;
        RECT 88.970 63.200 89.110 63.380 ;
        RECT 78.890 63.010 79.580 63.150 ;
        RECT 87.720 63.010 88.240 63.150 ;
        RECT 19.290 62.780 19.580 62.830 ;
        RECT 25.050 62.780 25.340 62.830 ;
        RECT 19.290 62.640 25.340 62.780 ;
        RECT 19.290 62.600 19.580 62.640 ;
        RECT 25.050 62.600 25.340 62.640 ;
        RECT 29.840 62.780 30.160 62.840 ;
        RECT 64.010 62.830 64.150 63.010 ;
        RECT 50.010 62.780 50.300 62.830 ;
        RECT 29.840 62.640 50.300 62.780 ;
        RECT 29.840 62.580 30.160 62.640 ;
        RECT 50.010 62.600 50.300 62.640 ;
        RECT 63.930 62.600 64.220 62.830 ;
        RECT 65.850 62.600 66.140 62.830 ;
        RECT 14.480 62.270 19.030 62.410 ;
        RECT 41.370 62.410 41.660 62.460 ;
        RECT 46.640 62.410 46.960 62.470 ;
        RECT 41.370 62.270 46.960 62.410 ;
        RECT 14.480 62.210 14.800 62.270 ;
        RECT 41.370 62.230 41.660 62.270 ;
        RECT 46.640 62.210 46.960 62.270 ;
        RECT 57.200 62.410 57.520 62.470 ;
        RECT 65.930 62.410 66.070 62.600 ;
        RECT 57.200 62.270 66.070 62.410 ;
        RECT 57.200 62.210 57.520 62.270 ;
        RECT 18.800 62.040 19.120 62.100 ;
        RECT 12.650 61.900 19.120 62.040 ;
        RECT 18.800 61.840 19.120 61.900 ;
        RECT 36.080 62.040 36.400 62.100 ;
        RECT 36.570 62.040 36.860 62.090 ;
        RECT 38.480 62.040 38.800 62.100 ;
        RECT 36.080 61.900 38.800 62.040 ;
        RECT 36.080 61.840 36.400 61.900 ;
        RECT 36.570 61.860 36.860 61.900 ;
        RECT 38.480 61.840 38.800 61.900 ;
        RECT 39.440 62.040 39.760 62.100 ;
        RECT 57.680 62.040 58.000 62.100 ;
        RECT 39.440 61.900 58.000 62.040 ;
        RECT 39.440 61.840 39.760 61.900 ;
        RECT 57.680 61.840 58.000 61.900 ;
        RECT 65.850 62.040 66.140 62.090 ;
        RECT 67.850 62.040 67.990 63.010 ;
        RECT 72.080 62.950 72.400 63.010 ;
        RECT 79.290 62.970 79.580 63.010 ;
        RECT 87.920 62.950 88.240 63.010 ;
        RECT 88.890 62.970 89.180 63.200 ;
        RECT 95.120 63.150 95.440 63.210 ;
        RECT 95.610 63.150 95.900 63.200 ;
        RECT 95.120 63.010 95.900 63.150 ;
        RECT 95.120 62.950 95.440 63.010 ;
        RECT 95.610 62.970 95.900 63.010 ;
        RECT 71.600 62.780 71.920 62.840 ;
        RECT 75.440 62.780 75.760 62.840 ;
        RECT 71.400 62.640 71.920 62.780 ;
        RECT 75.240 62.640 75.760 62.780 ;
        RECT 71.600 62.580 71.920 62.640 ;
        RECT 75.440 62.580 75.760 62.640 ;
        RECT 82.650 62.780 82.940 62.830 ;
        RECT 82.650 62.640 85.270 62.780 ;
        RECT 82.650 62.600 82.940 62.640 ;
        RECT 71.120 62.410 71.440 62.470 ;
        RECT 72.080 62.410 72.400 62.470 ;
        RECT 70.680 62.270 72.400 62.410 ;
        RECT 71.120 62.210 71.440 62.270 ;
        RECT 72.080 62.210 72.400 62.270 ;
        RECT 65.850 61.900 67.990 62.040 ;
        RECT 68.250 62.040 68.540 62.090 ;
        RECT 77.840 62.040 78.160 62.100 ;
        RECT 68.250 61.900 78.160 62.040 ;
        RECT 85.130 62.040 85.270 62.640 ;
        RECT 85.530 62.600 85.820 62.830 ;
        RECT 86.490 62.780 86.780 62.830 ;
        RECT 87.440 62.780 87.760 62.840 ;
        RECT 98.490 62.780 98.780 62.830 ;
        RECT 86.490 62.640 98.780 62.780 ;
        RECT 86.490 62.600 86.780 62.640 ;
        RECT 85.610 62.410 85.750 62.600 ;
        RECT 87.440 62.580 87.760 62.640 ;
        RECT 98.490 62.600 98.780 62.640 ;
        RECT 99.440 62.780 99.760 62.840 ;
        RECT 100.010 62.830 100.150 63.380 ;
        RECT 121.050 63.340 121.340 63.380 ;
      LAYER met1 ;
        RECT 108.100 63.160 108.390 63.200 ;
        RECT 110.500 63.160 110.790 63.200 ;
        RECT 115.780 63.160 116.070 63.200 ;
        RECT 108.100 63.020 116.070 63.160 ;
        RECT 108.100 62.970 108.390 63.020 ;
        RECT 110.500 62.970 110.790 63.020 ;
        RECT 115.780 62.970 116.070 63.020 ;
        RECT 125.380 63.160 125.670 63.200 ;
        RECT 127.780 63.160 128.070 63.200 ;
        RECT 133.060 63.160 133.350 63.200 ;
        RECT 125.380 63.020 133.350 63.160 ;
        RECT 125.380 62.970 125.670 63.020 ;
        RECT 127.780 62.970 128.070 63.020 ;
        RECT 133.060 62.970 133.350 63.020 ;
      LAYER met1 ;
        RECT 99.930 62.780 100.220 62.830 ;
        RECT 99.440 62.640 100.220 62.780 ;
        RECT 86.960 62.410 87.280 62.470 ;
        RECT 85.610 62.270 87.280 62.410 ;
        RECT 86.960 62.210 87.280 62.270 ;
        RECT 94.170 62.410 94.460 62.460 ;
        RECT 98.000 62.410 98.320 62.470 ;
        RECT 94.170 62.270 98.320 62.410 ;
        RECT 98.570 62.410 98.710 62.600 ;
        RECT 99.440 62.580 99.760 62.640 ;
        RECT 99.930 62.600 100.220 62.640 ;
        RECT 100.400 62.780 100.720 62.840 ;
        RECT 101.370 62.780 101.660 62.830 ;
        RECT 100.400 62.640 101.660 62.780 ;
        RECT 100.400 62.580 100.720 62.640 ;
        RECT 101.370 62.600 101.660 62.640 ;
        RECT 112.880 62.410 113.200 62.470 ;
        RECT 98.570 62.270 113.200 62.410 ;
        RECT 94.170 62.230 94.460 62.270 ;
        RECT 98.000 62.210 98.320 62.270 ;
        RECT 112.880 62.210 113.200 62.270 ;
        RECT 117.690 62.410 117.980 62.460 ;
        RECT 118.160 62.410 118.480 62.470 ;
        RECT 134.960 62.410 135.280 62.470 ;
        RECT 117.690 62.270 118.480 62.410 ;
        RECT 134.760 62.270 135.280 62.410 ;
        RECT 117.690 62.230 117.980 62.270 ;
        RECT 118.160 62.210 118.480 62.270 ;
        RECT 134.960 62.210 135.280 62.270 ;
        RECT 98.480 62.040 98.800 62.100 ;
        RECT 85.130 61.900 98.800 62.040 ;
        RECT 65.850 61.860 66.140 61.900 ;
        RECT 68.250 61.860 68.540 61.900 ;
        RECT 77.840 61.840 78.160 61.900 ;
        RECT 98.480 61.840 98.800 61.900 ;
        RECT 107.120 62.040 107.440 62.100 ;
        RECT 109.530 62.040 109.820 62.090 ;
        RECT 107.120 61.900 109.820 62.040 ;
        RECT 107.120 61.840 107.440 61.900 ;
        RECT 109.530 61.860 109.820 61.900 ;
        RECT 126.810 62.040 127.100 62.090 ;
        RECT 136.880 62.040 137.200 62.100 ;
        RECT 126.810 61.900 137.200 62.040 ;
        RECT 126.810 61.860 127.100 61.900 ;
        RECT 136.880 61.840 137.200 61.900 ;
        RECT 5.760 61.310 142.080 61.680 ;
        RECT 11.130 60.190 11.420 60.240 ;
        RECT 23.600 60.190 23.920 60.250 ;
        RECT 11.130 60.050 23.920 60.190 ;
        RECT 11.130 60.010 11.420 60.050 ;
        RECT 23.600 59.990 23.920 60.050 ;
        RECT 29.360 59.990 29.680 60.250 ;
        RECT 64.880 60.190 65.200 60.250 ;
        RECT 71.600 60.190 71.920 60.250 ;
        RECT 76.890 60.190 77.180 60.240 ;
        RECT 107.120 60.190 107.440 60.250 ;
        RECT 64.880 60.050 65.400 60.190 ;
        RECT 71.600 60.050 77.180 60.190 ;
        RECT 106.920 60.050 107.440 60.190 ;
        RECT 64.880 59.990 65.200 60.050 ;
        RECT 71.600 59.990 71.920 60.050 ;
        RECT 76.890 60.010 77.180 60.050 ;
        RECT 107.120 59.990 107.440 60.050 ;
        RECT 17.360 59.620 17.680 59.880 ;
        RECT 19.280 59.820 19.600 59.880 ;
        RECT 19.080 59.680 19.600 59.820 ;
        RECT 19.280 59.620 19.600 59.680 ;
        RECT 22.650 59.820 22.940 59.870 ;
        RECT 29.450 59.820 29.590 59.990 ;
        RECT 38.000 59.820 38.320 59.880 ;
        RECT 52.400 59.820 52.720 59.880 ;
        RECT 22.650 59.680 38.320 59.820 ;
        RECT 52.200 59.680 52.720 59.820 ;
        RECT 22.650 59.640 22.940 59.680 ;
        RECT 38.000 59.620 38.320 59.680 ;
        RECT 52.400 59.620 52.720 59.680 ;
        RECT 53.360 59.820 53.680 59.880 ;
        RECT 111.930 59.820 112.220 59.870 ;
        RECT 121.520 59.820 121.840 59.880 ;
        RECT 53.360 59.680 83.350 59.820 ;
        RECT 53.360 59.620 53.680 59.680 ;
        RECT 17.450 59.450 17.590 59.620 ;
        RECT 29.370 59.450 29.660 59.500 ;
        RECT 17.450 59.310 29.660 59.450 ;
        RECT 29.370 59.270 29.660 59.310 ;
        RECT 29.840 59.450 30.160 59.510 ;
        RECT 36.090 59.450 36.380 59.500 ;
        RECT 29.840 59.310 36.380 59.450 ;
        RECT 29.840 59.250 30.160 59.310 ;
        RECT 36.090 59.270 36.380 59.310 ;
        RECT 42.810 59.270 43.100 59.500 ;
        RECT 65.370 59.450 65.660 59.500 ;
        RECT 76.400 59.450 76.720 59.510 ;
        RECT 47.210 59.310 57.910 59.450 ;
      LAYER met1 ;
        RECT 9.700 59.080 9.990 59.130 ;
        RECT 12.100 59.080 12.390 59.130 ;
        RECT 17.380 59.080 17.670 59.130 ;
        RECT 9.700 58.940 17.670 59.080 ;
        RECT 9.700 58.900 9.990 58.940 ;
        RECT 12.100 58.900 12.390 58.940 ;
        RECT 17.380 58.900 17.670 58.940 ;
      LAYER met1 ;
        RECT 33.210 58.900 33.500 59.130 ;
        RECT 39.930 59.080 40.220 59.130 ;
        RECT 42.890 59.080 43.030 59.270 ;
        RECT 46.640 59.080 46.960 59.140 ;
        RECT 39.930 58.940 43.030 59.080 ;
        RECT 46.440 58.940 46.960 59.080 ;
        RECT 39.930 58.900 40.220 58.940 ;
        RECT 9.200 58.710 9.520 58.770 ;
        RECT 30.320 58.710 30.640 58.770 ;
        RECT 9.200 58.570 30.640 58.710 ;
        RECT 9.200 58.510 9.520 58.570 ;
        RECT 30.320 58.510 30.640 58.570 ;
        RECT 33.290 58.400 33.430 58.900 ;
        RECT 46.640 58.880 46.960 58.940 ;
        RECT 42.800 58.710 43.120 58.770 ;
        RECT 47.210 58.710 47.350 59.310 ;
        RECT 53.840 59.080 54.160 59.140 ;
        RECT 53.640 58.940 54.160 59.080 ;
        RECT 53.840 58.880 54.160 58.940 ;
        RECT 54.320 59.080 54.640 59.140 ;
        RECT 56.720 59.080 57.040 59.140 ;
        RECT 57.770 59.130 57.910 59.310 ;
        RECT 65.370 59.310 76.720 59.450 ;
        RECT 65.370 59.270 65.660 59.310 ;
        RECT 76.400 59.250 76.720 59.310 ;
        RECT 79.290 59.270 79.580 59.500 ;
        RECT 54.320 58.940 57.040 59.080 ;
        RECT 54.320 58.880 54.640 58.940 ;
        RECT 56.720 58.880 57.040 58.940 ;
        RECT 57.690 58.900 57.980 59.130 ;
      LAYER met1 ;
        RECT 63.940 59.080 64.230 59.130 ;
        RECT 66.340 59.080 66.630 59.130 ;
        RECT 71.620 59.080 71.910 59.130 ;
        RECT 63.940 58.940 71.910 59.080 ;
        RECT 63.940 58.900 64.230 58.940 ;
        RECT 66.340 58.900 66.630 58.940 ;
        RECT 71.620 58.900 71.910 58.940 ;
      LAYER met1 ;
        RECT 42.800 58.570 47.350 58.710 ;
        RECT 51.920 58.710 52.240 58.770 ;
        RECT 58.650 58.710 58.940 58.760 ;
        RECT 64.400 58.710 64.720 58.770 ;
        RECT 51.920 58.570 64.720 58.710 ;
        RECT 42.800 58.510 43.120 58.570 ;
        RECT 51.920 58.510 52.240 58.570 ;
        RECT 58.650 58.530 58.940 58.570 ;
        RECT 64.400 58.510 64.720 58.570 ;
        RECT 8.720 58.340 9.040 58.400 ;
        RECT 33.200 58.340 33.520 58.400 ;
        RECT 8.720 58.200 33.520 58.340 ;
        RECT 8.720 58.140 9.040 58.200 ;
        RECT 33.200 58.140 33.520 58.200 ;
        RECT 61.040 58.340 61.360 58.400 ;
        RECT 79.370 58.340 79.510 59.270 ;
        RECT 83.210 59.130 83.350 59.680 ;
        RECT 111.930 59.680 121.840 59.820 ;
        RECT 111.930 59.640 112.220 59.680 ;
        RECT 121.520 59.620 121.840 59.680 ;
        RECT 87.920 59.450 88.240 59.510 ;
        RECT 87.720 59.310 88.240 59.450 ;
        RECT 87.920 59.250 88.240 59.310 ;
        RECT 94.650 59.270 94.940 59.500 ;
        RECT 103.770 59.450 104.060 59.500 ;
        RECT 105.200 59.450 105.520 59.510 ;
        RECT 117.200 59.450 117.520 59.510 ;
        RECT 103.770 59.310 105.520 59.450 ;
        RECT 117.000 59.310 117.520 59.450 ;
        RECT 103.770 59.270 104.060 59.310 ;
        RECT 83.130 58.900 83.420 59.130 ;
        RECT 91.770 59.080 92.060 59.130 ;
        RECT 94.730 59.080 94.870 59.270 ;
        RECT 105.200 59.250 105.520 59.310 ;
        RECT 117.200 59.250 117.520 59.310 ;
        RECT 120.560 59.450 120.880 59.510 ;
        RECT 122.970 59.450 123.260 59.500 ;
        RECT 120.560 59.310 123.260 59.450 ;
        RECT 120.560 59.250 120.880 59.310 ;
        RECT 122.970 59.270 123.260 59.310 ;
        RECT 123.440 59.450 123.760 59.510 ;
        RECT 129.690 59.450 129.980 59.500 ;
        RECT 123.440 59.310 129.980 59.450 ;
        RECT 123.440 59.250 123.760 59.310 ;
        RECT 129.690 59.270 129.980 59.310 ;
        RECT 91.770 58.940 94.870 59.080 ;
        RECT 95.120 59.080 95.440 59.140 ;
        RECT 98.490 59.080 98.780 59.130 ;
        RECT 95.120 58.940 98.780 59.080 ;
        RECT 91.770 58.900 92.060 58.940 ;
        RECT 95.120 58.880 95.440 58.940 ;
        RECT 98.490 58.900 98.780 58.940 ;
        RECT 101.840 59.080 102.160 59.140 ;
        RECT 103.770 59.080 104.060 59.130 ;
        RECT 101.840 58.940 104.060 59.080 ;
        RECT 101.840 58.880 102.160 58.940 ;
        RECT 103.770 58.900 104.060 58.940 ;
        RECT 113.370 59.080 113.660 59.130 ;
        RECT 115.280 59.080 115.600 59.140 ;
        RECT 113.370 58.940 115.600 59.080 ;
        RECT 113.370 58.900 113.660 58.940 ;
        RECT 115.280 58.880 115.600 58.940 ;
        RECT 120.090 59.080 120.380 59.130 ;
        RECT 122.480 59.080 122.800 59.140 ;
        RECT 120.090 58.940 122.800 59.080 ;
        RECT 120.090 58.900 120.380 58.940 ;
        RECT 122.480 58.880 122.800 58.940 ;
        RECT 126.810 59.080 127.100 59.130 ;
        RECT 130.160 59.080 130.480 59.140 ;
        RECT 126.810 58.940 130.480 59.080 ;
        RECT 126.810 58.900 127.100 58.940 ;
        RECT 130.160 58.880 130.480 58.940 ;
        RECT 133.530 58.900 133.820 59.130 ;
        RECT 118.160 58.710 118.480 58.770 ;
        RECT 133.610 58.710 133.750 58.900 ;
        RECT 118.160 58.570 133.750 58.710 ;
        RECT 118.160 58.510 118.480 58.570 ;
        RECT 61.040 58.200 79.510 58.340 ;
        RECT 61.040 58.140 61.360 58.200 ;
        RECT 25.040 57.970 25.360 58.030 ;
        RECT 26.480 57.970 26.800 58.030 ;
        RECT 24.840 57.830 25.360 57.970 ;
        RECT 26.280 57.830 26.800 57.970 ;
        RECT 25.040 57.770 25.360 57.830 ;
        RECT 26.480 57.770 26.800 57.830 ;
        RECT 55.280 57.970 55.600 58.030 ;
        RECT 59.130 57.970 59.420 58.020 ;
        RECT 55.280 57.830 59.420 57.970 ;
        RECT 55.280 57.770 55.600 57.830 ;
        RECT 59.130 57.790 59.420 57.830 ;
        RECT 9.200 56.120 9.520 56.180 ;
        RECT 10.170 56.120 10.460 56.170 ;
        RECT 9.200 55.980 10.460 56.120 ;
        RECT 9.200 55.920 9.520 55.980 ;
        RECT 10.170 55.940 10.460 55.980 ;
        RECT 12.570 56.120 12.860 56.170 ;
        RECT 19.280 56.120 19.600 56.180 ;
        RECT 12.570 55.980 19.600 56.120 ;
        RECT 12.570 55.940 12.860 55.980 ;
        RECT 19.280 55.920 19.600 55.980 ;
        RECT 42.320 56.120 42.640 56.180 ;
        RECT 75.920 56.120 76.240 56.180 ;
        RECT 90.800 56.120 91.120 56.180 ;
        RECT 42.320 55.980 76.240 56.120 ;
        RECT 90.600 55.980 91.120 56.120 ;
        RECT 42.320 55.920 42.640 55.980 ;
        RECT 75.920 55.920 76.240 55.980 ;
        RECT 90.800 55.920 91.120 55.980 ;
        RECT 96.090 56.120 96.380 56.170 ;
        RECT 97.520 56.120 97.840 56.180 ;
        RECT 96.090 55.980 97.840 56.120 ;
        RECT 96.090 55.940 96.380 55.980 ;
        RECT 97.520 55.920 97.840 55.980 ;
        RECT 136.880 56.120 137.200 56.180 ;
        RECT 137.850 56.120 138.140 56.170 ;
        RECT 136.880 55.980 138.140 56.120 ;
        RECT 136.880 55.920 137.200 55.980 ;
        RECT 137.850 55.940 138.140 55.980 ;
        RECT 10.640 55.750 10.960 55.810 ;
        RECT 13.040 55.750 13.360 55.810 ;
        RECT 14.010 55.750 14.300 55.800 ;
        RECT 26.960 55.750 27.280 55.810 ;
        RECT 10.640 55.610 14.300 55.750 ;
        RECT 10.640 55.550 10.960 55.610 ;
        RECT 13.040 55.550 13.360 55.610 ;
        RECT 14.010 55.570 14.300 55.610 ;
        RECT 21.770 55.610 27.280 55.750 ;
        RECT 15.440 55.010 15.760 55.070 ;
        RECT 18.320 55.010 18.640 55.070 ;
        RECT 9.770 54.870 15.760 55.010 ;
        RECT 18.120 54.870 18.640 55.010 ;
        RECT 6.320 54.640 6.640 54.700 ;
        RECT 9.770 54.690 9.910 54.870 ;
        RECT 15.440 54.810 15.760 54.870 ;
        RECT 18.320 54.810 18.640 54.870 ;
        RECT 18.810 55.010 19.100 55.060 ;
        RECT 19.770 55.010 20.060 55.060 ;
        RECT 18.810 54.870 20.060 55.010 ;
        RECT 18.810 54.830 19.100 54.870 ;
        RECT 19.770 54.830 20.060 54.870 ;
        RECT 6.120 54.500 6.640 54.640 ;
        RECT 6.320 54.440 6.640 54.500 ;
        RECT 9.690 54.460 9.980 54.690 ;
        RECT 16.890 54.460 17.180 54.690 ;
        RECT 21.770 54.640 21.910 55.610 ;
        RECT 26.960 55.550 27.280 55.610 ;
        RECT 45.200 55.750 45.520 55.810 ;
        RECT 58.640 55.750 58.960 55.810 ;
        RECT 45.200 55.610 58.960 55.750 ;
        RECT 45.200 55.550 45.520 55.610 ;
        RECT 58.640 55.550 58.960 55.610 ;
        RECT 23.600 55.380 23.920 55.440 ;
        RECT 26.000 55.380 26.320 55.440 ;
        RECT 43.760 55.380 44.080 55.440 ;
        RECT 23.600 55.240 24.120 55.380 ;
        RECT 26.000 55.240 44.080 55.380 ;
        RECT 23.600 55.180 23.920 55.240 ;
        RECT 26.000 55.180 26.320 55.240 ;
        RECT 43.760 55.180 44.080 55.240 ;
        RECT 49.520 55.380 49.840 55.440 ;
        RECT 57.680 55.380 58.000 55.440 ;
        RECT 123.440 55.380 123.760 55.440 ;
        RECT 49.520 55.240 58.000 55.380 ;
        RECT 49.520 55.180 49.840 55.240 ;
        RECT 57.680 55.180 58.000 55.240 ;
        RECT 106.250 55.240 123.760 55.380 ;
        RECT 24.080 55.010 24.400 55.070 ;
        RECT 24.570 55.010 24.860 55.060 ;
        RECT 24.080 54.870 24.860 55.010 ;
        RECT 24.080 54.810 24.400 54.870 ;
        RECT 24.570 54.830 24.860 54.870 ;
        RECT 25.530 55.010 25.820 55.060 ;
        RECT 29.840 55.010 30.160 55.070 ;
        RECT 31.760 55.010 32.080 55.070 ;
        RECT 38.480 55.010 38.800 55.070 ;
        RECT 25.530 54.870 30.160 55.010 ;
        RECT 31.560 54.870 32.080 55.010 ;
        RECT 38.280 54.870 38.800 55.010 ;
        RECT 25.530 54.830 25.820 54.870 ;
        RECT 29.840 54.810 30.160 54.870 ;
        RECT 31.760 54.810 32.080 54.870 ;
        RECT 38.480 54.810 38.800 54.870 ;
        RECT 45.210 55.010 45.500 55.060 ;
        RECT 51.920 55.010 52.240 55.070 ;
        RECT 52.880 55.010 53.200 55.070 ;
        RECT 45.210 54.870 51.190 55.010 ;
        RECT 51.720 54.870 53.200 55.010 ;
        RECT 45.210 54.830 45.500 54.870 ;
        RECT 22.170 54.640 22.460 54.690 ;
        RECT 21.770 54.500 22.460 54.640 ;
        RECT 22.170 54.460 22.460 54.500 ;
        RECT 23.120 54.640 23.440 54.700 ;
        RECT 34.650 54.640 34.940 54.690 ;
        RECT 23.120 54.500 23.640 54.640 ;
        RECT 24.650 54.500 34.940 54.640 ;
        RECT 6.800 54.270 7.120 54.330 ;
        RECT 6.600 54.130 7.120 54.270 ;
        RECT 16.970 54.270 17.110 54.460 ;
        RECT 23.120 54.440 23.440 54.500 ;
        RECT 24.650 54.270 24.790 54.500 ;
        RECT 34.650 54.460 34.940 54.500 ;
        RECT 36.560 54.640 36.880 54.700 ;
        RECT 42.800 54.640 43.120 54.700 ;
        RECT 44.240 54.640 44.560 54.700 ;
        RECT 36.560 54.500 43.120 54.640 ;
        RECT 36.560 54.440 36.880 54.500 ;
        RECT 42.800 54.440 43.120 54.500 ;
        RECT 43.370 54.500 44.560 54.640 ;
        RECT 16.970 54.130 24.790 54.270 ;
        RECT 30.330 54.270 30.620 54.320 ;
        RECT 43.370 54.270 43.510 54.500 ;
        RECT 44.240 54.440 44.560 54.500 ;
        RECT 47.600 54.640 47.920 54.700 ;
        RECT 48.090 54.640 48.380 54.690 ;
        RECT 47.600 54.500 48.380 54.640 ;
        RECT 51.050 54.640 51.190 54.870 ;
        RECT 51.920 54.810 52.240 54.870 ;
        RECT 52.880 54.810 53.200 54.870 ;
        RECT 58.640 55.010 58.960 55.070 ;
        RECT 58.640 54.870 59.160 55.010 ;
        RECT 58.640 54.810 58.960 54.870 ;
        RECT 65.370 54.830 65.660 55.060 ;
        RECT 72.090 55.010 72.380 55.060 ;
        RECT 78.810 55.010 79.100 55.060 ;
        RECT 86.490 55.010 86.780 55.060 ;
        RECT 86.960 55.010 87.280 55.070 ;
        RECT 91.770 55.010 92.060 55.060 ;
        RECT 100.880 55.010 101.200 55.070 ;
        RECT 106.250 55.060 106.390 55.240 ;
        RECT 123.440 55.180 123.760 55.240 ;
        RECT 135.920 55.380 136.240 55.440 ;
        RECT 135.920 55.240 139.510 55.380 ;
        RECT 135.920 55.180 136.240 55.240 ;
        RECT 72.090 54.870 75.190 55.010 ;
        RECT 72.090 54.830 72.380 54.870 ;
        RECT 61.530 54.640 61.820 54.690 ;
        RECT 51.050 54.500 61.820 54.640 ;
        RECT 47.600 54.440 47.920 54.500 ;
        RECT 48.090 54.460 48.380 54.500 ;
        RECT 61.530 54.460 61.820 54.500 ;
        RECT 30.330 54.130 43.510 54.270 ;
        RECT 43.770 54.270 44.060 54.320 ;
        RECT 46.640 54.270 46.960 54.330 ;
        RECT 56.240 54.270 56.560 54.330 ;
        RECT 43.770 54.130 46.960 54.270 ;
        RECT 56.040 54.130 56.560 54.270 ;
        RECT 6.800 54.070 7.120 54.130 ;
        RECT 30.330 54.090 30.620 54.130 ;
        RECT 43.770 54.090 44.060 54.130 ;
        RECT 46.640 54.070 46.960 54.130 ;
        RECT 56.240 54.070 56.560 54.130 ;
        RECT 57.680 54.270 58.000 54.330 ;
        RECT 65.450 54.270 65.590 54.830 ;
        RECT 67.760 54.640 68.080 54.700 ;
        RECT 75.050 54.690 75.190 54.870 ;
        RECT 78.810 54.870 83.350 55.010 ;
        RECT 78.810 54.830 79.100 54.870 ;
        RECT 68.250 54.640 68.540 54.690 ;
        RECT 67.760 54.500 68.540 54.640 ;
        RECT 67.760 54.440 68.080 54.500 ;
        RECT 68.250 54.460 68.540 54.500 ;
        RECT 74.970 54.460 75.260 54.690 ;
        RECT 82.640 54.640 82.960 54.700 ;
        RECT 82.440 54.500 82.960 54.640 ;
        RECT 83.210 54.640 83.350 54.870 ;
        RECT 86.490 54.870 92.060 55.010 ;
        RECT 86.490 54.830 86.780 54.870 ;
        RECT 86.960 54.810 87.280 54.870 ;
        RECT 91.770 54.830 92.060 54.870 ;
        RECT 96.650 54.870 101.200 55.010 ;
        RECT 87.920 54.640 88.240 54.700 ;
        RECT 83.210 54.500 88.240 54.640 ;
        RECT 82.640 54.440 82.960 54.500 ;
        RECT 87.920 54.440 88.240 54.500 ;
        RECT 89.370 54.460 89.660 54.690 ;
        RECT 90.320 54.640 90.640 54.700 ;
        RECT 90.120 54.500 90.640 54.640 ;
        RECT 91.850 54.640 91.990 54.830 ;
        RECT 96.650 54.690 96.790 54.870 ;
        RECT 100.880 54.810 101.200 54.870 ;
        RECT 106.170 54.830 106.460 55.060 ;
        RECT 108.560 55.010 108.880 55.070 ;
        RECT 112.890 55.010 113.180 55.060 ;
        RECT 108.560 54.870 113.180 55.010 ;
        RECT 108.560 54.810 108.880 54.870 ;
        RECT 112.890 54.830 113.180 54.870 ;
        RECT 117.680 55.010 118.000 55.070 ;
        RECT 120.090 55.010 120.380 55.060 ;
        RECT 117.680 54.870 120.380 55.010 ;
        RECT 117.680 54.810 118.000 54.870 ;
        RECT 120.090 54.830 120.380 54.870 ;
        RECT 121.040 55.010 121.360 55.070 ;
        RECT 126.810 55.010 127.100 55.060 ;
        RECT 121.040 54.870 127.100 55.010 ;
        RECT 121.040 54.810 121.360 54.870 ;
        RECT 126.810 54.830 127.100 54.870 ;
        RECT 129.200 55.010 129.520 55.070 ;
        RECT 133.040 55.010 133.360 55.070 ;
        RECT 133.530 55.010 133.820 55.060 ;
        RECT 129.200 54.870 130.870 55.010 ;
        RECT 129.200 54.810 129.520 54.870 ;
        RECT 95.130 54.640 95.420 54.690 ;
        RECT 91.850 54.500 95.420 54.640 ;
        RECT 57.680 54.130 65.590 54.270 ;
        RECT 87.440 54.270 87.760 54.330 ;
        RECT 89.450 54.270 89.590 54.460 ;
        RECT 90.320 54.440 90.640 54.500 ;
        RECT 95.130 54.460 95.420 54.500 ;
        RECT 96.570 54.460 96.860 54.690 ;
        RECT 97.050 54.460 97.340 54.690 ;
        RECT 98.000 54.640 98.320 54.700 ;
        RECT 110.000 54.640 110.320 54.700 ;
        RECT 97.800 54.500 98.320 54.640 ;
        RECT 109.800 54.500 110.320 54.640 ;
        RECT 87.440 54.130 89.590 54.270 ;
        RECT 97.130 54.270 97.270 54.460 ;
        RECT 98.000 54.440 98.320 54.500 ;
        RECT 110.000 54.440 110.320 54.500 ;
        RECT 122.480 54.640 122.800 54.700 ;
        RECT 122.970 54.640 123.260 54.690 ;
        RECT 130.160 54.640 130.480 54.700 ;
        RECT 122.480 54.500 123.260 54.640 ;
        RECT 129.960 54.500 130.480 54.640 ;
        RECT 130.730 54.640 130.870 54.870 ;
        RECT 133.040 54.870 133.820 55.010 ;
        RECT 133.040 54.810 133.360 54.870 ;
        RECT 133.530 54.830 133.820 54.870 ;
        RECT 137.840 55.010 138.160 55.070 ;
        RECT 139.370 55.060 139.510 55.240 ;
        RECT 138.810 55.010 139.100 55.060 ;
        RECT 137.840 54.870 139.100 55.010 ;
        RECT 137.840 54.810 138.160 54.870 ;
        RECT 138.810 54.830 139.100 54.870 ;
        RECT 139.290 54.830 139.580 55.060 ;
        RECT 136.410 54.640 136.700 54.690 ;
        RECT 137.360 54.640 137.680 54.700 ;
        RECT 130.730 54.500 136.700 54.640 ;
        RECT 137.160 54.500 137.680 54.640 ;
        RECT 122.480 54.440 122.800 54.500 ;
        RECT 122.970 54.460 123.260 54.500 ;
        RECT 130.160 54.440 130.480 54.500 ;
        RECT 136.410 54.460 136.700 54.500 ;
        RECT 137.360 54.440 137.680 54.500 ;
        RECT 99.440 54.270 99.760 54.330 ;
        RECT 97.130 54.130 99.760 54.270 ;
        RECT 57.680 54.070 58.000 54.130 ;
        RECT 87.440 54.070 87.760 54.130 ;
        RECT 99.440 54.070 99.760 54.130 ;
        RECT 104.730 54.270 105.020 54.320 ;
        RECT 116.720 54.270 117.040 54.330 ;
        RECT 118.160 54.270 118.480 54.330 ;
        RECT 104.730 54.130 117.040 54.270 ;
        RECT 117.960 54.130 118.480 54.270 ;
        RECT 104.730 54.090 105.020 54.130 ;
        RECT 116.720 54.070 117.040 54.130 ;
        RECT 118.160 54.070 118.480 54.130 ;
        RECT 19.280 53.900 19.600 53.960 ;
        RECT 19.080 53.760 19.600 53.900 ;
        RECT 19.280 53.700 19.600 53.760 ;
        RECT 19.770 53.900 20.060 53.950 ;
        RECT 38.960 53.900 39.280 53.960 ;
        RECT 19.770 53.760 39.280 53.900 ;
        RECT 19.770 53.720 20.060 53.760 ;
        RECT 38.960 53.700 39.280 53.760 ;
        RECT 39.440 53.900 39.760 53.960 ;
        RECT 78.800 53.900 79.120 53.960 ;
        RECT 39.440 53.760 79.120 53.900 ;
        RECT 39.440 53.700 39.760 53.760 ;
        RECT 78.800 53.700 79.120 53.760 ;
        RECT 98.000 53.900 98.320 53.960 ;
        RECT 99.920 53.900 100.240 53.960 ;
        RECT 98.000 53.760 100.240 53.900 ;
        RECT 98.000 53.700 98.320 53.760 ;
        RECT 99.920 53.700 100.240 53.760 ;
        RECT 5.760 53.170 142.080 53.540 ;
        RECT 18.320 52.050 18.640 52.110 ;
        RECT 82.640 52.050 82.960 52.110 ;
        RECT 16.970 51.910 22.870 52.050 ;
        RECT 13.040 51.310 13.360 51.370 ;
        RECT 12.840 51.170 13.360 51.310 ;
        RECT 13.040 51.110 13.360 51.170 ;
        RECT 16.410 51.310 16.700 51.360 ;
        RECT 16.970 51.310 17.110 51.910 ;
        RECT 18.320 51.850 18.640 51.910 ;
        RECT 17.370 51.680 17.660 51.730 ;
        RECT 22.160 51.680 22.480 51.740 ;
        RECT 17.370 51.540 22.480 51.680 ;
        RECT 17.370 51.500 17.660 51.540 ;
        RECT 22.160 51.480 22.480 51.540 ;
        RECT 17.840 51.310 18.160 51.370 ;
        RECT 20.720 51.310 21.040 51.370 ;
        RECT 21.680 51.310 22.000 51.370 ;
        RECT 22.730 51.360 22.870 51.910 ;
        RECT 23.690 51.910 82.960 52.050 ;
        RECT 16.410 51.170 17.110 51.310 ;
        RECT 17.640 51.170 18.160 51.310 ;
        RECT 20.520 51.170 21.040 51.310 ;
        RECT 21.480 51.170 22.000 51.310 ;
        RECT 16.410 51.130 16.700 51.170 ;
        RECT 17.840 51.110 18.160 51.170 ;
        RECT 20.720 51.110 21.040 51.170 ;
        RECT 21.680 51.110 22.000 51.170 ;
        RECT 22.650 51.310 22.940 51.360 ;
        RECT 23.120 51.310 23.440 51.370 ;
        RECT 23.690 51.360 23.830 51.910 ;
        RECT 82.640 51.850 82.960 51.910 ;
        RECT 26.000 51.680 26.320 51.740 ;
        RECT 39.440 51.680 39.760 51.740 ;
        RECT 50.000 51.680 50.320 51.740 ;
        RECT 60.080 51.680 60.400 51.740 ;
        RECT 25.800 51.540 26.320 51.680 ;
        RECT 26.000 51.480 26.320 51.540 ;
        RECT 29.930 51.540 39.760 51.680 ;
        RECT 49.800 51.540 50.320 51.680 ;
        RECT 59.880 51.540 60.400 51.680 ;
        RECT 22.650 51.170 23.440 51.310 ;
        RECT 22.650 51.130 22.940 51.170 ;
        RECT 23.120 51.110 23.440 51.170 ;
        RECT 23.610 51.130 23.900 51.360 ;
        RECT 24.080 51.310 24.400 51.370 ;
        RECT 26.480 51.310 26.800 51.370 ;
        RECT 29.930 51.360 30.070 51.540 ;
        RECT 39.440 51.480 39.760 51.540 ;
        RECT 50.000 51.480 50.320 51.540 ;
        RECT 60.080 51.480 60.400 51.540 ;
        RECT 72.560 51.680 72.880 51.740 ;
        RECT 78.800 51.680 79.120 51.740 ;
        RECT 72.560 51.540 73.080 51.680 ;
        RECT 78.600 51.540 79.120 51.680 ;
        RECT 72.560 51.480 72.880 51.540 ;
        RECT 78.800 51.480 79.120 51.540 ;
        RECT 84.090 51.680 84.380 51.730 ;
        RECT 90.320 51.680 90.640 51.740 ;
        RECT 100.880 51.680 101.200 51.740 ;
        RECT 116.240 51.680 116.560 51.740 ;
        RECT 133.040 51.680 133.360 51.740 ;
        RECT 84.090 51.540 90.640 51.680 ;
        RECT 84.090 51.500 84.380 51.540 ;
        RECT 90.320 51.480 90.640 51.540 ;
        RECT 95.690 51.540 101.200 51.680 ;
        RECT 116.040 51.540 116.560 51.680 ;
        RECT 132.840 51.540 133.360 51.680 ;
        RECT 29.850 51.310 30.140 51.360 ;
        RECT 24.080 51.170 30.140 51.310 ;
        RECT 24.080 51.110 24.400 51.170 ;
        RECT 26.480 51.110 26.800 51.170 ;
        RECT 29.850 51.130 30.140 51.170 ;
        RECT 30.800 51.310 31.120 51.370 ;
        RECT 32.250 51.310 32.540 51.360 ;
        RECT 30.800 51.170 32.540 51.310 ;
        RECT 30.800 51.110 31.120 51.170 ;
        RECT 32.250 51.130 32.540 51.170 ;
        RECT 33.200 51.310 33.520 51.370 ;
        RECT 38.970 51.310 39.260 51.360 ;
        RECT 61.040 51.310 61.360 51.370 ;
        RECT 64.410 51.310 64.700 51.360 ;
        RECT 33.200 51.170 39.260 51.310 ;
        RECT 33.200 51.110 33.520 51.170 ;
        RECT 38.970 51.130 39.260 51.170 ;
        RECT 42.410 51.170 61.360 51.310 ;
        RECT 21.210 50.940 21.500 50.990 ;
        RECT 26.970 50.940 27.260 50.990 ;
        RECT 21.210 50.800 27.260 50.940 ;
        RECT 21.210 50.760 21.500 50.800 ;
        RECT 26.970 50.760 27.260 50.800 ;
        RECT 28.410 50.940 28.700 50.990 ;
        RECT 36.090 50.940 36.380 50.990 ;
        RECT 42.410 50.940 42.550 51.170 ;
        RECT 61.040 51.110 61.360 51.170 ;
        RECT 62.090 51.170 64.700 51.310 ;
        RECT 28.410 50.800 35.350 50.940 ;
        RECT 28.410 50.760 28.700 50.800 ;
        RECT 11.610 50.570 11.900 50.620 ;
        RECT 12.560 50.570 12.880 50.630 ;
        RECT 11.610 50.430 12.880 50.570 ;
        RECT 11.610 50.390 11.900 50.430 ;
        RECT 12.560 50.370 12.880 50.430 ;
        RECT 35.210 50.260 35.350 50.800 ;
        RECT 36.090 50.800 42.550 50.940 ;
        RECT 42.800 50.940 43.120 51.000 ;
        RECT 49.520 50.940 49.840 51.000 ;
        RECT 51.930 50.940 52.220 50.990 ;
        RECT 61.520 50.940 61.840 51.000 ;
        RECT 42.800 50.800 43.320 50.940 ;
        RECT 49.520 50.800 52.220 50.940 ;
        RECT 61.320 50.800 61.840 50.940 ;
        RECT 36.090 50.760 36.380 50.800 ;
        RECT 42.800 50.740 43.120 50.800 ;
        RECT 49.520 50.740 49.840 50.800 ;
        RECT 51.930 50.760 52.220 50.800 ;
        RECT 61.520 50.740 61.840 50.800 ;
        RECT 36.560 50.570 36.880 50.630 ;
        RECT 52.400 50.570 52.720 50.630 ;
        RECT 36.560 50.430 52.720 50.570 ;
        RECT 36.560 50.370 36.880 50.430 ;
        RECT 52.400 50.370 52.720 50.430 ;
        RECT 58.640 50.570 58.960 50.630 ;
        RECT 62.090 50.570 62.230 51.170 ;
        RECT 64.410 51.130 64.700 51.170 ;
        RECT 75.920 51.310 76.240 51.370 ;
        RECT 95.690 51.360 95.830 51.540 ;
        RECT 100.880 51.480 101.200 51.540 ;
        RECT 116.240 51.480 116.560 51.540 ;
        RECT 133.040 51.480 133.360 51.540 ;
        RECT 77.850 51.310 78.140 51.360 ;
        RECT 75.920 51.170 78.140 51.310 ;
        RECT 75.920 51.110 76.240 51.170 ;
        RECT 77.850 51.130 78.140 51.170 ;
        RECT 88.410 51.130 88.700 51.360 ;
        RECT 95.610 51.130 95.900 51.360 ;
        RECT 99.450 51.310 99.740 51.360 ;
        RECT 99.920 51.310 100.240 51.370 ;
        RECT 108.560 51.310 108.880 51.370 ;
        RECT 99.450 51.170 100.240 51.310 ;
        RECT 108.360 51.170 108.880 51.310 ;
        RECT 99.450 51.130 99.740 51.170 ;
        RECT 68.240 50.940 68.560 51.000 ;
        RECT 74.960 50.940 75.280 51.000 ;
        RECT 68.040 50.800 68.560 50.940 ;
        RECT 74.760 50.800 75.280 50.940 ;
        RECT 68.240 50.740 68.560 50.800 ;
        RECT 74.960 50.740 75.280 50.800 ;
        RECT 85.530 50.940 85.820 50.990 ;
        RECT 88.490 50.940 88.630 51.130 ;
        RECT 99.920 51.110 100.240 51.170 ;
        RECT 108.560 51.110 108.880 51.170 ;
        RECT 124.890 51.130 125.180 51.360 ;
        RECT 128.240 51.310 128.560 51.370 ;
        RECT 128.040 51.170 128.560 51.310 ;
        RECT 85.530 50.800 88.630 50.940 ;
        RECT 92.250 50.940 92.540 50.990 ;
        RECT 95.120 50.940 95.440 51.000 ;
        RECT 92.250 50.800 95.440 50.940 ;
        RECT 85.530 50.760 85.820 50.800 ;
        RECT 92.250 50.760 92.540 50.800 ;
        RECT 58.640 50.430 62.230 50.570 ;
        RECT 81.200 50.570 81.520 50.630 ;
        RECT 92.330 50.570 92.470 50.760 ;
        RECT 95.120 50.740 95.440 50.800 ;
        RECT 102.330 50.940 102.620 50.990 ;
        RECT 110.480 50.940 110.800 51.000 ;
        RECT 111.450 50.940 111.740 50.990 ;
        RECT 118.160 50.940 118.480 51.000 ;
        RECT 102.330 50.800 111.740 50.940 ;
        RECT 117.960 50.800 118.480 50.940 ;
        RECT 102.330 50.760 102.620 50.800 ;
        RECT 110.480 50.740 110.800 50.800 ;
        RECT 111.450 50.760 111.740 50.800 ;
        RECT 118.160 50.740 118.480 50.800 ;
        RECT 81.200 50.430 92.470 50.570 ;
        RECT 124.970 50.570 125.110 51.130 ;
        RECT 128.240 51.110 128.560 51.170 ;
        RECT 129.200 51.310 129.520 51.370 ;
        RECT 139.280 51.310 139.600 51.370 ;
        RECT 129.200 51.170 138.070 51.310 ;
        RECT 139.080 51.170 139.600 51.310 ;
        RECT 129.200 51.110 129.520 51.170 ;
        RECT 126.320 50.940 126.640 51.000 ;
        RECT 126.120 50.800 126.640 50.940 ;
        RECT 126.320 50.740 126.640 50.800 ;
        RECT 127.280 50.940 127.600 51.000 ;
        RECT 134.490 50.940 134.780 50.990 ;
        RECT 127.280 50.800 134.780 50.940 ;
        RECT 127.280 50.740 127.600 50.800 ;
        RECT 134.490 50.760 134.780 50.800 ;
        RECT 135.920 50.940 136.240 51.000 ;
        RECT 137.370 50.940 137.660 50.990 ;
        RECT 135.920 50.800 137.660 50.940 ;
        RECT 137.930 50.940 138.070 51.170 ;
        RECT 139.280 51.110 139.600 51.170 ;
        RECT 138.810 50.940 139.100 50.990 ;
        RECT 137.930 50.800 139.100 50.940 ;
        RECT 135.920 50.740 136.240 50.800 ;
        RECT 137.370 50.760 137.660 50.800 ;
        RECT 138.810 50.760 139.100 50.800 ;
        RECT 138.320 50.570 138.640 50.630 ;
        RECT 124.970 50.430 138.640 50.570 ;
        RECT 58.640 50.370 58.960 50.430 ;
        RECT 81.200 50.370 81.520 50.430 ;
        RECT 138.320 50.370 138.640 50.430 ;
        RECT 9.210 50.200 9.500 50.250 ;
        RECT 20.240 50.200 20.560 50.260 ;
        RECT 32.240 50.200 32.560 50.260 ;
        RECT 9.210 50.060 32.560 50.200 ;
        RECT 9.210 50.020 9.500 50.060 ;
        RECT 20.240 50.000 20.560 50.060 ;
        RECT 32.240 50.000 32.560 50.060 ;
        RECT 35.120 50.000 35.440 50.260 ;
        RECT 36.080 50.200 36.400 50.260 ;
        RECT 48.080 50.200 48.400 50.260 ;
        RECT 74.960 50.200 75.280 50.260 ;
        RECT 36.080 50.060 48.400 50.200 ;
        RECT 36.080 50.000 36.400 50.060 ;
        RECT 48.080 50.000 48.400 50.060 ;
        RECT 48.650 50.060 75.280 50.200 ;
        RECT 35.600 49.830 35.920 49.890 ;
        RECT 48.650 49.830 48.790 50.060 ;
        RECT 74.960 50.000 75.280 50.060 ;
        RECT 35.600 49.690 48.790 49.830 ;
        RECT 94.160 49.830 94.480 49.890 ;
        RECT 96.090 49.830 96.380 49.880 ;
        RECT 94.160 49.690 96.380 49.830 ;
        RECT 35.600 49.630 35.920 49.690 ;
        RECT 94.160 49.630 94.480 49.690 ;
        RECT 96.090 49.650 96.380 49.690 ;
        RECT 36.570 47.980 36.860 48.030 ;
        RECT 45.200 47.980 45.520 48.040 ;
        RECT 36.570 47.840 45.520 47.980 ;
        RECT 36.570 47.800 36.860 47.840 ;
        RECT 45.200 47.780 45.520 47.840 ;
        RECT 72.080 47.980 72.400 48.040 ;
        RECT 72.080 47.840 104.950 47.980 ;
        RECT 72.080 47.780 72.400 47.840 ;
        RECT 36.090 47.610 36.380 47.660 ;
        RECT 61.520 47.610 61.840 47.670 ;
        RECT 66.320 47.610 66.640 47.670 ;
        RECT 36.090 47.470 66.640 47.610 ;
        RECT 36.090 47.430 36.380 47.470 ;
        RECT 61.520 47.410 61.840 47.470 ;
        RECT 66.320 47.410 66.640 47.470 ;
        RECT 97.520 47.610 97.840 47.670 ;
        RECT 97.520 47.470 104.470 47.610 ;
        RECT 97.520 47.410 97.840 47.470 ;
        RECT 12.560 47.240 12.880 47.300 ;
        RECT 12.360 47.100 12.880 47.240 ;
        RECT 12.560 47.040 12.880 47.100 ;
        RECT 21.680 47.240 22.000 47.300 ;
        RECT 52.400 47.240 52.720 47.300 ;
        RECT 71.610 47.240 71.900 47.290 ;
        RECT 101.360 47.240 101.680 47.300 ;
        RECT 21.680 47.100 34.870 47.240 ;
        RECT 21.680 47.040 22.000 47.100 ;
      LAYER met1 ;
        RECT 11.620 46.880 11.910 46.920 ;
        RECT 14.020 46.880 14.310 46.920 ;
        RECT 19.300 46.880 19.590 46.920 ;
        RECT 11.620 46.740 19.590 46.880 ;
        RECT 11.620 46.690 11.910 46.740 ;
        RECT 14.020 46.690 14.310 46.740 ;
        RECT 19.300 46.690 19.590 46.740 ;
      LAYER met1 ;
        RECT 24.570 46.870 24.860 46.920 ;
        RECT 26.000 46.870 26.320 46.930 ;
        RECT 28.410 46.870 28.700 46.920 ;
        RECT 29.360 46.870 29.680 46.930 ;
        RECT 24.570 46.730 28.700 46.870 ;
        RECT 29.160 46.730 29.680 46.870 ;
        RECT 34.730 46.870 34.870 47.100 ;
        RECT 52.400 47.100 71.900 47.240 ;
        RECT 52.400 47.040 52.720 47.100 ;
        RECT 71.610 47.060 71.900 47.100 ;
        RECT 96.650 47.100 101.680 47.240 ;
        RECT 35.600 46.870 35.920 46.930 ;
        RECT 34.730 46.730 35.920 46.870 ;
        RECT 24.570 46.690 24.860 46.730 ;
        RECT 26.000 46.670 26.320 46.730 ;
        RECT 28.410 46.690 28.700 46.730 ;
        RECT 29.360 46.670 29.680 46.730 ;
        RECT 35.600 46.670 35.920 46.730 ;
        RECT 43.290 46.870 43.580 46.920 ;
        RECT 44.720 46.870 45.040 46.930 ;
        RECT 52.880 46.870 53.200 46.930 ;
        RECT 54.800 46.870 55.120 46.930 ;
        RECT 43.290 46.730 45.040 46.870 ;
        RECT 43.290 46.690 43.580 46.730 ;
        RECT 44.720 46.670 45.040 46.730 ;
        RECT 46.730 46.730 53.200 46.870 ;
        RECT 54.600 46.730 55.120 46.870 ;
        RECT 20.720 46.500 21.040 46.560 ;
        RECT 28.880 46.500 29.200 46.560 ;
        RECT 29.850 46.500 30.140 46.550 ;
        RECT 30.800 46.500 31.120 46.560 ;
        RECT 20.720 46.360 28.630 46.500 ;
        RECT 20.720 46.300 21.040 46.360 ;
        RECT 13.050 46.130 13.340 46.180 ;
        RECT 26.970 46.130 27.260 46.180 ;
        RECT 13.050 45.990 27.260 46.130 ;
        RECT 28.490 46.130 28.630 46.360 ;
        RECT 28.880 46.360 30.140 46.500 ;
        RECT 30.600 46.360 31.120 46.500 ;
        RECT 28.880 46.300 29.200 46.360 ;
        RECT 29.850 46.320 30.140 46.360 ;
        RECT 30.800 46.300 31.120 46.360 ;
        RECT 34.170 46.500 34.460 46.550 ;
        RECT 42.320 46.500 42.640 46.560 ;
        RECT 34.170 46.360 42.640 46.500 ;
        RECT 34.170 46.320 34.460 46.360 ;
        RECT 34.250 46.130 34.390 46.320 ;
        RECT 42.320 46.300 42.640 46.360 ;
        RECT 42.800 46.500 43.120 46.560 ;
        RECT 46.730 46.550 46.870 46.730 ;
        RECT 52.880 46.670 53.200 46.730 ;
        RECT 54.800 46.670 55.120 46.730 ;
        RECT 60.080 46.870 60.400 46.930 ;
        RECT 61.530 46.870 61.820 46.920 ;
        RECT 60.080 46.730 61.820 46.870 ;
        RECT 60.080 46.670 60.400 46.730 ;
        RECT 61.530 46.690 61.820 46.730 ;
        RECT 65.370 46.690 65.660 46.920 ;
        RECT 65.850 46.870 66.140 46.920 ;
        RECT 66.800 46.870 67.120 46.930 ;
        RECT 65.850 46.730 67.120 46.870 ;
        RECT 65.850 46.690 66.140 46.730 ;
        RECT 42.800 46.360 46.390 46.500 ;
        RECT 42.800 46.300 43.120 46.360 ;
        RECT 28.490 45.990 34.390 46.130 ;
        RECT 41.850 46.130 42.140 46.180 ;
        RECT 43.280 46.130 43.600 46.190 ;
        RECT 41.850 45.990 43.600 46.130 ;
        RECT 46.250 46.130 46.390 46.360 ;
        RECT 46.650 46.320 46.940 46.550 ;
        RECT 48.090 46.320 48.380 46.550 ;
        RECT 48.170 46.130 48.310 46.320 ;
        RECT 46.250 45.990 48.310 46.130 ;
        RECT 53.370 46.130 53.660 46.180 ;
        RECT 58.160 46.130 58.480 46.190 ;
        RECT 59.120 46.130 59.440 46.190 ;
        RECT 53.370 45.990 58.480 46.130 ;
        RECT 58.920 45.990 59.440 46.130 ;
        RECT 65.450 46.130 65.590 46.690 ;
        RECT 66.800 46.670 67.120 46.730 ;
      LAYER met1 ;
        RECT 70.660 46.880 70.950 46.920 ;
        RECT 73.060 46.880 73.350 46.920 ;
        RECT 78.340 46.880 78.630 46.920 ;
        RECT 70.660 46.740 78.630 46.880 ;
      LAYER met1 ;
        RECT 89.840 46.870 90.160 46.930 ;
        RECT 96.650 46.920 96.790 47.100 ;
        RECT 101.360 47.040 101.680 47.100 ;
      LAYER met1 ;
        RECT 70.660 46.690 70.950 46.740 ;
        RECT 73.060 46.690 73.350 46.740 ;
        RECT 78.340 46.690 78.630 46.740 ;
      LAYER met1 ;
        RECT 89.640 46.730 90.160 46.870 ;
        RECT 89.840 46.670 90.160 46.730 ;
        RECT 96.570 46.690 96.860 46.920 ;
        RECT 97.530 46.870 97.820 46.920 ;
        RECT 100.400 46.870 100.720 46.930 ;
        RECT 104.330 46.870 104.470 47.470 ;
        RECT 104.810 47.240 104.950 47.840 ;
        RECT 104.810 47.100 105.430 47.240 ;
        RECT 105.290 46.920 105.430 47.100 ;
        RECT 104.730 46.870 105.020 46.920 ;
        RECT 97.530 46.730 100.720 46.870 ;
        RECT 97.530 46.690 97.820 46.730 ;
        RECT 100.400 46.670 100.720 46.730 ;
        RECT 100.970 46.730 103.990 46.870 ;
        RECT 104.330 46.730 105.020 46.870 ;
        RECT 66.320 46.500 66.640 46.560 ;
        RECT 98.010 46.500 98.300 46.550 ;
        RECT 66.120 46.360 66.640 46.500 ;
        RECT 66.320 46.300 66.640 46.360 ;
        RECT 96.650 46.360 98.300 46.500 ;
        RECT 65.840 46.130 66.160 46.190 ;
        RECT 65.450 45.990 66.160 46.130 ;
        RECT 13.050 45.950 13.340 45.990 ;
        RECT 26.970 45.950 27.260 45.990 ;
        RECT 41.850 45.950 42.140 45.990 ;
        RECT 43.280 45.930 43.600 45.990 ;
        RECT 53.370 45.950 53.660 45.990 ;
        RECT 58.160 45.930 58.480 45.990 ;
        RECT 59.120 45.930 59.440 45.990 ;
        RECT 65.840 45.930 66.160 45.990 ;
        RECT 88.410 46.130 88.700 46.180 ;
        RECT 91.760 46.130 92.080 46.190 ;
        RECT 88.410 45.990 92.080 46.130 ;
        RECT 88.410 45.950 88.700 45.990 ;
        RECT 91.760 45.930 92.080 45.990 ;
        RECT 48.080 45.760 48.400 45.820 ;
        RECT 47.880 45.620 48.400 45.760 ;
        RECT 48.080 45.560 48.400 45.620 ;
        RECT 72.090 45.760 72.380 45.810 ;
        RECT 83.120 45.760 83.440 45.820 ;
        RECT 72.090 45.620 83.440 45.760 ;
        RECT 72.090 45.580 72.380 45.620 ;
        RECT 83.120 45.560 83.440 45.620 ;
        RECT 83.610 45.760 83.900 45.810 ;
        RECT 87.440 45.760 87.760 45.820 ;
        RECT 95.120 45.760 95.440 45.820 ;
        RECT 83.610 45.620 87.760 45.760 ;
        RECT 94.920 45.620 95.440 45.760 ;
        RECT 96.650 45.760 96.790 46.360 ;
        RECT 98.010 46.320 98.300 46.360 ;
        RECT 98.490 46.320 98.780 46.550 ;
        RECT 98.960 46.500 99.280 46.560 ;
        RECT 100.970 46.500 101.110 46.730 ;
        RECT 102.320 46.500 102.640 46.560 ;
        RECT 103.280 46.500 103.600 46.560 ;
        RECT 98.960 46.360 101.110 46.500 ;
        RECT 102.120 46.360 102.640 46.500 ;
        RECT 103.080 46.360 103.600 46.500 ;
        RECT 103.850 46.500 103.990 46.730 ;
        RECT 104.730 46.690 105.020 46.730 ;
        RECT 105.210 46.690 105.500 46.920 ;
        RECT 112.400 46.870 112.720 46.930 ;
        RECT 112.200 46.730 112.720 46.870 ;
        RECT 112.400 46.670 112.720 46.730 ;
        RECT 117.200 46.870 117.520 46.930 ;
        RECT 120.090 46.870 120.380 46.920 ;
        RECT 117.200 46.730 120.380 46.870 ;
        RECT 117.200 46.670 117.520 46.730 ;
        RECT 120.090 46.690 120.380 46.730 ;
      LAYER met1 ;
        RECT 126.820 46.880 127.110 46.920 ;
        RECT 129.220 46.880 129.510 46.920 ;
        RECT 134.500 46.880 134.790 46.920 ;
        RECT 126.820 46.740 134.790 46.880 ;
        RECT 126.820 46.690 127.110 46.740 ;
        RECT 129.220 46.690 129.510 46.740 ;
        RECT 134.500 46.690 134.790 46.740 ;
      LAYER met1 ;
        RECT 108.570 46.500 108.860 46.550 ;
        RECT 128.240 46.500 128.560 46.560 ;
        RECT 103.850 46.360 108.860 46.500 ;
        RECT 128.040 46.360 128.560 46.500 ;
        RECT 97.520 46.130 97.840 46.190 ;
        RECT 98.570 46.130 98.710 46.320 ;
        RECT 98.960 46.300 99.280 46.360 ;
        RECT 102.320 46.300 102.640 46.360 ;
        RECT 103.280 46.300 103.600 46.360 ;
        RECT 108.570 46.320 108.860 46.360 ;
        RECT 128.240 46.300 128.560 46.360 ;
        RECT 101.840 46.130 102.160 46.190 ;
        RECT 117.680 46.130 118.000 46.190 ;
        RECT 136.400 46.130 136.720 46.190 ;
        RECT 97.520 45.990 98.710 46.130 ;
        RECT 100.490 45.990 102.160 46.130 ;
        RECT 117.480 45.990 118.000 46.130 ;
        RECT 136.200 45.990 136.720 46.130 ;
        RECT 97.520 45.930 97.840 45.990 ;
        RECT 100.490 45.760 100.630 45.990 ;
        RECT 101.840 45.930 102.160 45.990 ;
        RECT 117.680 45.930 118.000 45.990 ;
        RECT 136.400 45.930 136.720 45.990 ;
        RECT 96.650 45.620 100.630 45.760 ;
        RECT 100.880 45.760 101.200 45.820 ;
        RECT 103.290 45.760 103.580 45.810 ;
        RECT 100.880 45.620 103.580 45.760 ;
        RECT 83.610 45.580 83.900 45.620 ;
        RECT 87.440 45.560 87.760 45.620 ;
        RECT 95.120 45.560 95.440 45.620 ;
        RECT 100.880 45.560 101.200 45.620 ;
        RECT 103.290 45.580 103.580 45.620 ;
        RECT 136.880 45.760 137.200 45.820 ;
        RECT 139.770 45.760 140.060 45.810 ;
        RECT 136.880 45.620 140.060 45.760 ;
        RECT 136.880 45.560 137.200 45.620 ;
        RECT 139.770 45.580 140.060 45.620 ;
        RECT 5.760 45.030 142.080 45.400 ;
        RECT 15.930 43.910 16.220 43.960 ;
        RECT 50.480 43.910 50.800 43.970 ;
        RECT 15.930 43.770 50.800 43.910 ;
        RECT 15.930 43.730 16.220 43.770 ;
        RECT 50.480 43.710 50.800 43.770 ;
        RECT 96.560 43.910 96.880 43.970 ;
        RECT 98.000 43.910 98.320 43.970 ;
        RECT 96.560 43.770 98.320 43.910 ;
        RECT 96.560 43.710 96.880 43.770 ;
        RECT 98.000 43.710 98.320 43.770 ;
        RECT 15.440 43.540 15.760 43.600 ;
        RECT 22.640 43.540 22.960 43.600 ;
        RECT 15.440 43.400 22.960 43.540 ;
        RECT 15.440 43.340 15.760 43.400 ;
        RECT 22.640 43.340 22.960 43.400 ;
        RECT 50.010 43.540 50.300 43.590 ;
        RECT 54.800 43.540 55.120 43.600 ;
        RECT 100.400 43.540 100.720 43.600 ;
        RECT 110.480 43.540 110.800 43.600 ;
        RECT 138.320 43.540 138.640 43.600 ;
        RECT 50.010 43.400 55.120 43.540 ;
        RECT 50.010 43.360 50.300 43.400 ;
        RECT 54.800 43.340 55.120 43.400 ;
        RECT 94.730 43.400 100.720 43.540 ;
        RECT 110.280 43.400 110.800 43.540 ;
        RECT 13.040 43.170 13.360 43.230 ;
        RECT 20.240 43.170 20.560 43.230 ;
        RECT 21.200 43.170 21.520 43.230 ;
        RECT 25.530 43.170 25.820 43.220 ;
        RECT 12.840 43.030 13.360 43.170 ;
        RECT 20.040 43.030 20.560 43.170 ;
        RECT 21.000 43.030 21.520 43.170 ;
        RECT 13.040 42.970 13.360 43.030 ;
        RECT 20.240 42.970 20.560 43.030 ;
        RECT 21.200 42.970 21.520 43.030 ;
        RECT 21.770 43.030 25.820 43.170 ;
        RECT 15.920 42.800 16.240 42.860 ;
        RECT 17.840 42.800 18.160 42.860 ;
        RECT 21.770 42.800 21.910 43.030 ;
        RECT 25.530 42.990 25.820 43.030 ;
        RECT 26.970 43.170 27.260 43.220 ;
        RECT 29.840 43.170 30.160 43.230 ;
        RECT 30.800 43.170 31.120 43.230 ;
        RECT 38.000 43.170 38.320 43.230 ;
        RECT 40.880 43.170 41.200 43.230 ;
        RECT 54.320 43.170 54.640 43.230 ;
        RECT 26.970 43.030 30.160 43.170 ;
        RECT 30.600 43.030 31.120 43.170 ;
        RECT 37.800 43.030 38.320 43.170 ;
        RECT 40.680 43.030 41.200 43.170 ;
        RECT 54.120 43.030 54.640 43.170 ;
        RECT 26.970 42.990 27.260 43.030 ;
        RECT 29.840 42.970 30.160 43.030 ;
        RECT 30.800 42.970 31.120 43.030 ;
        RECT 38.000 42.970 38.320 43.030 ;
        RECT 40.880 42.970 41.200 43.030 ;
        RECT 54.320 42.970 54.640 43.030 ;
        RECT 59.120 43.170 59.440 43.230 ;
        RECT 61.050 43.170 61.340 43.220 ;
        RECT 67.770 43.170 68.060 43.220 ;
        RECT 59.120 43.030 61.340 43.170 ;
        RECT 59.120 42.970 59.440 43.030 ;
        RECT 61.050 42.990 61.340 43.030 ;
        RECT 61.610 43.030 68.060 43.170 ;
        RECT 15.920 42.660 21.910 42.800 ;
        RECT 22.160 42.800 22.480 42.860 ;
        RECT 23.130 42.800 23.420 42.850 ;
        RECT 23.600 42.800 23.920 42.860 ;
        RECT 22.160 42.660 23.920 42.800 ;
        RECT 15.920 42.600 16.240 42.660 ;
        RECT 17.840 42.600 18.160 42.660 ;
        RECT 22.160 42.600 22.480 42.660 ;
        RECT 23.130 42.620 23.420 42.660 ;
        RECT 23.600 42.600 23.920 42.660 ;
        RECT 28.410 42.800 28.700 42.850 ;
        RECT 33.680 42.800 34.000 42.860 ;
        RECT 34.650 42.800 34.940 42.850 ;
        RECT 28.410 42.660 34.940 42.800 ;
        RECT 28.410 42.620 28.700 42.660 ;
        RECT 33.680 42.600 34.000 42.660 ;
        RECT 34.650 42.620 34.940 42.660 ;
        RECT 44.730 42.620 45.020 42.850 ;
        RECT 51.450 42.800 51.740 42.850 ;
        RECT 56.240 42.800 56.560 42.860 ;
        RECT 58.160 42.800 58.480 42.860 ;
        RECT 51.450 42.660 56.560 42.800 ;
        RECT 57.960 42.660 58.480 42.800 ;
        RECT 51.450 42.620 51.740 42.660 ;
        RECT 21.690 42.430 21.980 42.480 ;
        RECT 28.880 42.430 29.200 42.490 ;
        RECT 21.690 42.290 29.200 42.430 ;
        RECT 21.690 42.250 21.980 42.290 ;
        RECT 28.880 42.230 29.200 42.290 ;
        RECT 13.530 42.060 13.820 42.110 ;
        RECT 29.360 42.060 29.680 42.120 ;
        RECT 13.530 41.920 29.680 42.060 ;
        RECT 44.810 42.060 44.950 42.620 ;
        RECT 56.240 42.600 56.560 42.660 ;
        RECT 58.160 42.600 58.480 42.660 ;
        RECT 59.600 42.800 59.920 42.860 ;
        RECT 61.610 42.800 61.750 43.030 ;
        RECT 67.770 42.990 68.060 43.030 ;
        RECT 75.450 43.170 75.740 43.220 ;
        RECT 76.880 43.170 77.200 43.230 ;
        RECT 75.450 43.030 77.200 43.170 ;
        RECT 75.450 42.990 75.740 43.030 ;
        RECT 76.880 42.970 77.200 43.030 ;
        RECT 82.170 42.990 82.460 43.220 ;
        RECT 87.920 43.170 88.240 43.230 ;
        RECT 87.720 43.030 88.240 43.170 ;
        RECT 59.600 42.660 61.750 42.800 ;
        RECT 64.880 42.800 65.200 42.860 ;
        RECT 66.320 42.800 66.640 42.860 ;
        RECT 71.610 42.800 71.900 42.850 ;
        RECT 64.880 42.660 65.400 42.800 ;
        RECT 66.320 42.660 71.900 42.800 ;
        RECT 59.600 42.600 59.920 42.660 ;
        RECT 64.880 42.600 65.200 42.660 ;
        RECT 66.320 42.600 66.640 42.660 ;
        RECT 71.610 42.620 71.900 42.660 ;
        RECT 78.330 42.620 78.620 42.850 ;
        RECT 66.800 42.430 67.120 42.490 ;
        RECT 78.410 42.430 78.550 42.620 ;
        RECT 66.800 42.290 78.550 42.430 ;
        RECT 66.800 42.230 67.120 42.290 ;
        RECT 72.560 42.060 72.880 42.120 ;
        RECT 44.810 41.920 72.880 42.060 ;
        RECT 82.250 42.060 82.390 42.990 ;
        RECT 87.920 42.970 88.240 43.030 ;
        RECT 94.160 43.170 94.480 43.230 ;
        RECT 94.730 43.220 94.870 43.400 ;
        RECT 100.400 43.340 100.720 43.400 ;
        RECT 110.480 43.340 110.800 43.400 ;
        RECT 136.010 43.400 137.110 43.540 ;
        RECT 94.650 43.170 94.940 43.220 ;
        RECT 94.160 43.030 94.940 43.170 ;
        RECT 94.160 42.970 94.480 43.030 ;
        RECT 94.650 42.990 94.940 43.030 ;
        RECT 95.610 43.170 95.900 43.220 ;
        RECT 97.520 43.170 97.840 43.230 ;
        RECT 95.610 43.030 97.840 43.170 ;
        RECT 95.610 42.990 95.900 43.030 ;
        RECT 97.520 42.970 97.840 43.030 ;
        RECT 102.330 43.170 102.620 43.220 ;
        RECT 117.210 43.170 117.500 43.220 ;
        RECT 121.040 43.170 121.360 43.230 ;
        RECT 102.330 43.030 106.870 43.170 ;
        RECT 102.330 42.990 102.620 43.030 ;
        RECT 85.040 42.800 85.360 42.860 ;
        RECT 91.760 42.800 92.080 42.860 ;
        RECT 84.840 42.660 85.360 42.800 ;
        RECT 91.560 42.660 92.080 42.800 ;
        RECT 85.040 42.600 85.360 42.660 ;
        RECT 91.760 42.600 92.080 42.660 ;
        RECT 95.120 42.800 95.440 42.860 ;
        RECT 97.050 42.800 97.340 42.850 ;
        RECT 95.120 42.660 97.340 42.800 ;
        RECT 95.120 42.600 95.440 42.660 ;
        RECT 97.050 42.620 97.340 42.660 ;
        RECT 98.010 42.800 98.300 42.850 ;
        RECT 98.960 42.800 99.280 42.860 ;
        RECT 98.010 42.660 99.280 42.800 ;
        RECT 98.010 42.620 98.300 42.660 ;
        RECT 98.960 42.600 99.280 42.660 ;
        RECT 105.210 42.800 105.500 42.850 ;
        RECT 106.160 42.800 106.480 42.860 ;
        RECT 105.210 42.660 106.480 42.800 ;
        RECT 106.730 42.800 106.870 43.030 ;
        RECT 117.210 43.030 121.360 43.170 ;
        RECT 117.210 42.990 117.500 43.030 ;
        RECT 121.040 42.970 121.360 43.030 ;
        RECT 123.930 43.170 124.220 43.220 ;
        RECT 127.280 43.170 127.600 43.230 ;
        RECT 123.930 43.030 127.600 43.170 ;
        RECT 123.930 42.990 124.220 43.030 ;
        RECT 127.280 42.970 127.600 43.030 ;
        RECT 127.760 43.170 128.080 43.230 ;
        RECT 129.690 43.170 129.980 43.220 ;
        RECT 127.760 43.030 129.980 43.170 ;
        RECT 127.760 42.970 128.080 43.030 ;
        RECT 129.690 42.990 129.980 43.030 ;
        RECT 111.930 42.800 112.220 42.850 ;
        RECT 106.730 42.660 112.220 42.800 ;
        RECT 105.210 42.620 105.500 42.660 ;
        RECT 106.160 42.600 106.480 42.660 ;
        RECT 111.930 42.620 112.220 42.660 ;
        RECT 120.090 42.800 120.380 42.850 ;
        RECT 120.560 42.800 120.880 42.860 ;
        RECT 120.090 42.660 120.880 42.800 ;
        RECT 120.090 42.620 120.380 42.660 ;
        RECT 120.560 42.600 120.880 42.660 ;
        RECT 121.520 42.800 121.840 42.860 ;
        RECT 126.810 42.800 127.100 42.850 ;
        RECT 133.520 42.800 133.840 42.860 ;
        RECT 121.520 42.660 127.100 42.800 ;
        RECT 133.320 42.660 133.840 42.800 ;
        RECT 121.520 42.600 121.840 42.660 ;
        RECT 126.810 42.620 127.100 42.660 ;
        RECT 133.520 42.600 133.840 42.660 ;
        RECT 94.640 42.430 94.960 42.490 ;
        RECT 96.090 42.430 96.380 42.480 ;
        RECT 94.640 42.290 96.380 42.430 ;
        RECT 94.640 42.230 94.960 42.290 ;
        RECT 96.090 42.250 96.380 42.290 ;
        RECT 100.410 42.430 100.700 42.480 ;
        RECT 136.010 42.430 136.150 43.400 ;
        RECT 136.410 42.990 136.700 43.220 ;
        RECT 136.970 43.170 137.110 43.400 ;
        RECT 138.320 43.400 139.030 43.540 ;
        RECT 138.320 43.340 138.640 43.400 ;
        RECT 137.850 43.170 138.140 43.220 ;
        RECT 136.970 43.030 138.140 43.170 ;
        RECT 138.890 43.170 139.030 43.400 ;
        RECT 139.290 43.170 139.580 43.220 ;
        RECT 138.890 43.030 139.580 43.170 ;
        RECT 137.850 42.990 138.140 43.030 ;
        RECT 139.290 42.990 139.580 43.030 ;
        RECT 100.410 42.290 136.150 42.430 ;
        RECT 100.410 42.250 100.700 42.290 ;
        RECT 103.760 42.060 104.080 42.120 ;
        RECT 82.250 41.920 104.080 42.060 ;
        RECT 13.530 41.880 13.820 41.920 ;
        RECT 29.360 41.860 29.680 41.920 ;
        RECT 72.560 41.860 72.880 41.920 ;
        RECT 103.760 41.860 104.080 41.920 ;
        RECT 17.370 41.690 17.660 41.740 ;
        RECT 22.160 41.690 22.480 41.750 ;
        RECT 26.960 41.690 27.280 41.750 ;
        RECT 17.370 41.550 22.480 41.690 ;
        RECT 26.760 41.550 27.280 41.690 ;
        RECT 17.370 41.510 17.660 41.550 ;
        RECT 22.160 41.490 22.480 41.550 ;
        RECT 26.960 41.490 27.280 41.550 ;
        RECT 38.490 41.690 38.780 41.740 ;
        RECT 56.720 41.690 57.040 41.750 ;
        RECT 38.490 41.550 57.040 41.690 ;
        RECT 38.490 41.510 38.780 41.550 ;
        RECT 56.720 41.490 57.040 41.550 ;
        RECT 79.760 41.690 80.080 41.750 ;
        RECT 96.560 41.690 96.880 41.750 ;
        RECT 100.410 41.690 100.700 41.740 ;
        RECT 79.760 41.550 100.700 41.690 ;
        RECT 79.760 41.490 80.080 41.550 ;
        RECT 96.560 41.490 96.880 41.550 ;
        RECT 100.410 41.510 100.700 41.550 ;
        RECT 103.280 41.690 103.600 41.750 ;
        RECT 136.490 41.690 136.630 42.990 ;
        RECT 103.280 41.550 136.630 41.690 ;
        RECT 138.320 41.690 138.640 41.750 ;
        RECT 138.810 41.690 139.100 41.740 ;
        RECT 138.320 41.550 139.100 41.690 ;
        RECT 103.280 41.490 103.600 41.550 ;
        RECT 138.320 41.490 138.640 41.550 ;
        RECT 138.810 41.510 139.100 41.550 ;
        RECT 15.920 39.840 16.240 39.900 ;
        RECT 24.570 39.840 24.860 39.890 ;
        RECT 33.680 39.840 34.000 39.900 ;
        RECT 15.720 39.700 16.240 39.840 ;
        RECT 15.920 39.640 16.240 39.700 ;
        RECT 23.690 39.700 34.000 39.840 ;
        RECT 13.040 39.470 13.360 39.530 ;
        RECT 23.690 39.470 23.830 39.700 ;
        RECT 24.570 39.660 24.860 39.700 ;
        RECT 33.680 39.640 34.000 39.700 ;
        RECT 34.170 39.840 34.460 39.890 ;
        RECT 40.880 39.840 41.200 39.900 ;
        RECT 34.170 39.700 41.200 39.840 ;
        RECT 34.170 39.660 34.460 39.700 ;
        RECT 40.880 39.640 41.200 39.700 ;
        RECT 74.960 39.840 75.280 39.900 ;
        RECT 78.330 39.840 78.620 39.890 ;
        RECT 74.960 39.700 78.620 39.840 ;
        RECT 74.960 39.640 75.280 39.700 ;
        RECT 78.330 39.660 78.620 39.700 ;
        RECT 79.770 39.840 80.060 39.890 ;
        RECT 81.200 39.840 81.520 39.900 ;
        RECT 79.770 39.700 81.520 39.840 ;
        RECT 79.770 39.660 80.060 39.700 ;
        RECT 13.040 39.330 23.830 39.470 ;
        RECT 25.040 39.470 25.360 39.530 ;
        RECT 54.320 39.470 54.640 39.530 ;
        RECT 25.040 39.330 54.640 39.470 ;
        RECT 78.410 39.470 78.550 39.660 ;
        RECT 81.200 39.640 81.520 39.700 ;
        RECT 83.120 39.840 83.440 39.900 ;
        RECT 97.530 39.840 97.820 39.890 ;
        RECT 83.120 39.700 97.820 39.840 ;
        RECT 83.120 39.640 83.440 39.700 ;
        RECT 97.530 39.660 97.820 39.700 ;
        RECT 100.400 39.840 100.720 39.900 ;
        RECT 103.770 39.840 104.060 39.890 ;
        RECT 100.400 39.700 104.060 39.840 ;
        RECT 100.400 39.640 100.720 39.700 ;
        RECT 103.770 39.660 104.060 39.700 ;
        RECT 124.880 39.840 125.200 39.900 ;
        RECT 127.290 39.840 127.580 39.890 ;
        RECT 129.680 39.840 130.000 39.900 ;
        RECT 124.880 39.700 127.580 39.840 ;
        RECT 129.480 39.700 130.000 39.840 ;
        RECT 124.880 39.640 125.200 39.700 ;
        RECT 127.290 39.660 127.580 39.700 ;
        RECT 129.680 39.640 130.000 39.700 ;
        RECT 133.530 39.840 133.820 39.890 ;
        RECT 136.400 39.840 136.720 39.900 ;
        RECT 133.530 39.700 136.720 39.840 ;
        RECT 133.530 39.660 133.820 39.700 ;
        RECT 136.400 39.640 136.720 39.700 ;
        RECT 89.840 39.470 90.160 39.530 ;
        RECT 78.410 39.330 90.160 39.470 ;
        RECT 13.040 39.270 13.360 39.330 ;
        RECT 25.040 39.270 25.360 39.330 ;
        RECT 54.320 39.270 54.640 39.330 ;
        RECT 89.840 39.270 90.160 39.330 ;
        RECT 95.120 39.470 95.440 39.530 ;
        RECT 97.040 39.470 97.360 39.530 ;
        RECT 95.120 39.330 97.360 39.470 ;
        RECT 95.120 39.270 95.440 39.330 ;
        RECT 97.040 39.270 97.360 39.330 ;
        RECT 99.440 39.470 99.760 39.530 ;
        RECT 104.730 39.470 105.020 39.520 ;
        RECT 99.440 39.330 105.020 39.470 ;
        RECT 99.440 39.270 99.760 39.330 ;
        RECT 104.730 39.290 105.020 39.330 ;
        RECT 130.640 39.470 130.960 39.530 ;
        RECT 134.970 39.470 135.260 39.520 ;
        RECT 130.640 39.330 135.260 39.470 ;
        RECT 130.640 39.270 130.960 39.330 ;
        RECT 134.970 39.290 135.260 39.330 ;
        RECT 21.680 39.100 22.000 39.160 ;
        RECT 34.160 39.100 34.480 39.160 ;
        RECT 34.650 39.100 34.940 39.150 ;
        RECT 45.200 39.100 45.520 39.160 ;
        RECT 18.890 38.960 22.000 39.100 ;
        RECT 18.890 38.780 19.030 38.960 ;
        RECT 21.680 38.900 22.000 38.960 ;
        RECT 23.210 38.960 33.910 39.100 ;
        RECT 18.810 38.550 19.100 38.780 ;
        RECT 19.760 38.730 20.080 38.790 ;
        RECT 19.560 38.590 20.080 38.730 ;
        RECT 19.760 38.530 20.080 38.590 ;
        RECT 20.250 38.730 20.540 38.780 ;
        RECT 23.210 38.730 23.350 38.960 ;
        RECT 20.250 38.590 23.350 38.730 ;
        RECT 20.250 38.550 20.540 38.590 ;
        RECT 23.610 38.550 23.900 38.780 ;
        RECT 24.090 38.550 24.380 38.780 ;
        RECT 28.400 38.730 28.720 38.790 ;
        RECT 28.200 38.590 28.720 38.730 ;
        RECT 15.450 38.180 15.740 38.410 ;
        RECT 15.530 37.620 15.670 38.180 ;
        RECT 23.690 37.990 23.830 38.550 ;
        RECT 24.170 38.360 24.310 38.550 ;
        RECT 28.400 38.530 28.720 38.590 ;
        RECT 28.890 38.730 29.180 38.780 ;
        RECT 31.760 38.730 32.080 38.790 ;
        RECT 33.200 38.730 33.520 38.790 ;
        RECT 28.890 38.590 32.080 38.730 ;
        RECT 33.000 38.590 33.520 38.730 ;
        RECT 33.770 38.730 33.910 38.960 ;
        RECT 34.160 38.960 34.940 39.100 ;
        RECT 34.160 38.900 34.480 38.960 ;
        RECT 34.650 38.920 34.940 38.960 ;
        RECT 40.970 38.960 45.520 39.100 ;
        RECT 40.970 38.730 41.110 38.960 ;
        RECT 45.200 38.900 45.520 38.960 ;
        RECT 53.450 38.960 68.470 39.100 ;
        RECT 33.770 38.590 41.110 38.730 ;
        RECT 41.370 38.730 41.660 38.780 ;
        RECT 48.080 38.730 48.400 38.790 ;
        RECT 41.370 38.590 47.350 38.730 ;
        RECT 47.880 38.590 48.400 38.730 ;
        RECT 28.890 38.550 29.180 38.590 ;
        RECT 31.760 38.530 32.080 38.590 ;
        RECT 33.200 38.530 33.520 38.590 ;
        RECT 41.370 38.550 41.660 38.590 ;
        RECT 25.040 38.360 25.360 38.420 ;
        RECT 24.170 38.220 25.360 38.360 ;
        RECT 25.040 38.160 25.360 38.220 ;
        RECT 26.000 38.360 26.320 38.420 ;
        RECT 26.970 38.360 27.260 38.410 ;
        RECT 26.000 38.220 27.260 38.360 ;
        RECT 26.000 38.160 26.320 38.220 ;
        RECT 26.970 38.180 27.260 38.220 ;
        RECT 29.840 38.360 30.160 38.420 ;
        RECT 32.250 38.360 32.540 38.410 ;
        RECT 36.080 38.360 36.400 38.420 ;
        RECT 44.720 38.360 45.040 38.420 ;
        RECT 29.840 38.220 36.400 38.360 ;
        RECT 44.520 38.220 45.040 38.360 ;
        RECT 47.210 38.360 47.350 38.590 ;
        RECT 48.080 38.530 48.400 38.590 ;
        RECT 47.210 38.220 50.710 38.360 ;
        RECT 29.840 38.160 30.160 38.220 ;
        RECT 32.250 38.180 32.540 38.220 ;
        RECT 36.080 38.160 36.400 38.220 ;
        RECT 44.720 38.160 45.040 38.220 ;
        RECT 38.480 37.990 38.800 38.050 ;
        RECT 23.690 37.850 38.800 37.990 ;
        RECT 38.480 37.790 38.800 37.850 ;
        RECT 39.930 37.990 40.220 38.040 ;
        RECT 50.000 37.990 50.320 38.050 ;
        RECT 39.930 37.850 50.320 37.990 ;
        RECT 39.930 37.810 40.220 37.850 ;
        RECT 50.000 37.790 50.320 37.850 ;
        RECT 26.000 37.620 26.320 37.680 ;
        RECT 29.360 37.620 29.680 37.680 ;
        RECT 15.530 37.480 26.320 37.620 ;
        RECT 29.160 37.480 29.680 37.620 ;
        RECT 26.000 37.420 26.320 37.480 ;
        RECT 29.360 37.420 29.680 37.480 ;
        RECT 33.200 37.620 33.520 37.680 ;
        RECT 40.400 37.620 40.720 37.680 ;
        RECT 33.200 37.480 40.720 37.620 ;
        RECT 50.570 37.620 50.710 38.220 ;
        RECT 53.450 38.040 53.590 38.960 ;
        RECT 54.810 38.730 55.100 38.780 ;
        RECT 59.600 38.730 59.920 38.790 ;
        RECT 68.330 38.780 68.470 38.960 ;
        RECT 54.810 38.590 59.920 38.730 ;
        RECT 54.810 38.550 55.100 38.590 ;
        RECT 59.600 38.530 59.920 38.590 ;
        RECT 61.530 38.730 61.820 38.780 ;
        RECT 61.530 38.590 64.630 38.730 ;
        RECT 61.530 38.550 61.820 38.590 ;
        RECT 57.680 38.360 58.000 38.420 ;
        RECT 64.490 38.410 64.630 38.590 ;
        RECT 68.250 38.550 68.540 38.780 ;
        RECT 68.720 38.730 69.040 38.790 ;
        RECT 74.970 38.730 75.260 38.780 ;
        RECT 68.720 38.590 75.260 38.730 ;
        RECT 68.720 38.530 69.040 38.590 ;
        RECT 74.970 38.550 75.260 38.590 ;
        RECT 86.490 38.730 86.780 38.780 ;
        RECT 86.960 38.730 87.280 38.790 ;
        RECT 86.490 38.590 87.280 38.730 ;
        RECT 89.930 38.730 90.070 39.270 ;
        RECT 97.520 39.100 97.840 39.160 ;
        RECT 98.960 39.100 99.280 39.160 ;
        RECT 96.650 38.960 99.280 39.100 ;
        RECT 93.210 38.730 93.500 38.780 ;
        RECT 89.930 38.590 93.500 38.730 ;
        RECT 86.490 38.550 86.780 38.590 ;
        RECT 86.960 38.530 87.280 38.590 ;
        RECT 93.210 38.550 93.500 38.590 ;
        RECT 57.480 38.220 58.000 38.360 ;
        RECT 57.680 38.160 58.000 38.220 ;
        RECT 64.410 38.180 64.700 38.410 ;
        RECT 64.880 38.360 65.200 38.420 ;
        RECT 71.130 38.360 71.420 38.410 ;
        RECT 64.880 38.220 71.420 38.360 ;
        RECT 64.880 38.160 65.200 38.220 ;
        RECT 71.130 38.180 71.420 38.220 ;
        RECT 85.040 38.360 85.360 38.420 ;
        RECT 89.370 38.360 89.660 38.410 ;
        RECT 85.040 38.220 89.660 38.360 ;
        RECT 85.040 38.160 85.360 38.220 ;
        RECT 89.370 38.180 89.660 38.220 ;
        RECT 96.090 38.360 96.380 38.410 ;
        RECT 96.650 38.360 96.790 38.960 ;
        RECT 97.520 38.900 97.840 38.960 ;
        RECT 98.960 38.900 99.280 38.960 ;
        RECT 101.360 39.100 101.680 39.160 ;
        RECT 108.090 39.100 108.380 39.150 ;
        RECT 101.360 38.960 108.380 39.100 ;
        RECT 101.360 38.900 101.680 38.960 ;
        RECT 98.000 38.730 98.320 38.790 ;
        RECT 98.490 38.730 98.780 38.780 ;
        RECT 98.000 38.590 98.780 38.730 ;
        RECT 98.000 38.530 98.320 38.590 ;
        RECT 98.490 38.550 98.780 38.590 ;
        RECT 99.450 38.730 99.740 38.780 ;
        RECT 102.320 38.730 102.640 38.790 ;
        RECT 99.450 38.590 102.640 38.730 ;
        RECT 99.450 38.550 99.740 38.590 ;
        RECT 102.320 38.530 102.640 38.590 ;
        RECT 96.090 38.220 96.790 38.360 ;
        RECT 97.050 38.360 97.340 38.410 ;
        RECT 100.880 38.360 101.200 38.420 ;
        RECT 97.050 38.220 101.200 38.360 ;
        RECT 96.090 38.180 96.380 38.220 ;
        RECT 97.050 38.180 97.340 38.220 ;
        RECT 100.880 38.160 101.200 38.220 ;
        RECT 101.850 38.360 102.140 38.410 ;
        RECT 102.890 38.360 103.030 38.960 ;
        RECT 108.090 38.920 108.380 38.960 ;
        RECT 136.400 39.100 136.720 39.160 ;
        RECT 138.320 39.100 138.640 39.160 ;
        RECT 136.400 38.960 138.640 39.100 ;
        RECT 136.400 38.900 136.720 38.960 ;
        RECT 138.320 38.900 138.640 38.960 ;
        RECT 112.400 38.730 112.720 38.790 ;
        RECT 114.810 38.730 115.100 38.780 ;
        RECT 124.400 38.730 124.720 38.790 ;
        RECT 112.400 38.590 124.720 38.730 ;
        RECT 112.400 38.530 112.720 38.590 ;
        RECT 114.810 38.550 115.100 38.590 ;
        RECT 124.400 38.530 124.720 38.590 ;
        RECT 128.730 38.730 129.020 38.780 ;
        RECT 129.200 38.730 129.520 38.790 ;
        RECT 135.920 38.730 136.240 38.790 ;
        RECT 128.730 38.590 129.520 38.730 ;
        RECT 128.730 38.550 129.020 38.590 ;
        RECT 101.850 38.220 103.030 38.360 ;
        RECT 104.730 38.360 105.020 38.410 ;
        RECT 107.130 38.360 107.420 38.410 ;
        RECT 104.730 38.220 107.420 38.360 ;
        RECT 101.850 38.180 102.140 38.220 ;
        RECT 104.730 38.180 105.020 38.220 ;
        RECT 107.130 38.180 107.420 38.220 ;
        RECT 108.080 38.360 108.400 38.420 ;
        RECT 110.970 38.360 111.260 38.410 ;
        RECT 108.080 38.220 111.260 38.360 ;
        RECT 108.080 38.160 108.400 38.220 ;
        RECT 110.970 38.180 111.260 38.220 ;
        RECT 123.440 38.360 123.760 38.420 ;
        RECT 128.810 38.360 128.950 38.550 ;
        RECT 129.200 38.530 129.520 38.590 ;
        RECT 131.210 38.590 136.240 38.730 ;
        RECT 131.210 38.410 131.350 38.590 ;
        RECT 135.920 38.530 136.240 38.590 ;
        RECT 123.440 38.220 128.950 38.360 ;
        RECT 123.440 38.160 123.760 38.220 ;
        RECT 131.130 38.180 131.420 38.410 ;
        RECT 53.370 37.810 53.660 38.040 ;
        RECT 84.570 37.990 84.860 38.040 ;
        RECT 101.360 37.990 101.680 38.050 ;
        RECT 122.960 37.990 123.280 38.050 ;
        RECT 84.570 37.850 101.680 37.990 ;
        RECT 122.760 37.850 123.280 37.990 ;
        RECT 84.570 37.810 84.860 37.850 ;
        RECT 101.360 37.790 101.680 37.850 ;
        RECT 122.960 37.790 123.280 37.850 ;
        RECT 57.200 37.620 57.520 37.680 ;
        RECT 50.570 37.480 57.520 37.620 ;
        RECT 33.200 37.420 33.520 37.480 ;
        RECT 40.400 37.420 40.720 37.480 ;
        RECT 57.200 37.420 57.520 37.480 ;
        RECT 99.440 37.620 99.760 37.680 ;
        RECT 104.250 37.620 104.540 37.670 ;
        RECT 99.440 37.480 104.540 37.620 ;
        RECT 99.440 37.420 99.760 37.480 ;
        RECT 104.250 37.440 104.540 37.480 ;
        RECT 5.760 36.890 142.080 37.260 ;
        RECT 57.680 35.770 58.000 35.830 ;
        RECT 10.730 35.630 58.000 35.770 ;
        RECT 10.730 35.080 10.870 35.630 ;
        RECT 57.680 35.570 58.000 35.630 ;
        RECT 97.050 35.770 97.340 35.820 ;
        RECT 98.480 35.770 98.800 35.830 ;
        RECT 97.050 35.630 98.800 35.770 ;
        RECT 97.050 35.590 97.340 35.630 ;
        RECT 98.480 35.570 98.800 35.630 ;
        RECT 103.280 35.770 103.600 35.830 ;
        RECT 111.920 35.770 112.240 35.830 ;
        RECT 112.410 35.770 112.700 35.820 ;
        RECT 103.280 35.630 106.390 35.770 ;
        RECT 103.280 35.570 103.600 35.630 ;
        RECT 22.650 35.220 22.940 35.450 ;
        RECT 29.840 35.400 30.160 35.460 ;
        RECT 25.610 35.260 30.160 35.400 ;
        RECT 10.650 34.850 10.940 35.080 ;
        RECT 21.680 35.030 22.000 35.090 ;
        RECT 21.480 34.890 22.000 35.030 ;
        RECT 21.680 34.830 22.000 34.890 ;
        RECT 22.730 34.290 22.870 35.220 ;
        RECT 25.610 35.080 25.750 35.260 ;
        RECT 29.840 35.200 30.160 35.260 ;
        RECT 50.010 35.400 50.300 35.450 ;
        RECT 60.560 35.400 60.880 35.460 ;
        RECT 106.250 35.450 106.390 35.630 ;
        RECT 111.920 35.630 112.700 35.770 ;
        RECT 111.920 35.570 112.240 35.630 ;
        RECT 112.410 35.590 112.700 35.630 ;
        RECT 115.770 35.770 116.060 35.820 ;
        RECT 123.440 35.770 123.760 35.830 ;
        RECT 124.400 35.770 124.720 35.830 ;
        RECT 126.320 35.770 126.640 35.830 ;
        RECT 115.770 35.630 123.760 35.770 ;
        RECT 123.960 35.630 125.590 35.770 ;
        RECT 126.120 35.630 126.640 35.770 ;
        RECT 115.770 35.590 116.060 35.630 ;
        RECT 123.440 35.570 123.760 35.630 ;
        RECT 50.010 35.260 60.880 35.400 ;
        RECT 50.010 35.220 50.300 35.260 ;
        RECT 60.560 35.200 60.880 35.260 ;
        RECT 84.090 35.400 84.380 35.450 ;
        RECT 84.090 35.260 97.270 35.400 ;
        RECT 84.090 35.220 84.380 35.260 ;
        RECT 23.130 35.030 23.420 35.080 ;
        RECT 25.530 35.030 25.820 35.080 ;
        RECT 26.480 35.030 26.800 35.090 ;
        RECT 34.170 35.030 34.460 35.080 ;
        RECT 35.120 35.030 35.440 35.090 ;
        RECT 23.130 34.890 25.820 35.030 ;
        RECT 26.280 34.890 26.800 35.030 ;
        RECT 23.130 34.850 23.420 34.890 ;
        RECT 25.530 34.850 25.820 34.890 ;
        RECT 26.480 34.830 26.800 34.890 ;
        RECT 27.050 34.890 34.460 35.030 ;
        RECT 34.680 34.890 35.440 35.030 ;
        RECT 23.600 34.660 23.920 34.720 ;
        RECT 27.050 34.660 27.190 34.890 ;
        RECT 34.170 34.850 34.460 34.890 ;
        RECT 35.120 34.830 35.440 34.890 ;
        RECT 41.850 35.030 42.140 35.080 ;
        RECT 54.320 35.030 54.640 35.090 ;
        RECT 41.850 34.890 43.030 35.030 ;
        RECT 54.120 34.890 54.640 35.030 ;
        RECT 41.850 34.850 42.140 34.890 ;
        RECT 23.600 34.520 27.190 34.660 ;
        RECT 23.600 34.460 23.920 34.520 ;
        RECT 27.930 34.480 28.220 34.710 ;
        RECT 28.880 34.660 29.200 34.720 ;
        RECT 32.720 34.660 33.040 34.720 ;
        RECT 28.680 34.520 29.200 34.660 ;
        RECT 32.520 34.520 33.040 34.660 ;
        RECT 28.010 34.290 28.150 34.480 ;
        RECT 28.880 34.460 29.200 34.520 ;
        RECT 32.720 34.460 33.040 34.520 ;
        RECT 33.690 34.480 33.980 34.710 ;
        RECT 35.210 34.660 35.350 34.830 ;
        RECT 42.320 34.660 42.640 34.720 ;
        RECT 35.210 34.520 42.640 34.660 ;
        RECT 31.290 34.290 31.580 34.340 ;
        RECT 22.730 34.150 27.670 34.290 ;
        RECT 28.010 34.150 31.580 34.290 ;
        RECT 33.770 34.290 33.910 34.480 ;
        RECT 42.320 34.460 42.640 34.520 ;
        RECT 35.600 34.290 35.920 34.350 ;
        RECT 33.770 34.150 35.920 34.290 ;
        RECT 42.890 34.290 43.030 34.890 ;
        RECT 54.320 34.830 54.640 34.890 ;
        RECT 64.410 35.030 64.700 35.080 ;
        RECT 66.320 35.030 66.640 35.090 ;
        RECT 78.800 35.030 79.120 35.090 ;
        RECT 64.410 34.890 66.640 35.030 ;
        RECT 78.600 34.890 79.120 35.030 ;
        RECT 64.410 34.850 64.700 34.890 ;
        RECT 66.320 34.830 66.640 34.890 ;
        RECT 78.800 34.830 79.120 34.890 ;
        RECT 90.330 35.030 90.620 35.080 ;
        RECT 94.640 35.030 94.960 35.090 ;
        RECT 97.130 35.080 97.270 35.260 ;
        RECT 105.210 35.220 105.500 35.450 ;
        RECT 106.170 35.220 106.460 35.450 ;
        RECT 106.640 35.400 106.960 35.460 ;
        RECT 124.010 35.450 124.150 35.630 ;
        RECT 124.400 35.570 124.720 35.630 ;
        RECT 106.640 35.260 122.230 35.400 ;
        RECT 96.090 35.030 96.380 35.080 ;
        RECT 90.330 34.890 94.390 35.030 ;
        RECT 90.330 34.850 90.620 34.890 ;
        RECT 44.720 34.660 45.040 34.720 ;
        RECT 51.440 34.660 51.760 34.720 ;
        RECT 44.520 34.520 45.040 34.660 ;
        RECT 51.240 34.520 51.760 34.660 ;
        RECT 44.720 34.460 45.040 34.520 ;
        RECT 51.440 34.460 51.760 34.520 ;
        RECT 58.170 34.660 58.460 34.710 ;
        RECT 59.120 34.660 59.440 34.720 ;
        RECT 58.170 34.520 59.440 34.660 ;
        RECT 58.170 34.480 58.460 34.520 ;
        RECT 59.120 34.460 59.440 34.520 ;
      LAYER met1 ;
        RECT 62.980 34.660 63.270 34.710 ;
        RECT 65.380 34.660 65.670 34.710 ;
        RECT 70.660 34.660 70.950 34.710 ;
        RECT 62.980 34.520 70.950 34.660 ;
        RECT 62.980 34.480 63.270 34.520 ;
        RECT 65.380 34.480 65.670 34.520 ;
        RECT 70.660 34.480 70.950 34.520 ;
      LAYER met1 ;
        RECT 81.200 34.660 81.520 34.720 ;
        RECT 85.530 34.660 85.820 34.710 ;
        RECT 81.200 34.520 85.820 34.660 ;
        RECT 81.200 34.460 81.520 34.520 ;
        RECT 85.530 34.480 85.820 34.520 ;
        RECT 86.480 34.660 86.800 34.720 ;
        RECT 93.210 34.660 93.500 34.710 ;
        RECT 86.480 34.520 93.500 34.660 ;
        RECT 94.250 34.660 94.390 34.890 ;
        RECT 94.640 34.890 96.380 35.030 ;
        RECT 94.640 34.830 94.960 34.890 ;
        RECT 96.090 34.850 96.380 34.890 ;
        RECT 97.050 34.850 97.340 35.080 ;
        RECT 98.490 34.660 98.780 34.710 ;
        RECT 94.250 34.520 98.780 34.660 ;
        RECT 86.480 34.460 86.800 34.520 ;
        RECT 93.210 34.480 93.500 34.520 ;
        RECT 98.490 34.480 98.780 34.520 ;
        RECT 98.960 34.660 99.280 34.720 ;
        RECT 99.450 34.660 99.740 34.710 ;
        RECT 100.400 34.660 100.720 34.720 ;
        RECT 98.960 34.520 100.720 34.660 ;
        RECT 98.960 34.460 99.280 34.520 ;
        RECT 99.450 34.480 99.740 34.520 ;
        RECT 100.400 34.460 100.720 34.520 ;
        RECT 63.440 34.290 63.760 34.350 ;
        RECT 42.890 34.150 63.760 34.290 ;
        RECT 11.610 33.920 11.900 33.970 ;
        RECT 25.520 33.920 25.840 33.980 ;
        RECT 11.610 33.780 25.840 33.920 ;
        RECT 11.610 33.740 11.900 33.780 ;
        RECT 25.520 33.720 25.840 33.780 ;
        RECT 9.680 33.550 10.000 33.610 ;
        RECT 14.010 33.550 14.300 33.600 ;
        RECT 15.440 33.550 15.760 33.610 ;
        RECT 9.680 33.410 14.300 33.550 ;
        RECT 15.240 33.410 15.760 33.550 ;
        RECT 9.680 33.350 10.000 33.410 ;
        RECT 14.010 33.370 14.300 33.410 ;
        RECT 15.440 33.350 15.760 33.410 ;
        RECT 20.720 33.550 21.040 33.610 ;
        RECT 26.970 33.550 27.260 33.600 ;
        RECT 20.720 33.410 27.260 33.550 ;
        RECT 27.530 33.550 27.670 34.150 ;
        RECT 31.290 34.110 31.580 34.150 ;
        RECT 35.600 34.090 35.920 34.150 ;
        RECT 63.440 34.090 63.760 34.150 ;
        RECT 63.930 34.290 64.220 34.340 ;
        RECT 64.880 34.290 65.200 34.350 ;
        RECT 63.930 34.150 65.200 34.290 ;
        RECT 63.930 34.110 64.220 34.150 ;
        RECT 64.880 34.090 65.200 34.150 ;
        RECT 105.290 33.920 105.430 35.220 ;
        RECT 106.640 35.200 106.960 35.260 ;
        RECT 117.210 35.030 117.500 35.080 ;
        RECT 118.160 35.030 118.480 35.090 ;
        RECT 117.210 34.890 118.480 35.030 ;
        RECT 122.090 35.030 122.230 35.260 ;
        RECT 123.930 35.220 124.220 35.450 ;
        RECT 124.880 35.400 125.200 35.460 ;
        RECT 124.680 35.260 125.200 35.400 ;
        RECT 125.450 35.400 125.590 35.630 ;
        RECT 126.320 35.570 126.640 35.630 ;
        RECT 129.680 35.770 130.000 35.830 ;
        RECT 135.930 35.770 136.220 35.820 ;
        RECT 136.400 35.770 136.720 35.830 ;
        RECT 129.680 35.630 136.720 35.770 ;
        RECT 129.680 35.570 130.000 35.630 ;
        RECT 135.930 35.590 136.220 35.630 ;
        RECT 136.400 35.570 136.720 35.630 ;
        RECT 139.290 35.400 139.580 35.450 ;
        RECT 125.450 35.260 139.580 35.400 ;
        RECT 124.880 35.200 125.200 35.260 ;
        RECT 139.290 35.220 139.580 35.260 ;
        RECT 135.450 35.030 135.740 35.080 ;
        RECT 136.880 35.030 137.200 35.090 ;
        RECT 122.090 34.890 128.950 35.030 ;
        RECT 117.210 34.850 117.500 34.890 ;
        RECT 118.160 34.830 118.480 34.890 ;
        RECT 110.000 34.660 110.320 34.720 ;
        RECT 110.960 34.660 111.280 34.720 ;
        RECT 109.800 34.520 110.320 34.660 ;
        RECT 110.760 34.520 111.280 34.660 ;
        RECT 110.000 34.460 110.320 34.520 ;
        RECT 110.960 34.460 111.280 34.520 ;
        RECT 120.090 34.660 120.380 34.710 ;
        RECT 127.760 34.660 128.080 34.720 ;
        RECT 128.810 34.710 128.950 34.890 ;
        RECT 129.290 34.890 130.870 35.030 ;
        RECT 120.090 34.520 128.080 34.660 ;
        RECT 120.090 34.480 120.380 34.520 ;
        RECT 127.760 34.460 128.080 34.520 ;
        RECT 128.730 34.480 129.020 34.710 ;
        RECT 106.160 34.290 106.480 34.350 ;
        RECT 129.290 34.290 129.430 34.890 ;
        RECT 130.170 34.480 130.460 34.710 ;
        RECT 130.730 34.660 130.870 34.890 ;
        RECT 135.450 34.890 137.200 35.030 ;
        RECT 135.450 34.850 135.740 34.890 ;
        RECT 136.880 34.830 137.200 34.890 ;
        RECT 138.330 34.850 138.620 35.080 ;
        RECT 138.410 34.660 138.550 34.850 ;
        RECT 130.730 34.520 138.550 34.660 ;
        RECT 106.160 34.150 129.430 34.290 ;
        RECT 106.160 34.090 106.480 34.150 ;
        RECT 115.770 33.920 116.060 33.970 ;
        RECT 118.160 33.920 118.480 33.980 ;
        RECT 105.290 33.780 118.480 33.920 ;
        RECT 115.770 33.740 116.060 33.780 ;
        RECT 118.160 33.720 118.480 33.780 ;
        RECT 120.560 33.920 120.880 33.980 ;
        RECT 130.250 33.920 130.390 34.480 ;
        RECT 120.560 33.780 130.390 33.920 ;
        RECT 120.560 33.720 120.880 33.780 ;
        RECT 35.600 33.550 35.920 33.610 ;
        RECT 27.530 33.410 35.920 33.550 ;
        RECT 20.720 33.350 21.040 33.410 ;
        RECT 26.970 33.370 27.260 33.410 ;
        RECT 35.600 33.350 35.920 33.410 ;
        RECT 57.200 33.550 57.520 33.610 ;
        RECT 75.930 33.550 76.220 33.600 ;
        RECT 57.200 33.410 76.220 33.550 ;
        RECT 57.200 33.350 57.520 33.410 ;
        RECT 75.930 33.370 76.220 33.410 ;
        RECT 79.290 33.550 79.580 33.600 ;
        RECT 86.480 33.550 86.800 33.610 ;
        RECT 79.290 33.410 86.800 33.550 ;
        RECT 79.290 33.370 79.580 33.410 ;
        RECT 86.480 33.350 86.800 33.410 ;
        RECT 103.760 33.550 104.080 33.610 ;
        RECT 106.640 33.550 106.960 33.610 ;
        RECT 103.760 33.410 106.960 33.550 ;
        RECT 103.760 33.350 104.080 33.410 ;
        RECT 106.640 33.350 106.960 33.410 ;
        RECT 107.610 33.550 107.900 33.600 ;
        RECT 110.960 33.550 111.280 33.610 ;
        RECT 111.920 33.550 112.240 33.610 ;
        RECT 107.610 33.410 111.280 33.550 ;
        RECT 111.720 33.410 112.240 33.550 ;
        RECT 107.610 33.370 107.900 33.410 ;
        RECT 110.960 33.350 111.280 33.410 ;
        RECT 111.920 33.350 112.240 33.410 ;
        RECT 122.480 33.550 122.800 33.610 ;
        RECT 123.930 33.550 124.220 33.600 ;
        RECT 130.650 33.550 130.940 33.600 ;
        RECT 122.480 33.410 130.940 33.550 ;
        RECT 122.480 33.350 122.800 33.410 ;
        RECT 123.930 33.370 124.220 33.410 ;
        RECT 130.650 33.370 130.940 33.410 ;
        RECT 29.360 31.700 29.680 31.760 ;
        RECT 29.850 31.700 30.140 31.750 ;
        RECT 29.360 31.560 30.140 31.700 ;
        RECT 29.360 31.500 29.680 31.560 ;
        RECT 29.850 31.520 30.140 31.560 ;
        RECT 31.760 31.700 32.080 31.760 ;
        RECT 35.610 31.700 35.900 31.750 ;
        RECT 31.760 31.560 35.900 31.700 ;
        RECT 31.760 31.500 32.080 31.560 ;
        RECT 35.610 31.520 35.900 31.560 ;
        RECT 42.320 31.700 42.640 31.760 ;
        RECT 79.760 31.700 80.080 31.760 ;
        RECT 42.320 31.560 80.080 31.700 ;
        RECT 42.320 31.500 42.640 31.560 ;
        RECT 79.760 31.500 80.080 31.560 ;
        RECT 95.120 31.700 95.440 31.760 ;
        RECT 95.120 31.560 114.550 31.700 ;
        RECT 95.120 31.500 95.440 31.560 ;
        RECT 22.160 31.330 22.480 31.390 ;
        RECT 54.320 31.330 54.640 31.390 ;
        RECT 22.160 31.190 54.640 31.330 ;
        RECT 22.160 31.130 22.480 31.190 ;
        RECT 54.320 31.130 54.640 31.190 ;
        RECT 59.600 31.330 59.920 31.390 ;
        RECT 59.600 31.190 77.590 31.330 ;
        RECT 59.600 31.130 59.920 31.190 ;
        RECT 9.680 30.960 10.000 31.020 ;
        RECT 9.480 30.820 10.000 30.960 ;
        RECT 9.680 30.760 10.000 30.820 ;
        RECT 25.520 30.960 25.840 31.020 ;
        RECT 37.520 30.960 37.840 31.020 ;
        RECT 51.440 30.960 51.760 31.020 ;
        RECT 25.520 30.820 35.830 30.960 ;
        RECT 25.520 30.760 25.840 30.820 ;
      LAYER met1 ;
        RECT 8.740 30.600 9.030 30.640 ;
        RECT 11.140 30.600 11.430 30.640 ;
        RECT 16.420 30.600 16.710 30.640 ;
        RECT 8.740 30.460 16.710 30.600 ;
      LAYER met1 ;
        RECT 32.720 30.590 33.040 30.650 ;
        RECT 35.120 30.590 35.440 30.650 ;
      LAYER met1 ;
        RECT 8.740 30.410 9.030 30.460 ;
        RECT 11.140 30.410 11.430 30.460 ;
        RECT 16.420 30.410 16.710 30.460 ;
      LAYER met1 ;
        RECT 28.970 30.450 33.040 30.590 ;
        RECT 34.920 30.450 35.440 30.590 ;
        RECT 35.690 30.590 35.830 30.820 ;
        RECT 37.520 30.820 48.790 30.960 ;
        RECT 37.520 30.760 37.840 30.820 ;
        RECT 35.690 30.450 39.190 30.590 ;
        RECT 10.170 30.220 10.460 30.270 ;
        RECT 20.720 30.220 21.040 30.280 ;
        RECT 10.170 30.080 21.040 30.220 ;
        RECT 10.170 30.040 10.460 30.080 ;
        RECT 20.720 30.020 21.040 30.080 ;
        RECT 21.690 30.220 21.980 30.270 ;
        RECT 24.090 30.220 24.380 30.270 ;
        RECT 21.690 30.080 24.380 30.220 ;
        RECT 21.690 30.040 21.980 30.080 ;
        RECT 24.090 30.040 24.380 30.080 ;
        RECT 26.960 30.220 27.280 30.280 ;
        RECT 28.970 30.270 29.110 30.450 ;
        RECT 32.720 30.390 33.040 30.450 ;
        RECT 35.120 30.390 35.440 30.450 ;
        RECT 27.450 30.220 27.740 30.270 ;
        RECT 26.960 30.080 27.740 30.220 ;
        RECT 26.960 30.020 27.280 30.080 ;
        RECT 27.450 30.040 27.740 30.080 ;
        RECT 28.890 30.040 29.180 30.270 ;
        RECT 29.360 30.220 29.680 30.280 ;
        RECT 30.330 30.220 30.620 30.270 ;
        RECT 33.680 30.220 34.000 30.280 ;
        RECT 29.360 30.080 30.620 30.220 ;
        RECT 33.480 30.080 34.000 30.220 ;
        RECT 28.970 29.850 29.110 30.040 ;
        RECT 29.360 30.020 29.680 30.080 ;
        RECT 30.330 30.040 30.620 30.080 ;
        RECT 33.680 30.020 34.000 30.080 ;
        RECT 34.170 30.220 34.460 30.270 ;
        RECT 36.080 30.220 36.400 30.280 ;
        RECT 39.050 30.270 39.190 30.450 ;
        RECT 41.370 30.410 41.660 30.640 ;
        RECT 42.320 30.590 42.640 30.650 ;
        RECT 48.650 30.640 48.790 30.820 ;
        RECT 51.440 30.820 73.750 30.960 ;
        RECT 51.440 30.760 51.760 30.820 ;
        RECT 42.120 30.450 42.640 30.590 ;
        RECT 34.170 30.080 36.400 30.220 ;
        RECT 34.170 30.040 34.460 30.080 ;
        RECT 36.080 30.020 36.400 30.080 ;
        RECT 38.970 30.040 39.260 30.270 ;
        RECT 39.930 30.040 40.220 30.270 ;
        RECT 41.450 30.220 41.590 30.410 ;
        RECT 42.320 30.390 42.640 30.450 ;
        RECT 48.570 30.590 48.860 30.640 ;
        RECT 55.280 30.590 55.600 30.650 ;
        RECT 48.570 30.450 55.600 30.590 ;
        RECT 48.570 30.410 48.860 30.450 ;
        RECT 55.280 30.390 55.600 30.450 ;
        RECT 59.120 30.590 59.440 30.650 ;
        RECT 63.930 30.590 64.220 30.640 ;
        RECT 70.650 30.590 70.940 30.640 ;
        RECT 59.120 30.450 64.220 30.590 ;
        RECT 59.120 30.390 59.440 30.450 ;
        RECT 63.930 30.410 64.220 30.450 ;
        RECT 64.490 30.450 70.940 30.590 ;
        RECT 51.450 30.220 51.740 30.270 ;
        RECT 41.450 30.080 51.740 30.220 ;
        RECT 51.450 30.040 51.740 30.080 ;
        RECT 60.560 30.220 60.880 30.280 ;
        RECT 64.490 30.220 64.630 30.450 ;
        RECT 70.650 30.410 70.940 30.450 ;
        RECT 60.560 30.080 64.630 30.220 ;
        RECT 65.360 30.220 65.680 30.280 ;
        RECT 73.610 30.270 73.750 30.820 ;
        RECT 77.450 30.640 77.590 31.190 ;
        RECT 77.370 30.410 77.660 30.640 ;
        RECT 66.810 30.220 67.100 30.270 ;
        RECT 65.360 30.080 67.100 30.220 ;
        RECT 21.770 29.710 29.110 29.850 ;
        RECT 34.640 29.850 34.960 29.910 ;
        RECT 40.010 29.850 40.150 30.040 ;
        RECT 60.560 30.020 60.880 30.080 ;
        RECT 65.360 30.020 65.680 30.080 ;
        RECT 66.810 30.040 67.100 30.080 ;
        RECT 73.530 30.040 73.820 30.270 ;
        RECT 79.850 30.220 79.990 31.500 ;
        RECT 98.000 31.330 98.320 31.390 ;
        RECT 105.680 31.330 106.000 31.390 ;
        RECT 87.050 31.190 106.000 31.330 ;
        RECT 82.640 30.590 82.960 30.650 ;
        RECT 83.600 30.590 83.920 30.650 ;
        RECT 82.440 30.450 82.960 30.590 ;
        RECT 83.400 30.450 83.920 30.590 ;
        RECT 82.640 30.390 82.960 30.450 ;
        RECT 83.600 30.390 83.920 30.450 ;
        RECT 80.250 30.220 80.540 30.270 ;
        RECT 79.850 30.080 80.540 30.220 ;
        RECT 80.250 30.040 80.540 30.080 ;
        RECT 80.720 30.220 81.040 30.280 ;
        RECT 87.050 30.270 87.190 31.190 ;
        RECT 98.000 31.130 98.320 31.190 ;
        RECT 105.680 31.130 106.000 31.190 ;
        RECT 97.520 30.960 97.840 31.020 ;
        RECT 101.840 30.960 102.160 31.020 ;
        RECT 89.450 30.820 97.840 30.960 ;
        RECT 101.640 30.820 102.160 30.960 ;
        RECT 89.450 30.640 89.590 30.820 ;
        RECT 97.520 30.760 97.840 30.820 ;
        RECT 101.840 30.760 102.160 30.820 ;
        RECT 110.960 30.960 111.280 31.020 ;
        RECT 110.960 30.820 113.590 30.960 ;
        RECT 110.960 30.760 111.280 30.820 ;
        RECT 88.410 30.410 88.700 30.640 ;
        RECT 89.370 30.410 89.660 30.640 ;
        RECT 94.160 30.590 94.480 30.650 ;
        RECT 93.960 30.450 94.480 30.590 ;
        RECT 81.210 30.220 81.500 30.270 ;
        RECT 80.720 30.080 81.500 30.220 ;
        RECT 80.720 30.020 81.040 30.080 ;
        RECT 81.210 30.040 81.500 30.080 ;
        RECT 86.010 30.040 86.300 30.270 ;
        RECT 86.970 30.040 87.260 30.270 ;
        RECT 88.490 30.220 88.630 30.410 ;
        RECT 94.160 30.390 94.480 30.450 ;
        RECT 94.650 30.590 94.940 30.640 ;
        RECT 100.880 30.590 101.200 30.650 ;
        RECT 94.650 30.450 101.200 30.590 ;
        RECT 94.650 30.410 94.940 30.450 ;
        RECT 100.880 30.390 101.200 30.450 ;
        RECT 107.130 30.410 107.420 30.640 ;
        RECT 108.080 30.590 108.400 30.650 ;
        RECT 113.450 30.640 113.590 30.820 ;
        RECT 107.880 30.450 108.400 30.590 ;
        RECT 91.770 30.220 92.060 30.270 ;
        RECT 95.120 30.220 95.440 30.280 ;
        RECT 88.490 30.080 92.060 30.220 ;
        RECT 94.920 30.080 95.440 30.220 ;
        RECT 91.770 30.040 92.060 30.080 ;
        RECT 34.640 29.710 40.150 29.850 ;
        RECT 47.130 29.850 47.420 29.900 ;
        RECT 48.080 29.850 48.400 29.910 ;
        RECT 62.480 29.850 62.800 29.910 ;
        RECT 47.130 29.710 48.400 29.850 ;
        RECT 62.280 29.710 62.800 29.850 ;
        RECT 86.090 29.850 86.230 30.040 ;
        RECT 95.120 30.020 95.440 30.080 ;
        RECT 96.090 30.220 96.380 30.270 ;
        RECT 98.960 30.220 99.280 30.280 ;
        RECT 96.090 30.080 99.280 30.220 ;
        RECT 96.090 30.040 96.380 30.080 ;
        RECT 98.960 30.020 99.280 30.080 ;
        RECT 104.730 30.040 105.020 30.270 ;
        RECT 105.680 30.220 106.000 30.280 ;
        RECT 105.480 30.080 106.000 30.220 ;
        RECT 107.210 30.220 107.350 30.410 ;
        RECT 108.080 30.390 108.400 30.450 ;
        RECT 112.890 30.410 113.180 30.640 ;
        RECT 113.370 30.410 113.660 30.640 ;
        RECT 110.490 30.220 110.780 30.270 ;
        RECT 107.210 30.080 110.780 30.220 ;
        RECT 93.680 29.850 94.000 29.910 ;
        RECT 99.440 29.850 99.760 29.910 ;
        RECT 86.090 29.710 94.000 29.850 ;
        RECT 99.240 29.710 99.760 29.850 ;
        RECT 21.770 29.540 21.910 29.710 ;
        RECT 34.640 29.650 34.960 29.710 ;
        RECT 47.130 29.670 47.420 29.710 ;
        RECT 48.080 29.650 48.400 29.710 ;
        RECT 62.480 29.650 62.800 29.710 ;
        RECT 93.680 29.650 94.000 29.710 ;
        RECT 99.440 29.650 99.760 29.710 ;
        RECT 100.410 29.850 100.700 29.900 ;
        RECT 103.280 29.850 103.600 29.910 ;
        RECT 100.410 29.710 103.600 29.850 ;
        RECT 104.810 29.850 104.950 30.040 ;
        RECT 105.680 30.020 106.000 30.080 ;
        RECT 110.490 30.040 110.780 30.080 ;
        RECT 111.440 29.850 111.760 29.910 ;
        RECT 104.810 29.710 111.760 29.850 ;
        RECT 100.410 29.670 100.700 29.710 ;
        RECT 103.280 29.650 103.600 29.710 ;
        RECT 111.440 29.650 111.760 29.710 ;
        RECT 21.680 29.280 22.000 29.540 ;
        RECT 25.050 29.480 25.340 29.530 ;
        RECT 29.840 29.480 30.160 29.540 ;
        RECT 33.680 29.480 34.000 29.540 ;
        RECT 25.050 29.340 34.000 29.480 ;
        RECT 25.050 29.300 25.340 29.340 ;
        RECT 29.840 29.280 30.160 29.340 ;
        RECT 33.680 29.280 34.000 29.340 ;
        RECT 39.930 29.480 40.220 29.530 ;
        RECT 47.600 29.480 47.920 29.540 ;
        RECT 39.930 29.340 47.920 29.480 ;
        RECT 39.930 29.300 40.220 29.340 ;
        RECT 47.600 29.280 47.920 29.340 ;
        RECT 72.080 29.480 72.400 29.540 ;
        RECT 81.210 29.480 81.500 29.530 ;
        RECT 72.080 29.340 81.500 29.480 ;
        RECT 72.080 29.280 72.400 29.340 ;
        RECT 81.210 29.300 81.500 29.340 ;
        RECT 86.000 29.480 86.320 29.540 ;
        RECT 86.970 29.480 87.260 29.530 ;
        RECT 105.680 29.480 106.000 29.540 ;
        RECT 86.000 29.340 87.260 29.480 ;
        RECT 105.480 29.340 106.000 29.480 ;
        RECT 112.970 29.480 113.110 30.410 ;
        RECT 114.410 30.270 114.550 31.560 ;
        RECT 121.040 31.330 121.360 31.390 ;
        RECT 137.840 31.330 138.160 31.390 ;
        RECT 121.040 31.190 138.160 31.330 ;
        RECT 121.040 31.130 121.360 31.190 ;
        RECT 137.840 31.130 138.160 31.190 ;
        RECT 119.690 30.820 127.990 30.960 ;
        RECT 114.330 30.040 114.620 30.270 ;
        RECT 119.690 30.220 119.830 30.820 ;
        RECT 122.250 30.590 122.540 30.640 ;
        RECT 122.960 30.590 123.280 30.650 ;
        RECT 121.610 30.450 122.540 30.590 ;
        RECT 122.760 30.450 123.280 30.590 ;
        RECT 120.090 30.220 120.380 30.270 ;
        RECT 121.040 30.220 121.360 30.280 ;
        RECT 116.330 30.080 120.380 30.220 ;
        RECT 120.840 30.080 121.360 30.220 ;
        RECT 121.610 30.220 121.750 30.450 ;
        RECT 122.250 30.410 122.540 30.450 ;
        RECT 122.960 30.390 123.280 30.450 ;
        RECT 127.850 30.590 127.990 30.820 ;
        RECT 133.530 30.590 133.820 30.640 ;
        RECT 127.850 30.450 133.820 30.590 ;
        RECT 123.440 30.220 123.760 30.280 ;
        RECT 127.850 30.270 127.990 30.450 ;
        RECT 133.530 30.410 133.820 30.450 ;
        RECT 121.610 30.080 123.760 30.220 ;
        RECT 113.850 29.850 114.140 29.900 ;
        RECT 115.280 29.850 115.600 29.910 ;
        RECT 116.330 29.850 116.470 30.080 ;
        RECT 120.090 30.040 120.380 30.080 ;
        RECT 121.040 30.020 121.360 30.080 ;
        RECT 123.440 30.020 123.760 30.080 ;
        RECT 125.850 30.040 126.140 30.270 ;
        RECT 127.770 30.040 128.060 30.270 ;
        RECT 133.050 30.220 133.340 30.270 ;
        RECT 136.880 30.220 137.200 30.280 ;
        RECT 133.050 30.080 137.200 30.220 ;
        RECT 133.050 30.040 133.340 30.080 ;
        RECT 113.850 29.710 116.470 29.850 ;
        RECT 116.720 29.850 117.040 29.910 ;
        RECT 125.930 29.850 126.070 30.040 ;
        RECT 136.880 30.020 137.200 30.080 ;
        RECT 127.280 29.850 127.600 29.910 ;
        RECT 116.720 29.710 126.070 29.850 ;
        RECT 127.080 29.710 127.600 29.850 ;
        RECT 113.850 29.670 114.140 29.710 ;
        RECT 115.280 29.650 115.600 29.710 ;
        RECT 116.720 29.650 117.040 29.710 ;
        RECT 127.280 29.650 127.600 29.710 ;
        RECT 117.680 29.480 118.000 29.540 ;
        RECT 112.970 29.340 118.000 29.480 ;
        RECT 86.000 29.280 86.320 29.340 ;
        RECT 86.970 29.300 87.260 29.340 ;
        RECT 105.680 29.280 106.000 29.340 ;
        RECT 117.680 29.280 118.000 29.340 ;
        RECT 121.050 29.480 121.340 29.530 ;
        RECT 125.360 29.480 125.680 29.540 ;
        RECT 121.050 29.340 125.680 29.480 ;
        RECT 121.050 29.300 121.340 29.340 ;
        RECT 125.360 29.280 125.680 29.340 ;
        RECT 5.760 28.750 142.080 29.120 ;
        RECT 15.930 27.630 16.220 27.680 ;
        RECT 21.680 27.630 22.000 27.690 ;
        RECT 33.680 27.630 34.000 27.690 ;
        RECT 15.930 27.490 22.000 27.630 ;
        RECT 15.930 27.450 16.220 27.490 ;
        RECT 21.680 27.430 22.000 27.490 ;
        RECT 22.250 27.490 31.990 27.630 ;
        RECT 33.480 27.490 34.000 27.630 ;
        RECT 19.280 27.260 19.600 27.320 ;
        RECT 22.250 27.260 22.390 27.490 ;
        RECT 19.280 27.120 22.390 27.260 ;
        RECT 26.000 27.260 26.320 27.320 ;
        RECT 26.000 27.120 31.510 27.260 ;
        RECT 19.280 27.060 19.600 27.120 ;
        RECT 26.000 27.060 26.320 27.120 ;
        RECT 15.450 26.890 15.740 26.940 ;
        RECT 26.480 26.890 26.800 26.950 ;
        RECT 31.370 26.940 31.510 27.120 ;
        RECT 28.890 26.890 29.180 26.940 ;
        RECT 15.450 26.750 26.230 26.890 ;
        RECT 15.450 26.710 15.740 26.750 ;
        RECT 19.290 26.340 19.580 26.570 ;
        RECT 19.760 26.520 20.080 26.580 ;
        RECT 26.090 26.520 26.230 26.750 ;
        RECT 26.480 26.750 29.180 26.890 ;
        RECT 26.480 26.690 26.800 26.750 ;
        RECT 28.890 26.710 29.180 26.750 ;
        RECT 31.290 26.710 31.580 26.940 ;
        RECT 31.850 26.890 31.990 27.490 ;
        RECT 33.680 27.430 34.000 27.490 ;
        RECT 41.850 27.630 42.140 27.680 ;
        RECT 102.330 27.630 102.620 27.680 ;
        RECT 103.280 27.630 103.600 27.690 ;
        RECT 106.640 27.630 106.960 27.690 ;
        RECT 41.850 27.490 46.870 27.630 ;
        RECT 41.850 27.450 42.140 27.490 ;
        RECT 32.720 27.260 33.040 27.320 ;
        RECT 33.210 27.260 33.500 27.310 ;
        RECT 32.720 27.120 33.500 27.260 ;
        RECT 32.720 27.060 33.040 27.120 ;
        RECT 33.210 27.080 33.500 27.120 ;
        RECT 43.760 27.260 44.080 27.320 ;
        RECT 46.730 27.310 46.870 27.490 ;
        RECT 54.890 27.490 66.550 27.630 ;
        RECT 54.890 27.310 55.030 27.490 ;
        RECT 45.210 27.260 45.500 27.310 ;
        RECT 43.760 27.120 45.500 27.260 ;
        RECT 43.760 27.060 44.080 27.120 ;
        RECT 45.210 27.080 45.500 27.120 ;
        RECT 46.650 27.080 46.940 27.310 ;
        RECT 54.810 27.080 55.100 27.310 ;
        RECT 38.010 26.890 38.300 26.940 ;
        RECT 31.850 26.750 38.300 26.890 ;
        RECT 38.010 26.710 38.300 26.750 ;
        RECT 38.480 26.890 38.800 26.950 ;
        RECT 48.090 26.890 48.380 26.940 ;
        RECT 38.480 26.750 48.380 26.890 ;
        RECT 38.480 26.690 38.800 26.750 ;
        RECT 48.090 26.710 48.380 26.750 ;
        RECT 60.570 26.890 60.860 26.940 ;
        RECT 60.570 26.750 61.750 26.890 ;
        RECT 60.570 26.710 60.860 26.750 ;
        RECT 26.970 26.520 27.260 26.570 ;
        RECT 19.760 26.380 20.280 26.520 ;
        RECT 26.090 26.380 27.260 26.520 ;
        RECT 19.370 26.150 19.510 26.340 ;
        RECT 19.760 26.320 20.080 26.380 ;
        RECT 26.970 26.340 27.260 26.380 ;
        RECT 27.440 26.520 27.760 26.580 ;
        RECT 28.410 26.520 28.700 26.570 ;
        RECT 27.440 26.380 28.700 26.520 ;
        RECT 22.160 26.150 22.480 26.210 ;
        RECT 24.080 26.150 24.400 26.210 ;
        RECT 19.370 26.010 22.480 26.150 ;
        RECT 23.880 26.010 24.400 26.150 ;
        RECT 27.050 26.150 27.190 26.340 ;
        RECT 27.440 26.320 27.760 26.380 ;
        RECT 28.410 26.340 28.700 26.380 ;
        RECT 36.080 26.520 36.400 26.580 ;
        RECT 39.440 26.520 39.760 26.580 ;
        RECT 40.400 26.520 40.720 26.580 ;
        RECT 56.240 26.520 56.560 26.580 ;
        RECT 36.080 26.380 39.760 26.520 ;
        RECT 40.200 26.380 56.560 26.520 ;
        RECT 36.080 26.320 36.400 26.380 ;
        RECT 39.440 26.320 39.760 26.380 ;
        RECT 40.400 26.320 40.720 26.380 ;
        RECT 56.240 26.320 56.560 26.380 ;
        RECT 56.730 26.520 57.020 26.570 ;
        RECT 58.640 26.520 58.960 26.580 ;
        RECT 56.730 26.380 58.960 26.520 ;
        RECT 56.730 26.340 57.020 26.380 ;
        RECT 58.640 26.320 58.960 26.380 ;
        RECT 35.120 26.150 35.440 26.210 ;
        RECT 27.050 26.010 35.440 26.150 ;
        RECT 22.160 25.950 22.480 26.010 ;
        RECT 24.080 25.950 24.400 26.010 ;
        RECT 35.120 25.950 35.440 26.010 ;
        RECT 35.600 26.150 35.920 26.210 ;
        RECT 41.370 26.150 41.660 26.200 ;
        RECT 35.600 26.010 41.660 26.150 ;
        RECT 61.610 26.150 61.750 26.750 ;
        RECT 63.450 26.520 63.740 26.570 ;
        RECT 65.360 26.520 65.680 26.580 ;
        RECT 63.450 26.380 65.680 26.520 ;
        RECT 66.410 26.520 66.550 27.490 ;
        RECT 102.330 27.490 103.600 27.630 ;
        RECT 106.440 27.490 106.960 27.630 ;
        RECT 102.330 27.450 102.620 27.490 ;
        RECT 103.280 27.430 103.600 27.490 ;
        RECT 106.640 27.430 106.960 27.490 ;
        RECT 111.440 27.630 111.760 27.690 ;
        RECT 124.880 27.630 125.200 27.690 ;
        RECT 126.810 27.630 127.100 27.680 ;
        RECT 111.440 27.490 113.110 27.630 ;
        RECT 111.440 27.430 111.760 27.490 ;
        RECT 68.720 27.260 69.040 27.320 ;
        RECT 96.080 27.260 96.400 27.320 ;
        RECT 68.520 27.120 69.040 27.260 ;
        RECT 95.880 27.120 96.400 27.260 ;
        RECT 68.720 27.060 69.040 27.120 ;
        RECT 96.080 27.060 96.400 27.120 ;
        RECT 111.920 27.260 112.240 27.320 ;
        RECT 112.410 27.260 112.700 27.310 ;
        RECT 111.920 27.120 112.700 27.260 ;
        RECT 111.920 27.060 112.240 27.120 ;
        RECT 112.410 27.080 112.700 27.120 ;
        RECT 112.970 27.260 113.110 27.490 ;
        RECT 117.290 27.490 127.100 27.630 ;
        RECT 117.290 27.260 117.430 27.490 ;
        RECT 124.880 27.430 125.200 27.490 ;
        RECT 126.810 27.450 127.100 27.490 ;
        RECT 112.970 27.120 117.430 27.260 ;
        RECT 68.240 26.890 68.560 26.950 ;
        RECT 73.050 26.890 73.340 26.940 ;
        RECT 68.240 26.750 73.340 26.890 ;
        RECT 68.240 26.690 68.560 26.750 ;
        RECT 73.050 26.710 73.340 26.750 ;
        RECT 83.610 26.890 83.900 26.940 ;
        RECT 86.480 26.890 86.800 26.950 ;
        RECT 83.610 26.750 90.550 26.890 ;
        RECT 83.610 26.710 83.900 26.750 ;
        RECT 86.480 26.690 86.800 26.750 ;
        RECT 70.170 26.520 70.460 26.570 ;
        RECT 76.880 26.520 77.200 26.580 ;
        RECT 90.410 26.570 90.550 26.750 ;
        RECT 95.130 26.710 95.420 26.940 ;
        RECT 96.570 26.890 96.860 26.940 ;
        RECT 97.520 26.890 97.840 26.950 ;
        RECT 98.970 26.890 99.260 26.940 ;
        RECT 103.760 26.890 104.080 26.950 ;
        RECT 96.570 26.750 99.260 26.890 ;
        RECT 103.560 26.750 104.080 26.890 ;
        RECT 96.570 26.710 96.860 26.750 ;
        RECT 66.410 26.380 70.460 26.520 ;
        RECT 76.680 26.380 77.200 26.520 ;
        RECT 63.450 26.340 63.740 26.380 ;
        RECT 65.360 26.320 65.680 26.380 ;
        RECT 70.170 26.340 70.460 26.380 ;
        RECT 76.880 26.320 77.200 26.380 ;
        RECT 89.850 26.340 90.140 26.570 ;
        RECT 90.330 26.340 90.620 26.570 ;
        RECT 94.640 26.520 94.960 26.580 ;
        RECT 95.210 26.520 95.350 26.710 ;
        RECT 97.520 26.690 97.840 26.750 ;
        RECT 98.970 26.710 99.260 26.750 ;
        RECT 103.760 26.690 104.080 26.750 ;
        RECT 108.090 26.890 108.380 26.940 ;
        RECT 108.560 26.890 108.880 26.950 ;
        RECT 112.970 26.940 113.110 27.120 ;
        RECT 108.090 26.750 108.880 26.890 ;
        RECT 108.090 26.710 108.380 26.750 ;
        RECT 108.560 26.690 108.880 26.750 ;
        RECT 111.450 26.710 111.740 26.940 ;
        RECT 112.890 26.710 113.180 26.940 ;
        RECT 99.440 26.520 99.760 26.580 ;
        RECT 94.640 26.380 99.760 26.520 ;
        RECT 111.530 26.520 111.670 26.710 ;
        RECT 115.280 26.520 115.600 26.580 ;
        RECT 116.720 26.520 117.040 26.580 ;
        RECT 117.290 26.570 117.430 27.120 ;
        RECT 117.690 27.260 117.980 27.310 ;
        RECT 118.160 27.260 118.480 27.320 ;
        RECT 127.280 27.260 127.600 27.320 ;
        RECT 117.690 27.120 118.480 27.260 ;
        RECT 117.690 27.080 117.980 27.120 ;
        RECT 118.160 27.060 118.480 27.120 ;
        RECT 121.610 27.120 127.600 27.260 ;
        RECT 121.610 26.940 121.750 27.120 ;
        RECT 127.280 27.060 127.600 27.120 ;
        RECT 121.530 26.710 121.820 26.940 ;
        RECT 122.010 26.890 122.300 26.940 ;
        RECT 122.480 26.890 122.800 26.950 ;
        RECT 123.440 26.890 123.760 26.950 ;
        RECT 122.010 26.750 122.800 26.890 ;
        RECT 123.240 26.750 123.760 26.890 ;
        RECT 122.010 26.710 122.300 26.750 ;
        RECT 122.480 26.690 122.800 26.750 ;
        RECT 123.440 26.690 123.760 26.750 ;
        RECT 125.850 26.710 126.140 26.940 ;
        RECT 130.640 26.890 130.960 26.950 ;
        RECT 130.440 26.750 130.960 26.890 ;
        RECT 111.530 26.380 115.800 26.520 ;
        RECT 116.520 26.380 117.040 26.520 ;
        RECT 82.640 26.150 82.960 26.210 ;
        RECT 61.610 26.010 82.960 26.150 ;
        RECT 89.930 26.150 90.070 26.340 ;
        RECT 94.640 26.320 94.960 26.380 ;
        RECT 99.440 26.320 99.760 26.380 ;
        RECT 115.280 26.320 115.600 26.380 ;
        RECT 116.720 26.320 117.040 26.380 ;
        RECT 117.210 26.340 117.500 26.570 ;
        RECT 118.160 26.520 118.480 26.580 ;
        RECT 125.930 26.520 126.070 26.710 ;
        RECT 130.640 26.690 130.960 26.750 ;
        RECT 118.160 26.380 126.070 26.520 ;
        RECT 118.160 26.320 118.480 26.380 ;
        RECT 93.680 26.150 94.000 26.210 ;
        RECT 99.930 26.150 100.220 26.200 ;
        RECT 89.930 26.010 100.220 26.150 ;
        RECT 35.600 25.950 35.920 26.010 ;
        RECT 41.370 25.970 41.660 26.010 ;
        RECT 82.640 25.950 82.960 26.010 ;
        RECT 93.680 25.950 94.000 26.010 ;
        RECT 99.930 25.970 100.220 26.010 ;
        RECT 19.760 25.780 20.080 25.840 ;
        RECT 22.650 25.780 22.940 25.830 ;
        RECT 64.880 25.780 65.200 25.840 ;
        RECT 19.760 25.640 22.390 25.780 ;
        RECT 19.760 25.580 20.080 25.640 ;
        RECT 20.240 25.410 20.560 25.470 ;
        RECT 20.040 25.270 20.560 25.410 ;
        RECT 22.250 25.410 22.390 25.640 ;
        RECT 22.650 25.640 65.200 25.780 ;
        RECT 22.650 25.600 22.940 25.640 ;
        RECT 64.880 25.580 65.200 25.640 ;
        RECT 90.810 25.780 91.100 25.830 ;
        RECT 110.000 25.780 110.320 25.840 ;
        RECT 122.970 25.780 123.260 25.830 ;
        RECT 90.810 25.640 123.260 25.780 ;
        RECT 90.810 25.600 91.100 25.640 ;
        RECT 110.000 25.580 110.320 25.640 ;
        RECT 122.970 25.600 123.260 25.640 ;
        RECT 34.170 25.410 34.460 25.460 ;
        RECT 34.640 25.410 34.960 25.470 ;
        RECT 22.250 25.270 34.960 25.410 ;
        RECT 20.240 25.210 20.560 25.270 ;
        RECT 34.170 25.230 34.460 25.270 ;
        RECT 34.640 25.210 34.960 25.270 ;
        RECT 38.010 25.410 38.300 25.460 ;
        RECT 45.210 25.410 45.500 25.460 ;
        RECT 38.010 25.270 45.500 25.410 ;
        RECT 38.010 25.230 38.300 25.270 ;
        RECT 45.210 25.230 45.500 25.270 ;
        RECT 82.170 25.410 82.460 25.460 ;
        RECT 86.960 25.410 87.280 25.470 ;
        RECT 129.200 25.410 129.520 25.470 ;
        RECT 82.170 25.270 87.280 25.410 ;
        RECT 129.000 25.270 129.520 25.410 ;
        RECT 82.170 25.230 82.460 25.270 ;
        RECT 86.960 25.210 87.280 25.270 ;
        RECT 129.200 25.210 129.520 25.270 ;
        RECT 20.240 23.560 20.560 23.620 ;
        RECT 67.280 23.560 67.600 23.620 ;
        RECT 78.800 23.560 79.120 23.620 ;
        RECT 82.650 23.560 82.940 23.610 ;
        RECT 86.960 23.560 87.280 23.620 ;
        RECT 20.240 23.420 67.600 23.560 ;
        RECT 78.600 23.420 82.940 23.560 ;
        RECT 86.760 23.420 87.280 23.560 ;
        RECT 20.240 23.360 20.560 23.420 ;
        RECT 67.280 23.360 67.600 23.420 ;
        RECT 78.800 23.360 79.120 23.420 ;
        RECT 82.650 23.380 82.940 23.420 ;
        RECT 86.960 23.360 87.280 23.420 ;
        RECT 92.730 23.560 93.020 23.610 ;
        RECT 94.160 23.560 94.480 23.620 ;
        RECT 92.730 23.420 94.480 23.560 ;
        RECT 92.730 23.380 93.020 23.420 ;
        RECT 94.160 23.360 94.480 23.420 ;
        RECT 117.680 23.560 118.000 23.620 ;
        RECT 119.610 23.560 119.900 23.610 ;
        RECT 136.880 23.560 137.200 23.620 ;
        RECT 117.680 23.420 119.900 23.560 ;
        RECT 136.680 23.420 137.200 23.560 ;
        RECT 117.680 23.360 118.000 23.420 ;
        RECT 119.610 23.380 119.900 23.420 ;
        RECT 136.880 23.360 137.200 23.420 ;
        RECT 35.120 23.190 35.440 23.250 ;
        RECT 40.890 23.190 41.180 23.240 ;
        RECT 35.120 23.050 41.180 23.190 ;
        RECT 35.120 22.990 35.440 23.050 ;
        RECT 40.890 23.010 41.180 23.050 ;
        RECT 42.800 23.190 43.120 23.250 ;
        RECT 59.610 23.190 59.900 23.240 ;
        RECT 42.800 23.050 59.900 23.190 ;
        RECT 42.800 22.990 43.120 23.050 ;
        RECT 59.610 23.010 59.900 23.050 ;
        RECT 64.880 23.190 65.200 23.250 ;
        RECT 66.800 23.190 67.120 23.250 ;
        RECT 81.200 23.190 81.520 23.250 ;
        RECT 64.880 23.050 67.120 23.190 ;
        RECT 81.000 23.050 81.520 23.190 ;
        RECT 64.880 22.990 65.200 23.050 ;
        RECT 66.800 22.990 67.120 23.050 ;
        RECT 81.200 22.990 81.520 23.050 ;
        RECT 87.440 23.190 87.760 23.250 ;
        RECT 103.760 23.190 104.080 23.250 ;
        RECT 130.640 23.190 130.960 23.250 ;
        RECT 87.440 23.050 104.080 23.190 ;
        RECT 87.440 22.990 87.760 23.050 ;
        RECT 103.760 22.990 104.080 23.050 ;
        RECT 110.570 23.050 130.960 23.190 ;
        RECT 52.880 22.820 53.200 22.880 ;
        RECT 67.760 22.820 68.080 22.880 ;
        RECT 97.520 22.820 97.840 22.880 ;
        RECT 52.880 22.680 68.080 22.820 ;
        RECT 52.880 22.620 53.200 22.680 ;
        RECT 67.760 22.620 68.080 22.680 ;
        RECT 91.850 22.680 97.840 22.820 ;
        RECT 91.850 22.500 91.990 22.680 ;
        RECT 97.520 22.620 97.840 22.680 ;
        RECT 98.970 22.820 99.260 22.870 ;
        RECT 108.570 22.820 108.860 22.870 ;
        RECT 98.970 22.680 108.860 22.820 ;
        RECT 98.970 22.640 99.260 22.680 ;
        RECT 108.570 22.640 108.860 22.680 ;
      LAYER met1 ;
        RECT 27.940 22.460 28.230 22.500 ;
        RECT 30.340 22.460 30.630 22.500 ;
        RECT 35.620 22.460 35.910 22.500 ;
        RECT 27.940 22.320 35.910 22.460 ;
        RECT 27.940 22.270 28.230 22.320 ;
        RECT 30.340 22.270 30.630 22.320 ;
        RECT 35.620 22.270 35.910 22.320 ;
        RECT 65.860 22.460 66.150 22.500 ;
        RECT 68.260 22.460 68.550 22.500 ;
        RECT 73.540 22.460 73.830 22.500 ;
        RECT 65.860 22.320 73.830 22.460 ;
        RECT 65.860 22.270 66.150 22.320 ;
        RECT 68.260 22.270 68.550 22.320 ;
        RECT 73.540 22.270 73.830 22.320 ;
      LAYER met1 ;
        RECT 91.770 22.270 92.060 22.500 ;
        RECT 92.250 22.450 92.540 22.500 ;
        RECT 94.640 22.450 94.960 22.510 ;
        RECT 110.570 22.500 110.710 23.050 ;
        RECT 130.640 22.990 130.960 23.050 ;
        RECT 115.280 22.820 115.600 22.880 ;
        RECT 114.410 22.680 115.600 22.820 ;
        RECT 114.410 22.500 114.550 22.680 ;
        RECT 115.280 22.620 115.600 22.680 ;
        RECT 124.890 22.820 125.180 22.870 ;
        RECT 129.200 22.820 129.520 22.880 ;
        RECT 124.890 22.680 129.520 22.820 ;
        RECT 124.890 22.640 125.180 22.680 ;
        RECT 129.200 22.620 129.520 22.680 ;
        RECT 92.250 22.310 94.960 22.450 ;
        RECT 92.250 22.270 92.540 22.310 ;
        RECT 94.640 22.250 94.960 22.310 ;
        RECT 96.570 22.450 96.860 22.500 ;
        RECT 110.490 22.450 110.780 22.500 ;
        RECT 96.570 22.310 110.780 22.450 ;
        RECT 96.570 22.270 96.860 22.310 ;
        RECT 110.490 22.270 110.780 22.310 ;
        RECT 114.330 22.270 114.620 22.500 ;
        RECT 114.810 22.450 115.100 22.500 ;
        RECT 116.720 22.450 117.040 22.510 ;
        RECT 118.160 22.450 118.480 22.510 ;
        RECT 114.810 22.310 117.040 22.450 ;
        RECT 117.960 22.310 118.480 22.450 ;
        RECT 114.810 22.270 115.100 22.310 ;
        RECT 29.360 22.080 29.680 22.140 ;
        RECT 47.600 22.080 47.920 22.140 ;
        RECT 29.160 21.940 29.680 22.080 ;
        RECT 47.400 21.940 47.920 22.080 ;
        RECT 29.360 21.880 29.680 21.940 ;
        RECT 47.600 21.880 47.920 21.940 ;
        RECT 67.290 22.080 67.580 22.130 ;
        RECT 72.080 22.080 72.400 22.140 ;
        RECT 67.290 21.940 72.400 22.080 ;
        RECT 67.290 21.900 67.580 21.940 ;
        RECT 72.080 21.880 72.400 21.940 ;
        RECT 96.080 22.080 96.400 22.140 ;
        RECT 98.970 22.080 99.260 22.130 ;
        RECT 99.450 22.080 99.740 22.130 ;
        RECT 101.360 22.080 101.680 22.140 ;
        RECT 103.760 22.080 104.080 22.140 ;
        RECT 105.690 22.080 105.980 22.130 ;
        RECT 96.080 21.940 99.740 22.080 ;
        RECT 101.160 21.940 101.680 22.080 ;
        RECT 103.560 21.940 104.080 22.080 ;
        RECT 96.080 21.880 96.400 21.940 ;
        RECT 98.970 21.900 99.260 21.940 ;
        RECT 99.450 21.900 99.740 21.940 ;
        RECT 101.360 21.880 101.680 21.940 ;
        RECT 103.760 21.880 104.080 21.940 ;
        RECT 104.330 21.940 105.980 22.080 ;
        RECT 99.920 21.510 100.240 21.770 ;
        RECT 100.880 21.710 101.200 21.770 ;
        RECT 104.330 21.710 104.470 21.940 ;
        RECT 105.690 21.900 105.980 21.940 ;
        RECT 108.570 22.080 108.860 22.130 ;
        RECT 114.890 22.080 115.030 22.270 ;
        RECT 116.720 22.250 117.040 22.310 ;
        RECT 118.160 22.250 118.480 22.310 ;
        RECT 119.130 22.450 119.420 22.500 ;
        RECT 120.560 22.450 120.880 22.510 ;
        RECT 119.130 22.310 120.880 22.450 ;
        RECT 119.130 22.270 119.420 22.310 ;
        RECT 108.570 21.940 115.030 22.080 ;
        RECT 115.290 22.080 115.580 22.130 ;
        RECT 119.210 22.080 119.350 22.270 ;
        RECT 120.560 22.250 120.880 22.310 ;
      LAYER met1 ;
        RECT 123.940 22.460 124.230 22.500 ;
        RECT 126.340 22.460 126.630 22.500 ;
        RECT 131.620 22.460 131.910 22.500 ;
        RECT 123.940 22.320 131.910 22.460 ;
        RECT 123.940 22.270 124.230 22.320 ;
        RECT 126.340 22.270 126.630 22.320 ;
        RECT 131.620 22.270 131.910 22.320 ;
      LAYER met1 ;
        RECT 125.360 22.080 125.680 22.140 ;
        RECT 115.290 21.940 119.350 22.080 ;
        RECT 125.160 21.940 125.680 22.080 ;
        RECT 108.570 21.900 108.860 21.940 ;
        RECT 115.290 21.900 115.580 21.940 ;
        RECT 125.360 21.880 125.680 21.940 ;
        RECT 105.200 21.710 105.520 21.770 ;
        RECT 100.680 21.570 101.200 21.710 ;
        RECT 100.880 21.510 101.200 21.570 ;
        RECT 101.450 21.570 104.470 21.710 ;
        RECT 105.000 21.570 105.520 21.710 ;
        RECT 28.890 21.340 29.180 21.390 ;
        RECT 33.200 21.340 33.520 21.400 ;
        RECT 53.360 21.340 53.680 21.400 ;
        RECT 66.800 21.340 67.120 21.400 ;
        RECT 28.890 21.200 33.520 21.340 ;
        RECT 53.160 21.200 53.680 21.340 ;
        RECT 66.600 21.200 67.120 21.340 ;
        RECT 28.890 21.160 29.180 21.200 ;
        RECT 33.200 21.140 33.520 21.200 ;
        RECT 53.360 21.140 53.680 21.200 ;
        RECT 66.800 21.140 67.120 21.200 ;
        RECT 69.680 21.340 70.000 21.400 ;
        RECT 83.600 21.340 83.920 21.400 ;
        RECT 85.530 21.340 85.820 21.390 ;
        RECT 69.680 21.200 85.820 21.340 ;
        RECT 69.680 21.140 70.000 21.200 ;
        RECT 83.600 21.140 83.920 21.200 ;
        RECT 85.530 21.160 85.820 21.200 ;
        RECT 94.160 21.340 94.480 21.400 ;
        RECT 95.130 21.340 95.420 21.390 ;
        RECT 94.160 21.200 95.420 21.340 ;
        RECT 100.010 21.340 100.150 21.510 ;
        RECT 101.450 21.340 101.590 21.570 ;
        RECT 105.200 21.510 105.520 21.570 ;
        RECT 109.040 21.340 109.360 21.400 ;
        RECT 100.010 21.200 101.590 21.340 ;
        RECT 108.840 21.200 109.360 21.340 ;
        RECT 94.160 21.140 94.480 21.200 ;
        RECT 95.130 21.160 95.420 21.200 ;
        RECT 109.040 21.140 109.360 21.200 ;
        RECT 5.760 20.610 142.080 20.980 ;
        RECT 24.570 19.490 24.860 19.540 ;
        RECT 53.360 19.490 53.680 19.550 ;
        RECT 24.570 19.350 53.680 19.490 ;
        RECT 24.570 19.310 24.860 19.350 ;
        RECT 53.360 19.290 53.680 19.350 ;
        RECT 56.240 19.490 56.560 19.550 ;
        RECT 57.210 19.490 57.500 19.540 ;
        RECT 65.840 19.490 66.160 19.550 ;
        RECT 56.240 19.350 66.160 19.490 ;
        RECT 56.240 19.290 56.560 19.350 ;
        RECT 57.210 19.310 57.500 19.350 ;
        RECT 65.840 19.290 66.160 19.350 ;
        RECT 66.320 19.490 66.640 19.550 ;
        RECT 67.290 19.490 67.580 19.540 ;
        RECT 66.320 19.350 67.580 19.490 ;
        RECT 66.320 19.290 66.640 19.350 ;
        RECT 67.290 19.310 67.580 19.350 ;
        RECT 72.090 19.490 72.380 19.540 ;
        RECT 72.560 19.490 72.880 19.550 ;
        RECT 76.400 19.490 76.720 19.550 ;
        RECT 86.000 19.490 86.320 19.550 ;
        RECT 97.520 19.490 97.840 19.550 ;
        RECT 72.090 19.350 72.880 19.490 ;
        RECT 76.200 19.350 76.720 19.490 ;
        RECT 85.800 19.350 86.320 19.490 ;
        RECT 97.320 19.350 97.840 19.490 ;
        RECT 72.090 19.310 72.380 19.350 ;
        RECT 72.560 19.290 72.880 19.350 ;
        RECT 76.400 19.290 76.720 19.350 ;
        RECT 86.000 19.290 86.320 19.350 ;
        RECT 97.520 19.290 97.840 19.350 ;
        RECT 105.680 19.490 106.000 19.550 ;
        RECT 106.170 19.490 106.460 19.540 ;
        RECT 105.680 19.350 106.460 19.490 ;
        RECT 105.680 19.290 106.000 19.350 ;
        RECT 106.170 19.310 106.460 19.350 ;
        RECT 117.690 19.490 117.980 19.540 ;
        RECT 118.160 19.490 118.480 19.550 ;
        RECT 117.690 19.350 118.480 19.490 ;
        RECT 117.690 19.310 117.980 19.350 ;
        RECT 118.160 19.290 118.480 19.350 ;
        RECT 28.890 19.120 29.180 19.170 ;
        RECT 64.400 19.120 64.720 19.180 ;
        RECT 94.160 19.120 94.480 19.180 ;
        RECT 28.890 18.980 64.720 19.120 ;
        RECT 93.960 18.980 94.480 19.120 ;
        RECT 28.890 18.940 29.180 18.980 ;
        RECT 64.400 18.920 64.720 18.980 ;
        RECT 94.160 18.920 94.480 18.980 ;
        RECT 109.040 19.120 109.360 19.180 ;
        RECT 114.330 19.120 114.620 19.170 ;
        RECT 109.040 18.980 114.620 19.120 ;
        RECT 109.040 18.920 109.360 18.980 ;
        RECT 114.330 18.940 114.620 18.980 ;
        RECT 38.010 18.570 38.300 18.800 ;
        RECT 56.730 18.750 57.020 18.800 ;
        RECT 57.200 18.750 57.520 18.810 ;
        RECT 59.600 18.750 59.920 18.810 ;
        RECT 56.730 18.610 57.520 18.750 ;
        RECT 59.400 18.610 59.920 18.750 ;
        RECT 56.730 18.570 57.020 18.610 ;
        RECT 33.200 18.380 33.520 18.440 ;
        RECT 33.000 18.240 33.520 18.380 ;
        RECT 33.200 18.180 33.520 18.240 ;
        RECT 37.520 18.380 37.840 18.440 ;
        RECT 38.090 18.380 38.230 18.570 ;
        RECT 57.200 18.550 57.520 18.610 ;
        RECT 59.600 18.550 59.920 18.610 ;
        RECT 65.840 18.750 66.160 18.810 ;
        RECT 66.330 18.750 66.620 18.800 ;
        RECT 67.280 18.750 67.600 18.810 ;
        RECT 77.840 18.750 78.160 18.810 ;
        RECT 65.840 18.610 66.620 18.750 ;
        RECT 67.080 18.610 67.600 18.750 ;
        RECT 77.640 18.610 78.160 18.750 ;
        RECT 65.840 18.550 66.160 18.610 ;
        RECT 66.330 18.570 66.620 18.610 ;
        RECT 67.280 18.550 67.600 18.610 ;
        RECT 77.840 18.550 78.160 18.610 ;
        RECT 37.520 18.240 38.230 18.380 ;
        RECT 39.440 18.380 39.760 18.440 ;
        RECT 41.370 18.380 41.660 18.430 ;
        RECT 45.690 18.380 45.980 18.430 ;
        RECT 39.440 18.240 45.980 18.380 ;
        RECT 37.520 18.180 37.840 18.240 ;
        RECT 39.440 18.180 39.760 18.240 ;
        RECT 41.370 18.200 41.660 18.240 ;
        RECT 15.440 17.640 15.760 17.700 ;
        RECT 34.650 17.640 34.940 17.690 ;
        RECT 42.800 17.640 43.120 17.700 ;
        RECT 15.440 17.500 34.940 17.640 ;
        RECT 42.600 17.500 43.120 17.640 ;
        RECT 15.440 17.440 15.760 17.500 ;
        RECT 34.650 17.460 34.940 17.500 ;
        RECT 42.800 17.440 43.120 17.500 ;
        RECT 24.080 17.270 24.400 17.330 ;
        RECT 26.010 17.270 26.300 17.320 ;
        RECT 30.330 17.270 30.620 17.320 ;
        RECT 24.080 17.130 30.620 17.270 ;
        RECT 24.080 17.070 24.400 17.130 ;
        RECT 26.010 17.090 26.300 17.130 ;
        RECT 30.330 17.090 30.620 17.130 ;
        RECT 38.970 17.270 39.260 17.320 ;
        RECT 41.840 17.270 42.160 17.330 ;
        RECT 38.970 17.130 42.160 17.270 ;
        RECT 44.810 17.270 44.950 18.240 ;
        RECT 45.690 18.200 45.980 18.240 ;
        RECT 46.170 18.200 46.460 18.430 ;
        RECT 48.570 18.380 48.860 18.430 ;
        RECT 50.970 18.380 51.260 18.430 ;
        RECT 48.570 18.240 51.260 18.380 ;
        RECT 48.570 18.200 48.860 18.240 ;
        RECT 50.970 18.200 51.260 18.240 ;
        RECT 51.440 18.380 51.760 18.440 ;
        RECT 52.880 18.380 53.200 18.440 ;
        RECT 63.440 18.380 63.760 18.440 ;
        RECT 68.720 18.380 69.040 18.440 ;
        RECT 69.680 18.380 70.000 18.440 ;
        RECT 51.440 18.240 51.960 18.380 ;
        RECT 52.680 18.240 53.200 18.380 ;
        RECT 63.240 18.240 63.760 18.380 ;
        RECT 68.520 18.240 69.040 18.380 ;
        RECT 69.480 18.240 70.000 18.380 ;
        RECT 45.200 18.010 45.520 18.070 ;
        RECT 46.250 18.010 46.390 18.200 ;
        RECT 51.440 18.180 51.760 18.240 ;
        RECT 52.880 18.180 53.200 18.240 ;
        RECT 63.440 18.180 63.760 18.240 ;
        RECT 68.720 18.180 69.040 18.240 ;
        RECT 69.680 18.180 70.000 18.240 ;
      LAYER met1 ;
        RECT 84.580 18.380 84.870 18.430 ;
        RECT 86.980 18.380 87.270 18.430 ;
        RECT 92.260 18.380 92.550 18.430 ;
        RECT 84.580 18.240 92.550 18.380 ;
        RECT 84.580 18.200 84.870 18.240 ;
        RECT 86.980 18.200 87.270 18.240 ;
        RECT 92.260 18.200 92.550 18.240 ;
        RECT 104.740 18.380 105.030 18.430 ;
        RECT 107.140 18.380 107.430 18.430 ;
        RECT 112.420 18.380 112.710 18.430 ;
        RECT 104.740 18.240 112.710 18.380 ;
        RECT 104.740 18.200 105.030 18.240 ;
        RECT 107.140 18.200 107.430 18.240 ;
        RECT 112.420 18.200 112.710 18.240 ;
      LAYER met1 ;
        RECT 45.200 17.870 46.390 18.010 ;
        RECT 48.090 18.010 48.380 18.060 ;
        RECT 48.090 17.870 86.230 18.010 ;
        RECT 45.200 17.810 45.520 17.870 ;
        RECT 48.090 17.830 48.380 17.870 ;
        RECT 45.680 17.640 46.000 17.700 ;
        RECT 47.610 17.640 47.900 17.690 ;
        RECT 45.680 17.500 47.900 17.640 ;
        RECT 45.680 17.440 46.000 17.500 ;
        RECT 47.610 17.460 47.900 17.500 ;
        RECT 64.400 17.640 64.720 17.700 ;
        RECT 66.800 17.640 67.120 17.700 ;
        RECT 64.400 17.500 67.120 17.640 ;
        RECT 86.090 17.640 86.230 17.870 ;
        RECT 106.160 17.640 106.480 17.700 ;
        RECT 86.090 17.500 106.480 17.640 ;
        RECT 64.400 17.440 64.720 17.500 ;
        RECT 66.800 17.440 67.120 17.500 ;
        RECT 106.160 17.440 106.480 17.500 ;
        RECT 48.570 17.270 48.860 17.320 ;
        RECT 44.810 17.130 48.860 17.270 ;
        RECT 38.970 17.090 39.260 17.130 ;
        RECT 41.840 17.070 42.160 17.130 ;
        RECT 48.570 17.090 48.860 17.130 ;
        RECT 53.370 17.270 53.660 17.320 ;
        RECT 53.840 17.270 54.160 17.330 ;
        RECT 53.370 17.130 54.160 17.270 ;
        RECT 53.370 17.090 53.660 17.130 ;
        RECT 53.840 17.070 54.160 17.130 ;
        RECT 41.840 15.790 42.160 15.850 ;
        RECT 64.400 15.790 64.720 15.850 ;
        RECT 41.840 15.650 64.720 15.790 ;
        RECT 41.840 15.590 42.160 15.650 ;
        RECT 64.400 15.590 64.720 15.650 ;
      LAYER via ;
        RECT 32.750 143.980 33.010 144.240 ;
        RECT 49.550 143.980 49.810 144.240 ;
        RECT 77.870 143.980 78.130 144.240 ;
        RECT 117.230 144.720 117.490 144.980 ;
        RECT 64.910 143.610 65.170 143.870 ;
        RECT 99.470 143.980 99.730 144.240 ;
        RECT 30.830 143.240 31.090 143.500 ;
        RECT 36.590 143.240 36.850 143.500 ;
        RECT 50.030 143.240 50.290 143.500 ;
        RECT 70.670 143.240 70.930 143.500 ;
        RECT 86.030 143.240 86.290 143.500 ;
        RECT 98.510 143.240 98.770 143.500 ;
        RECT 106.670 143.240 106.930 143.500 ;
        RECT 36.590 141.390 36.850 141.650 ;
        RECT 50.030 141.390 50.290 141.650 ;
        RECT 64.910 141.390 65.170 141.650 ;
        RECT 86.030 141.390 86.290 141.650 ;
        RECT 98.510 141.020 98.770 141.280 ;
        RECT 106.670 141.020 106.930 141.280 ;
        RECT 33.710 140.650 33.970 140.910 ;
        RECT 44.270 140.650 44.530 140.910 ;
        RECT 77.870 140.650 78.130 140.910 ;
        RECT 86.990 140.650 87.250 140.910 ;
        RECT 101.390 140.650 101.650 140.910 ;
        RECT 78.350 139.540 78.610 139.800 ;
        RECT 66.350 139.170 66.610 139.430 ;
        RECT 74.990 139.170 75.250 139.430 ;
        RECT 99.470 139.540 99.730 139.800 ;
        RECT 93.710 139.170 93.970 139.430 ;
        RECT 100.910 139.170 101.170 139.430 ;
        RECT 66.350 137.320 66.610 137.580 ;
        RECT 99.470 136.950 99.730 137.210 ;
        RECT 30.830 136.580 31.090 136.840 ;
        RECT 70.670 136.580 70.930 136.840 ;
        RECT 86.990 136.580 87.250 136.840 ;
        RECT 49.550 136.210 49.810 136.470 ;
        RECT 36.110 135.100 36.370 135.360 ;
        RECT 77.390 135.840 77.650 136.100 ;
        RECT 78.350 136.210 78.610 136.470 ;
        RECT 85.070 135.840 85.330 136.100 ;
        RECT 93.710 136.210 93.970 136.470 ;
        RECT 94.190 135.840 94.450 136.100 ;
        RECT 101.390 136.580 101.650 136.840 ;
        RECT 110.990 136.580 111.250 136.840 ;
        RECT 100.910 136.210 101.170 136.470 ;
        RECT 102.830 136.210 103.090 136.470 ;
        RECT 101.870 135.840 102.130 136.100 ;
        RECT 111.470 135.840 111.730 136.100 ;
        RECT 117.230 135.840 117.490 136.100 ;
        RECT 118.670 135.840 118.930 136.100 ;
        RECT 102.350 135.470 102.610 135.730 ;
        RECT 107.630 135.100 107.890 135.360 ;
        RECT 118.190 135.100 118.450 135.360 ;
        RECT 32.750 133.250 33.010 133.510 ;
        RECT 101.870 133.250 102.130 133.510 ;
        RECT 107.630 133.250 107.890 133.510 ;
        RECT 118.190 133.250 118.450 133.510 ;
        RECT 29.390 132.510 29.650 132.770 ;
        RECT 39.470 132.510 39.730 132.770 ;
        RECT 36.110 132.140 36.370 132.400 ;
        RECT 79.310 132.140 79.570 132.400 ;
        RECT 80.270 132.140 80.530 132.400 ;
        RECT 87.950 132.140 88.210 132.400 ;
        RECT 93.710 132.510 93.970 132.770 ;
        RECT 99.950 132.140 100.210 132.400 ;
        RECT 101.390 132.510 101.650 132.770 ;
        RECT 102.350 132.510 102.610 132.770 ;
        RECT 102.830 132.140 103.090 132.400 ;
        RECT 103.310 132.140 103.570 132.400 ;
        RECT 36.590 131.770 36.850 132.030 ;
        RECT 83.630 131.400 83.890 131.660 ;
        RECT 107.630 132.140 107.890 132.400 ;
        RECT 110.990 132.140 111.250 132.400 ;
        RECT 76.430 131.030 76.690 131.290 ;
        RECT 81.230 131.030 81.490 131.290 ;
        RECT 33.710 129.180 33.970 129.440 ;
        RECT 36.590 129.180 36.850 129.440 ;
        RECT 87.950 129.180 88.210 129.440 ;
        RECT 101.390 129.180 101.650 129.440 ;
        RECT 110.990 129.180 111.250 129.440 ;
        RECT 36.590 128.440 36.850 128.700 ;
        RECT 42.830 128.440 43.090 128.700 ;
        RECT 16.910 127.700 17.170 127.960 ;
        RECT 39.470 127.700 39.730 127.960 ;
        RECT 26.030 127.330 26.290 127.590 ;
        RECT 47.630 127.330 47.890 127.590 ;
        RECT 75.470 127.700 75.730 127.960 ;
        RECT 79.310 128.070 79.570 128.330 ;
        RECT 83.630 128.070 83.890 128.330 ;
        RECT 95.150 128.070 95.410 128.330 ;
        RECT 100.910 128.440 101.170 128.700 ;
        RECT 100.430 128.070 100.690 128.330 ;
        RECT 103.310 128.070 103.570 128.330 ;
        RECT 83.150 127.700 83.410 127.960 ;
        RECT 100.910 127.700 101.170 127.960 ;
        RECT 118.190 127.700 118.450 127.960 ;
        RECT 15.470 126.960 15.730 127.220 ;
        RECT 31.790 126.960 32.050 127.220 ;
        RECT 58.190 126.960 58.450 127.220 ;
        RECT 80.270 126.960 80.530 127.220 ;
        RECT 111.950 126.960 112.210 127.220 ;
        RECT 118.670 126.960 118.930 127.220 ;
        RECT 15.470 125.110 15.730 125.370 ;
        RECT 44.270 125.110 44.530 125.370 ;
        RECT 58.190 125.110 58.450 125.370 ;
        RECT 77.390 125.110 77.650 125.370 ;
        RECT 94.190 125.110 94.450 125.370 ;
        RECT 118.670 125.110 118.930 125.370 ;
        RECT 38.030 124.740 38.290 125.000 ;
        RECT 20.270 124.370 20.530 124.630 ;
        RECT 29.870 124.370 30.130 124.630 ;
        RECT 41.390 124.370 41.650 124.630 ;
        RECT 47.630 124.370 47.890 124.630 ;
        RECT 42.830 124.000 43.090 124.260 ;
        RECT 75.470 124.000 75.730 124.260 ;
        RECT 81.230 124.370 81.490 124.630 ;
        RECT 89.870 124.370 90.130 124.630 ;
        RECT 98.030 124.370 98.290 124.630 ;
        RECT 101.390 124.370 101.650 124.630 ;
        RECT 101.870 124.370 102.130 124.630 ;
        RECT 107.630 124.740 107.890 125.000 ;
        RECT 111.950 124.740 112.210 125.000 ;
        RECT 76.430 124.000 76.690 124.260 ;
        RECT 95.150 124.000 95.410 124.260 ;
        RECT 97.550 124.000 97.810 124.260 ;
        RECT 100.430 124.000 100.690 124.260 ;
        RECT 103.790 124.000 104.050 124.260 ;
        RECT 104.750 124.000 105.010 124.260 ;
        RECT 114.830 124.370 115.090 124.630 ;
        RECT 112.910 123.260 113.170 123.520 ;
        RECT 25.070 122.890 25.330 123.150 ;
        RECT 41.390 122.890 41.650 123.150 ;
        RECT 57.710 122.890 57.970 123.150 ;
        RECT 108.110 122.890 108.370 123.150 ;
        RECT 20.270 121.040 20.530 121.300 ;
        RECT 29.870 121.040 30.130 121.300 ;
        RECT 38.030 121.040 38.290 121.300 ;
        RECT 49.550 121.040 49.810 121.300 ;
        RECT 88.430 121.040 88.690 121.300 ;
        RECT 103.790 121.040 104.050 121.300 ;
        RECT 114.830 121.040 115.090 121.300 ;
        RECT 33.710 120.670 33.970 120.930 ;
        RECT 57.710 120.670 57.970 120.930 ;
        RECT 74.990 120.670 75.250 120.930 ;
        RECT 86.030 120.670 86.290 120.930 ;
        RECT 16.910 120.300 17.170 120.560 ;
        RECT 40.910 120.300 41.170 120.560 ;
        RECT 68.750 120.300 69.010 120.560 ;
        RECT 26.990 119.930 27.250 120.190 ;
        RECT 25.070 119.560 25.330 119.820 ;
        RECT 31.790 119.560 32.050 119.820 ;
        RECT 41.390 119.930 41.650 120.190 ;
        RECT 78.350 119.930 78.610 120.190 ;
        RECT 79.790 119.930 80.050 120.190 ;
        RECT 94.670 120.300 94.930 120.560 ;
        RECT 25.550 119.190 25.810 119.450 ;
        RECT 62.510 119.560 62.770 119.820 ;
        RECT 78.830 119.560 79.090 119.820 ;
        RECT 85.550 119.560 85.810 119.820 ;
        RECT 94.190 119.560 94.450 119.820 ;
        RECT 95.150 119.560 95.410 119.820 ;
        RECT 101.870 120.670 102.130 120.930 ;
        RECT 102.350 120.300 102.610 120.560 ;
        RECT 89.870 119.190 90.130 119.450 ;
        RECT 93.710 119.190 93.970 119.450 ;
        RECT 97.550 119.560 97.810 119.820 ;
        RECT 106.670 119.930 106.930 120.190 ;
        RECT 107.150 119.930 107.410 120.190 ;
        RECT 23.150 118.820 23.410 119.080 ;
        RECT 60.590 118.820 60.850 119.080 ;
        RECT 71.630 118.820 71.890 119.080 ;
        RECT 81.710 118.820 81.970 119.080 ;
        RECT 95.150 118.820 95.410 119.080 ;
        RECT 108.110 119.190 108.370 119.450 ;
        RECT 108.590 118.820 108.850 119.080 ;
        RECT 60.590 116.970 60.850 117.230 ;
        RECT 86.030 116.970 86.290 117.230 ;
        RECT 106.670 116.970 106.930 117.230 ;
        RECT 47.630 116.600 47.890 116.860 ;
        RECT 52.430 116.600 52.690 116.860 ;
        RECT 71.630 116.600 71.890 116.860 ;
        RECT 88.430 116.600 88.690 116.860 ;
        RECT 111.950 116.600 112.210 116.860 ;
        RECT 16.910 116.230 17.170 116.490 ;
        RECT 23.150 116.230 23.410 116.490 ;
        RECT 25.070 116.230 25.330 116.490 ;
        RECT 29.390 116.230 29.650 116.490 ;
        RECT 43.790 116.230 44.050 116.490 ;
        RECT 61.550 116.230 61.810 116.490 ;
        RECT 82.670 116.230 82.930 116.490 ;
        RECT 89.870 116.230 90.130 116.490 ;
        RECT 56.750 115.860 57.010 116.120 ;
        RECT 57.710 115.860 57.970 116.120 ;
        RECT 95.150 115.860 95.410 116.120 ;
        RECT 96.110 115.860 96.370 116.120 ;
        RECT 101.870 116.230 102.130 116.490 ;
        RECT 104.750 116.230 105.010 116.490 ;
        RECT 110.990 116.230 111.250 116.490 ;
        RECT 124.430 116.230 124.690 116.490 ;
        RECT 37.550 115.490 37.810 115.750 ;
        RECT 42.830 115.490 43.090 115.750 ;
        RECT 61.070 115.490 61.330 115.750 ;
        RECT 72.110 115.490 72.370 115.750 ;
        RECT 85.070 115.490 85.330 115.750 ;
        RECT 101.390 115.860 101.650 116.120 ;
        RECT 52.910 115.120 53.170 115.380 ;
        RECT 64.910 115.120 65.170 115.380 ;
        RECT 71.630 115.120 71.890 115.380 ;
        RECT 14.030 114.750 14.290 115.010 ;
        RECT 87.950 114.750 88.210 115.010 ;
        RECT 97.550 115.120 97.810 115.380 ;
        RECT 108.590 115.860 108.850 116.120 ;
        RECT 110.030 114.750 110.290 115.010 ;
        RECT 117.230 114.750 117.490 115.010 ;
        RECT 118.190 114.750 118.450 115.010 ;
        RECT 25.070 112.900 25.330 113.160 ;
        RECT 72.110 112.900 72.370 113.160 ;
        RECT 82.670 112.900 82.930 113.160 ;
        RECT 93.710 112.900 93.970 113.160 ;
        RECT 124.430 112.900 124.690 113.160 ;
        RECT 14.030 112.160 14.290 112.420 ;
        RECT 86.030 112.160 86.290 112.420 ;
        RECT 26.510 111.790 26.770 112.050 ;
        RECT 26.990 111.790 27.250 112.050 ;
        RECT 29.390 111.790 29.650 112.050 ;
        RECT 25.070 111.420 25.330 111.680 ;
        RECT 52.430 111.790 52.690 112.050 ;
        RECT 66.350 111.790 66.610 112.050 ;
        RECT 74.990 111.790 75.250 112.050 ;
        RECT 37.550 110.680 37.810 110.940 ;
        RECT 64.430 111.420 64.690 111.680 ;
        RECT 82.190 111.420 82.450 111.680 ;
        RECT 44.750 111.050 45.010 111.310 ;
        RECT 62.030 111.050 62.290 111.310 ;
        RECT 65.390 111.050 65.650 111.310 ;
        RECT 80.750 111.050 81.010 111.310 ;
        RECT 85.070 111.050 85.330 111.310 ;
        RECT 86.510 111.420 86.770 111.680 ;
        RECT 107.150 112.160 107.410 112.420 ;
        RECT 91.790 111.420 92.050 111.680 ;
        RECT 96.110 111.420 96.370 111.680 ;
        RECT 100.430 111.790 100.690 112.050 ;
        RECT 110.030 111.790 110.290 112.050 ;
        RECT 112.910 111.420 113.170 111.680 ;
        RECT 105.710 111.050 105.970 111.310 ;
        RECT 117.230 111.050 117.490 111.310 ;
        RECT 52.430 110.680 52.690 110.940 ;
        RECT 79.310 110.680 79.570 110.940 ;
        RECT 52.910 108.830 53.170 109.090 ;
        RECT 83.630 108.830 83.890 109.090 ;
        RECT 85.070 108.830 85.330 109.090 ;
        RECT 61.070 108.460 61.330 108.720 ;
        RECT 69.230 108.460 69.490 108.720 ;
        RECT 23.150 108.090 23.410 108.350 ;
        RECT 24.110 108.090 24.370 108.350 ;
        RECT 26.990 108.090 27.250 108.350 ;
        RECT 31.790 108.090 32.050 108.350 ;
        RECT 32.270 108.090 32.530 108.350 ;
        RECT 26.510 107.720 26.770 107.980 ;
        RECT 65.390 107.720 65.650 107.980 ;
        RECT 79.310 108.090 79.570 108.350 ;
        RECT 82.670 108.090 82.930 108.350 ;
        RECT 87.950 108.090 88.210 108.350 ;
        RECT 107.150 108.830 107.410 109.090 ;
        RECT 113.870 108.830 114.130 109.090 ;
        RECT 118.190 108.830 118.450 109.090 ;
        RECT 91.790 108.460 92.050 108.720 ;
        RECT 108.590 108.460 108.850 108.720 ;
        RECT 123.950 108.460 124.210 108.720 ;
        RECT 109.070 108.090 109.330 108.350 ;
        RECT 61.550 106.980 61.810 107.240 ;
        RECT 80.750 107.720 81.010 107.980 ;
        RECT 81.710 107.720 81.970 107.980 ;
        RECT 85.550 107.720 85.810 107.980 ;
        RECT 86.030 107.720 86.290 107.980 ;
        RECT 94.670 107.720 94.930 107.980 ;
        RECT 100.430 107.720 100.690 107.980 ;
        RECT 102.350 107.720 102.610 107.980 ;
        RECT 103.310 107.720 103.570 107.980 ;
        RECT 85.070 107.350 85.330 107.610 ;
        RECT 13.070 106.610 13.330 106.870 ;
        RECT 55.310 106.610 55.570 106.870 ;
        RECT 72.110 106.610 72.370 106.870 ;
        RECT 79.790 106.610 80.050 106.870 ;
        RECT 86.510 106.980 86.770 107.240 ;
        RECT 109.070 106.610 109.330 106.870 ;
        RECT 117.710 106.610 117.970 106.870 ;
        RECT 26.510 104.760 26.770 105.020 ;
        RECT 32.270 104.760 32.530 105.020 ;
        RECT 37.550 104.760 37.810 105.020 ;
        RECT 61.550 104.760 61.810 105.020 ;
        RECT 85.550 104.760 85.810 105.020 ;
        RECT 98.030 104.760 98.290 105.020 ;
        RECT 13.070 103.280 13.330 103.540 ;
        RECT 43.790 103.650 44.050 103.910 ;
        RECT 44.750 103.650 45.010 103.910 ;
        RECT 52.430 103.650 52.690 103.910 ;
        RECT 40.910 103.280 41.170 103.540 ;
        RECT 54.350 103.280 54.610 103.540 ;
        RECT 21.230 102.910 21.490 103.170 ;
        RECT 57.230 102.910 57.490 103.170 ;
        RECT 117.710 104.020 117.970 104.280 ;
        RECT 85.070 103.650 85.330 103.910 ;
        RECT 92.750 103.650 93.010 103.910 ;
        RECT 94.190 103.650 94.450 103.910 ;
        RECT 109.550 103.650 109.810 103.910 ;
        RECT 117.230 103.650 117.490 103.910 ;
        RECT 125.390 103.650 125.650 103.910 ;
        RECT 58.190 102.910 58.450 103.170 ;
        RECT 79.790 103.280 80.050 103.540 ;
        RECT 82.190 103.280 82.450 103.540 ;
        RECT 85.550 103.280 85.810 103.540 ;
        RECT 101.390 103.280 101.650 103.540 ;
        RECT 102.350 103.280 102.610 103.540 ;
        RECT 105.710 103.280 105.970 103.540 ;
        RECT 111.470 103.280 111.730 103.540 ;
        RECT 65.390 102.910 65.650 103.170 ;
        RECT 76.430 102.910 76.690 103.170 ;
        RECT 124.910 102.910 125.170 103.170 ;
        RECT 21.230 100.690 21.490 100.950 ;
        RECT 65.390 100.690 65.650 100.950 ;
        RECT 78.350 100.690 78.610 100.950 ;
        RECT 81.230 100.690 81.490 100.950 ;
        RECT 83.150 100.690 83.410 100.950 ;
        RECT 31.790 100.320 32.050 100.580 ;
        RECT 43.310 100.320 43.570 100.580 ;
        RECT 53.870 100.320 54.130 100.580 ;
        RECT 74.990 100.320 75.250 100.580 ;
        RECT 22.190 99.950 22.450 100.210 ;
        RECT 33.710 99.950 33.970 100.210 ;
        RECT 52.430 99.950 52.690 100.210 ;
        RECT 56.750 99.950 57.010 100.210 ;
        RECT 57.710 99.580 57.970 99.840 ;
        RECT 61.070 99.950 61.330 100.210 ;
        RECT 62.030 99.950 62.290 100.210 ;
        RECT 62.510 99.580 62.770 99.840 ;
        RECT 54.350 99.210 54.610 99.470 ;
        RECT 57.230 99.210 57.490 99.470 ;
        RECT 68.750 99.580 69.010 99.840 ;
        RECT 72.590 99.580 72.850 99.840 ;
        RECT 75.470 99.950 75.730 100.210 ;
        RECT 100.910 100.320 101.170 100.580 ;
        RECT 102.350 100.320 102.610 100.580 ;
        RECT 101.390 99.950 101.650 100.210 ;
        RECT 110.990 100.320 111.250 100.580 ;
        RECT 104.270 99.950 104.530 100.210 ;
        RECT 107.630 99.950 107.890 100.210 ;
        RECT 113.870 99.950 114.130 100.210 ;
        RECT 118.190 99.950 118.450 100.210 ;
        RECT 125.390 99.950 125.650 100.210 ;
        RECT 67.310 99.210 67.570 99.470 ;
        RECT 101.870 99.580 102.130 99.840 ;
        RECT 123.950 99.580 124.210 99.840 ;
        RECT 93.230 99.210 93.490 99.470 ;
        RECT 116.750 99.210 117.010 99.470 ;
        RECT 58.190 98.840 58.450 99.100 ;
        RECT 100.430 98.840 100.690 99.100 ;
        RECT 14.510 98.470 14.770 98.730 ;
        RECT 23.150 98.470 23.410 98.730 ;
        RECT 30.350 98.470 30.610 98.730 ;
        RECT 54.830 98.470 55.090 98.730 ;
        RECT 69.230 98.470 69.490 98.730 ;
        RECT 117.230 98.840 117.490 99.100 ;
        RECT 22.190 96.620 22.450 96.880 ;
        RECT 33.710 96.620 33.970 96.880 ;
        RECT 43.790 96.620 44.050 96.880 ;
        RECT 54.830 96.620 55.090 96.880 ;
        RECT 30.350 96.250 30.610 96.510 ;
        RECT 56.750 96.250 57.010 96.510 ;
        RECT 66.350 96.620 66.610 96.880 ;
        RECT 67.310 96.620 67.570 96.880 ;
        RECT 76.430 96.620 76.690 96.880 ;
        RECT 101.390 96.620 101.650 96.880 ;
        RECT 103.310 96.620 103.570 96.880 ;
        RECT 104.270 96.620 104.530 96.880 ;
        RECT 116.750 96.620 117.010 96.880 ;
        RECT 117.230 96.620 117.490 96.880 ;
        RECT 64.430 96.250 64.690 96.510 ;
        RECT 86.030 96.250 86.290 96.510 ;
        RECT 23.150 95.880 23.410 96.140 ;
        RECT 24.110 95.510 24.370 95.770 ;
        RECT 25.550 95.140 25.810 95.400 ;
        RECT 26.990 95.510 27.250 95.770 ;
        RECT 61.070 95.880 61.330 96.140 ;
        RECT 89.870 96.250 90.130 96.510 ;
        RECT 43.310 95.510 43.570 95.770 ;
        RECT 52.430 95.510 52.690 95.770 ;
        RECT 52.910 95.510 53.170 95.770 ;
        RECT 28.430 95.140 28.690 95.400 ;
        RECT 36.590 95.140 36.850 95.400 ;
        RECT 57.710 95.510 57.970 95.770 ;
        RECT 86.990 95.880 87.250 96.140 ;
        RECT 72.110 95.140 72.370 95.400 ;
        RECT 52.910 94.770 53.170 95.030 ;
        RECT 57.230 94.770 57.490 95.030 ;
        RECT 8.750 94.400 9.010 94.660 ;
        RECT 36.110 94.400 36.370 94.660 ;
        RECT 62.030 94.400 62.290 94.660 ;
        RECT 79.310 95.140 79.570 95.400 ;
        RECT 78.830 94.770 79.090 95.030 ;
        RECT 81.230 94.770 81.490 95.030 ;
        RECT 84.110 94.400 84.370 94.660 ;
        RECT 90.350 95.510 90.610 95.770 ;
        RECT 93.230 95.510 93.490 95.770 ;
        RECT 86.510 95.140 86.770 95.400 ;
        RECT 87.950 94.770 88.210 95.030 ;
        RECT 93.230 94.770 93.490 95.030 ;
        RECT 108.110 95.510 108.370 95.770 ;
        RECT 108.590 95.510 108.850 95.770 ;
        RECT 107.630 95.140 107.890 95.400 ;
        RECT 123.950 95.510 124.210 95.770 ;
        RECT 100.910 94.770 101.170 95.030 ;
        RECT 109.550 94.770 109.810 95.030 ;
        RECT 132.110 94.770 132.370 95.030 ;
        RECT 8.750 92.550 9.010 92.810 ;
        RECT 21.710 92.550 21.970 92.810 ;
        RECT 36.110 92.550 36.370 92.810 ;
        RECT 25.550 92.180 25.810 92.440 ;
        RECT 24.110 91.810 24.370 92.070 ;
        RECT 28.430 91.810 28.690 92.070 ;
        RECT 26.990 91.440 27.250 91.700 ;
        RECT 62.030 92.180 62.290 92.440 ;
        RECT 92.750 92.550 93.010 92.810 ;
        RECT 101.870 92.550 102.130 92.810 ;
        RECT 107.150 92.550 107.410 92.810 ;
        RECT 90.350 92.180 90.610 92.440 ;
        RECT 53.390 91.810 53.650 92.070 ;
        RECT 57.710 91.810 57.970 92.070 ;
        RECT 79.310 91.810 79.570 92.070 ;
        RECT 97.550 91.810 97.810 92.070 ;
        RECT 102.350 91.810 102.610 92.070 ;
        RECT 110.990 92.550 111.250 92.810 ;
        RECT 123.950 92.180 124.210 92.440 ;
        RECT 117.710 91.810 117.970 92.070 ;
        RECT 72.110 91.440 72.370 91.700 ;
        RECT 79.790 91.440 80.050 91.700 ;
        RECT 85.550 91.440 85.810 91.700 ;
        RECT 92.270 91.440 92.530 91.700 ;
        RECT 92.750 91.440 93.010 91.700 ;
        RECT 29.390 91.070 29.650 91.330 ;
        RECT 35.150 91.070 35.410 91.330 ;
        RECT 63.950 91.070 64.210 91.330 ;
        RECT 108.110 91.440 108.370 91.700 ;
        RECT 124.910 91.440 125.170 91.700 ;
        RECT 110.510 91.070 110.770 91.330 ;
        RECT 28.430 90.700 28.690 90.960 ;
        RECT 120.590 90.700 120.850 90.960 ;
        RECT 14.510 90.330 14.770 90.590 ;
        RECT 34.670 90.330 34.930 90.590 ;
        RECT 71.150 90.330 71.410 90.590 ;
        RECT 26.990 88.480 27.250 88.740 ;
        RECT 53.390 88.480 53.650 88.740 ;
        RECT 57.710 88.480 57.970 88.740 ;
        RECT 63.950 88.480 64.210 88.740 ;
        RECT 64.430 88.480 64.690 88.740 ;
        RECT 86.510 88.480 86.770 88.740 ;
        RECT 107.150 88.480 107.410 88.740 ;
        RECT 118.190 88.480 118.450 88.740 ;
        RECT 29.390 88.110 29.650 88.370 ;
        RECT 29.390 87.370 29.650 87.630 ;
        RECT 33.710 87.740 33.970 88.000 ;
        RECT 31.790 87.000 32.050 87.260 ;
        RECT 49.070 87.370 49.330 87.630 ;
        RECT 53.870 87.370 54.130 87.630 ;
        RECT 55.310 87.370 55.570 87.630 ;
        RECT 59.150 87.370 59.410 87.630 ;
        RECT 34.670 86.630 34.930 86.890 ;
        RECT 35.150 86.630 35.410 86.890 ;
        RECT 52.910 87.000 53.170 87.260 ;
        RECT 60.110 87.000 60.370 87.260 ;
        RECT 98.990 87.740 99.250 88.000 ;
        RECT 86.510 87.370 86.770 87.630 ;
        RECT 87.950 87.370 88.210 87.630 ;
        RECT 97.550 87.370 97.810 87.630 ;
        RECT 103.310 87.370 103.570 87.630 ;
        RECT 26.030 86.260 26.290 86.520 ;
        RECT 71.150 86.630 71.410 86.890 ;
        RECT 92.270 87.000 92.530 87.260 ;
        RECT 100.430 87.000 100.690 87.260 ;
        RECT 110.510 87.370 110.770 87.630 ;
        RECT 120.590 87.000 120.850 87.260 ;
        RECT 80.270 86.630 80.530 86.890 ;
        RECT 74.990 86.260 75.250 86.520 ;
        RECT 104.270 86.260 104.530 86.520 ;
        RECT 113.390 86.260 113.650 86.520 ;
        RECT 21.710 84.410 21.970 84.670 ;
        RECT 24.110 84.410 24.370 84.670 ;
        RECT 19.310 84.040 19.570 84.300 ;
        RECT 19.790 84.040 20.050 84.300 ;
        RECT 49.550 84.410 49.810 84.670 ;
        RECT 32.270 84.040 32.530 84.300 ;
        RECT 72.110 84.040 72.370 84.300 ;
        RECT 29.870 83.670 30.130 83.930 ;
        RECT 34.670 83.670 34.930 83.930 ;
        RECT 36.590 83.670 36.850 83.930 ;
        RECT 45.230 83.670 45.490 83.930 ;
        RECT 74.990 84.040 75.250 84.300 ;
        RECT 31.790 83.300 32.050 83.560 ;
        RECT 35.150 83.300 35.410 83.560 ;
        RECT 44.270 83.300 44.530 83.560 ;
        RECT 59.630 83.300 59.890 83.560 ;
        RECT 79.310 84.040 79.570 84.300 ;
        RECT 107.630 84.410 107.890 84.670 ;
        RECT 113.390 84.410 113.650 84.670 ;
        RECT 86.510 84.040 86.770 84.300 ;
        RECT 84.590 83.670 84.850 83.930 ;
        RECT 111.950 84.040 112.210 84.300 ;
        RECT 114.830 84.040 115.090 84.300 ;
        RECT 101.390 83.670 101.650 83.930 ;
        RECT 31.310 82.560 31.570 82.820 ;
        RECT 50.510 82.560 50.770 82.820 ;
        RECT 91.790 83.300 92.050 83.560 ;
        RECT 85.070 82.930 85.330 83.190 ;
        RECT 91.790 82.560 92.050 82.820 ;
        RECT 30.830 82.190 31.090 82.450 ;
        RECT 35.150 82.190 35.410 82.450 ;
        RECT 36.110 82.190 36.370 82.450 ;
        RECT 64.910 82.190 65.170 82.450 ;
        RECT 79.790 82.190 80.050 82.450 ;
        RECT 90.830 82.190 91.090 82.450 ;
        RECT 19.310 80.340 19.570 80.600 ;
        RECT 29.390 80.340 29.650 80.600 ;
        RECT 60.110 80.340 60.370 80.600 ;
        RECT 79.790 80.340 80.050 80.600 ;
        RECT 103.310 80.340 103.570 80.600 ;
        RECT 114.830 80.340 115.090 80.600 ;
        RECT 116.270 80.340 116.530 80.600 ;
        RECT 72.110 79.970 72.370 80.230 ;
        RECT 95.150 79.970 95.410 80.230 ;
        RECT 101.390 79.970 101.650 80.230 ;
        RECT 35.150 79.600 35.410 79.860 ;
        RECT 70.670 79.230 70.930 79.490 ;
        RECT 104.270 79.600 104.530 79.860 ;
        RECT 14.510 78.860 14.770 79.120 ;
        RECT 22.670 78.860 22.930 79.120 ;
        RECT 30.830 78.860 31.090 79.120 ;
        RECT 31.310 78.860 31.570 79.120 ;
        RECT 70.190 78.860 70.450 79.120 ;
        RECT 71.630 78.860 71.890 79.120 ;
        RECT 72.590 78.490 72.850 78.750 ;
        RECT 85.070 79.230 85.330 79.490 ;
        RECT 91.790 79.230 92.050 79.490 ;
        RECT 95.150 79.230 95.410 79.490 ;
        RECT 100.430 79.230 100.690 79.490 ;
        RECT 130.670 79.600 130.930 79.860 ;
        RECT 84.110 78.490 84.370 78.750 ;
        RECT 91.790 78.490 92.050 78.750 ;
        RECT 21.710 78.120 21.970 78.380 ;
        RECT 45.710 78.120 45.970 78.380 ;
        RECT 84.590 78.120 84.850 78.380 ;
        RECT 102.350 78.490 102.610 78.750 ;
        RECT 116.270 79.230 116.530 79.490 ;
        RECT 107.150 78.490 107.410 78.750 ;
        RECT 108.110 78.120 108.370 78.380 ;
        RECT 114.830 78.120 115.090 78.380 ;
        RECT 119.150 78.120 119.410 78.380 ;
        RECT 123.470 78.120 123.730 78.380 ;
        RECT 21.710 76.270 21.970 76.530 ;
        RECT 45.710 76.270 45.970 76.530 ;
        RECT 65.390 76.270 65.650 76.530 ;
        RECT 31.790 75.900 32.050 76.160 ;
        RECT 43.790 75.900 44.050 76.160 ;
        RECT 71.150 75.900 71.410 76.160 ;
        RECT 72.590 75.900 72.850 76.160 ;
        RECT 114.830 76.270 115.090 76.530 ;
        RECT 119.150 76.270 119.410 76.530 ;
        RECT 82.670 75.900 82.930 76.160 ;
        RECT 44.750 75.530 45.010 75.790 ;
        RECT 47.630 75.530 47.890 75.790 ;
        RECT 60.110 75.530 60.370 75.790 ;
        RECT 79.310 75.530 79.570 75.790 ;
        RECT 84.590 75.530 84.850 75.790 ;
        RECT 101.390 75.900 101.650 76.160 ;
        RECT 104.270 75.900 104.530 76.160 ;
        RECT 123.470 75.900 123.730 76.160 ;
        RECT 93.710 75.530 93.970 75.790 ;
        RECT 96.590 75.530 96.850 75.790 ;
        RECT 108.110 75.530 108.370 75.790 ;
        RECT 110.030 75.530 110.290 75.790 ;
        RECT 116.750 75.530 117.010 75.790 ;
        RECT 29.390 75.160 29.650 75.420 ;
        RECT 36.590 75.160 36.850 75.420 ;
        RECT 43.310 75.160 43.570 75.420 ;
        RECT 58.190 75.160 58.450 75.420 ;
        RECT 85.070 75.160 85.330 75.420 ;
        RECT 85.550 75.160 85.810 75.420 ;
        RECT 90.830 75.160 91.090 75.420 ;
        RECT 98.990 75.160 99.250 75.420 ;
        RECT 100.430 75.160 100.690 75.420 ;
        RECT 102.350 74.790 102.610 75.050 ;
        RECT 116.270 74.790 116.530 75.050 ;
        RECT 116.750 74.790 117.010 75.050 ;
        RECT 137.390 74.790 137.650 75.050 ;
        RECT 22.670 74.050 22.930 74.310 ;
        RECT 55.790 74.050 56.050 74.310 ;
        RECT 79.310 74.050 79.570 74.310 ;
        RECT 90.830 74.050 91.090 74.310 ;
        RECT 10.670 72.200 10.930 72.460 ;
        RECT 19.790 72.200 20.050 72.460 ;
        RECT 36.110 72.200 36.370 72.460 ;
        RECT 85.070 72.200 85.330 72.460 ;
        RECT 93.710 72.200 93.970 72.460 ;
        RECT 102.350 72.200 102.610 72.460 ;
        RECT 47.630 71.830 47.890 72.090 ;
        RECT 57.230 71.830 57.490 72.090 ;
        RECT 29.870 71.460 30.130 71.720 ;
        RECT 21.710 70.350 21.970 70.610 ;
        RECT 26.510 70.720 26.770 70.980 ;
        RECT 30.350 71.090 30.610 71.350 ;
        RECT 45.230 71.460 45.490 71.720 ;
        RECT 46.670 71.460 46.930 71.720 ;
        RECT 49.070 71.460 49.330 71.720 ;
        RECT 32.750 70.720 33.010 70.980 ;
        RECT 43.790 71.090 44.050 71.350 ;
        RECT 54.350 71.090 54.610 71.350 ;
        RECT 48.110 70.720 48.370 70.980 ;
        RECT 64.430 71.090 64.690 71.350 ;
        RECT 74.990 71.090 75.250 71.350 ;
        RECT 79.310 71.090 79.570 71.350 ;
        RECT 68.270 70.720 68.530 70.980 ;
        RECT 70.670 70.720 70.930 70.980 ;
        RECT 76.910 70.720 77.170 70.980 ;
        RECT 30.830 70.350 31.090 70.610 ;
        RECT 31.310 70.350 31.570 70.610 ;
        RECT 19.310 69.980 19.570 70.240 ;
        RECT 47.630 69.980 47.890 70.240 ;
        RECT 49.550 70.350 49.810 70.610 ;
        RECT 61.550 70.350 61.810 70.610 ;
        RECT 84.110 70.350 84.370 70.610 ;
        RECT 59.630 69.980 59.890 70.240 ;
        RECT 86.990 71.090 87.250 71.350 ;
        RECT 103.310 71.460 103.570 71.720 ;
        RECT 105.710 71.460 105.970 71.720 ;
        RECT 101.390 71.090 101.650 71.350 ;
        RECT 99.950 70.720 100.210 70.980 ;
        RECT 101.870 70.720 102.130 70.980 ;
        RECT 102.830 70.720 103.090 70.980 ;
        RECT 106.670 71.830 106.930 72.090 ;
        RECT 130.670 71.830 130.930 72.090 ;
        RECT 108.590 71.090 108.850 71.350 ;
        RECT 91.790 70.350 92.050 70.610 ;
        RECT 98.510 70.350 98.770 70.610 ;
        RECT 113.390 71.090 113.650 71.350 ;
        RECT 112.910 70.720 113.170 70.980 ;
        RECT 115.790 70.720 116.050 70.980 ;
        RECT 120.590 70.720 120.850 70.980 ;
        RECT 133.070 70.350 133.330 70.610 ;
        RECT 93.230 69.980 93.490 70.240 ;
        RECT 106.670 69.980 106.930 70.240 ;
        RECT 117.230 69.980 117.490 70.240 ;
        RECT 118.190 69.980 118.450 70.240 ;
        RECT 134.990 69.980 135.250 70.240 ;
        RECT 10.670 67.390 10.930 67.650 ;
        RECT 19.310 68.130 19.570 68.390 ;
        RECT 69.710 68.130 69.970 68.390 ;
        RECT 79.310 68.130 79.570 68.390 ;
        RECT 82.670 68.130 82.930 68.390 ;
        RECT 85.550 68.130 85.810 68.390 ;
        RECT 21.230 67.760 21.490 68.020 ;
        RECT 42.830 67.760 43.090 68.020 ;
        RECT 53.870 67.760 54.130 68.020 ;
        RECT 58.190 67.760 58.450 68.020 ;
        RECT 15.470 67.390 15.730 67.650 ;
        RECT 18.830 67.390 19.090 67.650 ;
        RECT 26.030 67.020 26.290 67.280 ;
        RECT 26.990 67.390 27.250 67.650 ;
        RECT 35.630 67.390 35.890 67.650 ;
        RECT 36.590 67.390 36.850 67.650 ;
        RECT 38.990 67.390 39.250 67.650 ;
        RECT 57.710 67.390 57.970 67.650 ;
        RECT 80.270 67.760 80.530 68.020 ;
        RECT 32.750 67.020 33.010 67.280 ;
        RECT 42.830 67.020 43.090 67.280 ;
        RECT 50.030 67.020 50.290 67.280 ;
        RECT 61.550 67.020 61.810 67.280 ;
        RECT 76.910 67.390 77.170 67.650 ;
        RECT 74.990 67.020 75.250 67.280 ;
        RECT 84.110 67.390 84.370 67.650 ;
        RECT 97.550 68.130 97.810 68.390 ;
        RECT 108.590 68.130 108.850 68.390 ;
        RECT 110.990 68.130 111.250 68.390 ;
        RECT 113.390 68.130 113.650 68.390 ;
        RECT 130.670 68.130 130.930 68.390 ;
        RECT 90.830 67.760 91.090 68.020 ;
        RECT 102.830 67.760 103.090 68.020 ;
        RECT 107.150 67.760 107.410 68.020 ;
        RECT 94.670 67.390 94.930 67.650 ;
        RECT 135.950 67.760 136.210 68.020 ;
        RECT 19.310 66.280 19.570 66.540 ;
        RECT 75.470 66.650 75.730 66.910 ;
        RECT 92.750 66.650 93.010 66.910 ;
        RECT 95.150 66.650 95.410 66.910 ;
        RECT 115.310 67.390 115.570 67.650 ;
        RECT 117.230 67.390 117.490 67.650 ;
        RECT 132.110 67.390 132.370 67.650 ;
        RECT 138.350 67.390 138.610 67.650 ;
        RECT 53.390 66.280 53.650 66.540 ;
        RECT 80.270 66.280 80.530 66.540 ;
        RECT 111.950 66.280 112.210 66.540 ;
        RECT 116.750 67.020 117.010 67.280 ;
        RECT 139.310 67.020 139.570 67.280 ;
        RECT 129.710 66.280 129.970 66.540 ;
        RECT 21.710 65.910 21.970 66.170 ;
        RECT 50.510 65.910 50.770 66.170 ;
        RECT 100.910 65.910 101.170 66.170 ;
        RECT 124.910 65.910 125.170 66.170 ;
        RECT 129.230 65.910 129.490 66.170 ;
        RECT 6.350 63.320 6.610 63.580 ;
        RECT 13.070 63.320 13.330 63.580 ;
        RECT 8.750 62.950 9.010 63.210 ;
        RECT 9.230 62.950 9.490 63.210 ;
        RECT 55.790 64.060 56.050 64.320 ;
        RECT 68.270 64.060 68.530 64.320 ;
        RECT 69.710 64.060 69.970 64.320 ;
        RECT 70.190 64.060 70.450 64.320 ;
        RECT 14.030 62.580 14.290 62.840 ;
        RECT 17.390 62.580 17.650 62.840 ;
        RECT 26.510 63.690 26.770 63.950 ;
        RECT 19.310 63.320 19.570 63.580 ;
        RECT 50.510 63.320 50.770 63.580 ;
        RECT 14.510 62.210 14.770 62.470 ;
        RECT 23.150 62.950 23.410 63.210 ;
        RECT 38.030 62.950 38.290 63.210 ;
        RECT 71.630 63.690 71.890 63.950 ;
        RECT 29.870 62.580 30.130 62.840 ;
        RECT 46.670 62.210 46.930 62.470 ;
        RECT 57.230 62.210 57.490 62.470 ;
        RECT 18.830 61.840 19.090 62.100 ;
        RECT 36.110 61.840 36.370 62.100 ;
        RECT 38.510 61.840 38.770 62.100 ;
        RECT 39.470 61.840 39.730 62.100 ;
        RECT 57.710 61.840 57.970 62.100 ;
        RECT 72.110 62.950 72.370 63.210 ;
        RECT 82.670 64.060 82.930 64.320 ;
        RECT 86.990 64.060 87.250 64.320 ;
        RECT 100.910 64.060 101.170 64.320 ;
        RECT 138.350 64.060 138.610 64.320 ;
        RECT 87.950 62.950 88.210 63.210 ;
        RECT 95.150 62.950 95.410 63.210 ;
        RECT 71.630 62.580 71.890 62.840 ;
        RECT 75.470 62.580 75.730 62.840 ;
        RECT 71.150 62.210 71.410 62.470 ;
        RECT 72.110 62.210 72.370 62.470 ;
        RECT 77.870 61.840 78.130 62.100 ;
        RECT 87.470 62.580 87.730 62.840 ;
        RECT 86.990 62.210 87.250 62.470 ;
        RECT 98.030 62.210 98.290 62.470 ;
        RECT 99.470 62.580 99.730 62.840 ;
        RECT 100.430 62.580 100.690 62.840 ;
        RECT 112.910 62.210 113.170 62.470 ;
        RECT 118.190 62.210 118.450 62.470 ;
        RECT 134.990 62.210 135.250 62.470 ;
        RECT 98.510 61.840 98.770 62.100 ;
        RECT 107.150 61.840 107.410 62.100 ;
        RECT 136.910 61.840 137.170 62.100 ;
        RECT 23.630 59.990 23.890 60.250 ;
        RECT 29.390 59.990 29.650 60.250 ;
        RECT 64.910 59.990 65.170 60.250 ;
        RECT 71.630 59.990 71.890 60.250 ;
        RECT 107.150 59.990 107.410 60.250 ;
        RECT 17.390 59.620 17.650 59.880 ;
        RECT 19.310 59.620 19.570 59.880 ;
        RECT 38.030 59.620 38.290 59.880 ;
        RECT 52.430 59.620 52.690 59.880 ;
        RECT 53.390 59.620 53.650 59.880 ;
        RECT 29.870 59.250 30.130 59.510 ;
        RECT 9.230 58.510 9.490 58.770 ;
        RECT 30.350 58.510 30.610 58.770 ;
        RECT 46.670 58.880 46.930 59.140 ;
        RECT 42.830 58.510 43.090 58.770 ;
        RECT 53.870 58.880 54.130 59.140 ;
        RECT 54.350 58.880 54.610 59.140 ;
        RECT 56.750 58.880 57.010 59.140 ;
        RECT 76.430 59.250 76.690 59.510 ;
        RECT 51.950 58.510 52.210 58.770 ;
        RECT 64.430 58.510 64.690 58.770 ;
        RECT 8.750 58.140 9.010 58.400 ;
        RECT 33.230 58.140 33.490 58.400 ;
        RECT 61.070 58.140 61.330 58.400 ;
        RECT 121.550 59.620 121.810 59.880 ;
        RECT 87.950 59.250 88.210 59.510 ;
        RECT 105.230 59.250 105.490 59.510 ;
        RECT 117.230 59.250 117.490 59.510 ;
        RECT 120.590 59.250 120.850 59.510 ;
        RECT 123.470 59.250 123.730 59.510 ;
        RECT 95.150 58.880 95.410 59.140 ;
        RECT 101.870 58.880 102.130 59.140 ;
        RECT 115.310 58.880 115.570 59.140 ;
        RECT 122.510 58.880 122.770 59.140 ;
        RECT 130.190 58.880 130.450 59.140 ;
        RECT 118.190 58.510 118.450 58.770 ;
        RECT 25.070 57.770 25.330 58.030 ;
        RECT 26.510 57.770 26.770 58.030 ;
        RECT 55.310 57.770 55.570 58.030 ;
        RECT 9.230 55.920 9.490 56.180 ;
        RECT 19.310 55.920 19.570 56.180 ;
        RECT 42.350 55.920 42.610 56.180 ;
        RECT 75.950 55.920 76.210 56.180 ;
        RECT 90.830 55.920 91.090 56.180 ;
        RECT 97.550 55.920 97.810 56.180 ;
        RECT 136.910 55.920 137.170 56.180 ;
        RECT 10.670 55.550 10.930 55.810 ;
        RECT 13.070 55.550 13.330 55.810 ;
        RECT 6.350 54.440 6.610 54.700 ;
        RECT 15.470 54.810 15.730 55.070 ;
        RECT 18.350 54.810 18.610 55.070 ;
        RECT 26.990 55.550 27.250 55.810 ;
        RECT 45.230 55.550 45.490 55.810 ;
        RECT 58.670 55.550 58.930 55.810 ;
        RECT 23.630 55.180 23.890 55.440 ;
        RECT 26.030 55.180 26.290 55.440 ;
        RECT 43.790 55.180 44.050 55.440 ;
        RECT 49.550 55.180 49.810 55.440 ;
        RECT 57.710 55.180 57.970 55.440 ;
        RECT 24.110 54.810 24.370 55.070 ;
        RECT 29.870 54.810 30.130 55.070 ;
        RECT 31.790 54.810 32.050 55.070 ;
        RECT 38.510 54.810 38.770 55.070 ;
        RECT 6.830 54.070 7.090 54.330 ;
        RECT 23.150 54.440 23.410 54.700 ;
        RECT 36.590 54.440 36.850 54.700 ;
        RECT 42.830 54.440 43.090 54.700 ;
        RECT 44.270 54.440 44.530 54.700 ;
        RECT 47.630 54.440 47.890 54.700 ;
        RECT 51.950 54.810 52.210 55.070 ;
        RECT 52.910 54.810 53.170 55.070 ;
        RECT 58.670 54.810 58.930 55.070 ;
        RECT 46.670 54.070 46.930 54.330 ;
        RECT 56.270 54.070 56.530 54.330 ;
        RECT 57.710 54.070 57.970 54.330 ;
        RECT 67.790 54.440 68.050 54.700 ;
        RECT 82.670 54.440 82.930 54.700 ;
        RECT 86.990 54.810 87.250 55.070 ;
        RECT 87.950 54.440 88.210 54.700 ;
        RECT 87.470 54.070 87.730 54.330 ;
        RECT 90.350 54.440 90.610 54.700 ;
        RECT 100.910 54.810 101.170 55.070 ;
        RECT 123.470 55.180 123.730 55.440 ;
        RECT 135.950 55.180 136.210 55.440 ;
        RECT 108.590 54.810 108.850 55.070 ;
        RECT 117.710 54.810 117.970 55.070 ;
        RECT 121.070 54.810 121.330 55.070 ;
        RECT 129.230 54.810 129.490 55.070 ;
        RECT 98.030 54.440 98.290 54.700 ;
        RECT 110.030 54.440 110.290 54.700 ;
        RECT 122.510 54.440 122.770 54.700 ;
        RECT 130.190 54.440 130.450 54.700 ;
        RECT 133.070 54.810 133.330 55.070 ;
        RECT 137.870 54.810 138.130 55.070 ;
        RECT 137.390 54.440 137.650 54.700 ;
        RECT 99.470 54.070 99.730 54.330 ;
        RECT 116.750 54.070 117.010 54.330 ;
        RECT 118.190 54.070 118.450 54.330 ;
        RECT 19.310 53.700 19.570 53.960 ;
        RECT 38.990 53.700 39.250 53.960 ;
        RECT 39.470 53.700 39.730 53.960 ;
        RECT 78.830 53.700 79.090 53.960 ;
        RECT 98.030 53.700 98.290 53.960 ;
        RECT 99.950 53.700 100.210 53.960 ;
        RECT 13.070 51.110 13.330 51.370 ;
        RECT 18.350 51.850 18.610 52.110 ;
        RECT 22.190 51.480 22.450 51.740 ;
        RECT 17.870 51.110 18.130 51.370 ;
        RECT 20.750 51.110 21.010 51.370 ;
        RECT 21.710 51.110 21.970 51.370 ;
        RECT 23.150 51.110 23.410 51.370 ;
        RECT 82.670 51.850 82.930 52.110 ;
        RECT 26.030 51.480 26.290 51.740 ;
        RECT 24.110 51.110 24.370 51.370 ;
        RECT 26.510 51.110 26.770 51.370 ;
        RECT 39.470 51.480 39.730 51.740 ;
        RECT 50.030 51.480 50.290 51.740 ;
        RECT 60.110 51.480 60.370 51.740 ;
        RECT 72.590 51.480 72.850 51.740 ;
        RECT 78.830 51.480 79.090 51.740 ;
        RECT 90.350 51.480 90.610 51.740 ;
        RECT 30.830 51.110 31.090 51.370 ;
        RECT 33.230 51.110 33.490 51.370 ;
        RECT 61.070 51.110 61.330 51.370 ;
        RECT 12.590 50.370 12.850 50.630 ;
        RECT 42.830 50.740 43.090 51.000 ;
        RECT 49.550 50.740 49.810 51.000 ;
        RECT 61.550 50.740 61.810 51.000 ;
        RECT 36.590 50.370 36.850 50.630 ;
        RECT 52.430 50.370 52.690 50.630 ;
        RECT 58.670 50.370 58.930 50.630 ;
        RECT 75.950 51.110 76.210 51.370 ;
        RECT 100.910 51.480 101.170 51.740 ;
        RECT 116.270 51.480 116.530 51.740 ;
        RECT 133.070 51.480 133.330 51.740 ;
        RECT 68.270 50.740 68.530 51.000 ;
        RECT 74.990 50.740 75.250 51.000 ;
        RECT 99.950 51.110 100.210 51.370 ;
        RECT 108.590 51.110 108.850 51.370 ;
        RECT 81.230 50.370 81.490 50.630 ;
        RECT 95.150 50.740 95.410 51.000 ;
        RECT 110.510 50.740 110.770 51.000 ;
        RECT 118.190 50.740 118.450 51.000 ;
        RECT 128.270 51.110 128.530 51.370 ;
        RECT 129.230 51.110 129.490 51.370 ;
        RECT 126.350 50.740 126.610 51.000 ;
        RECT 127.310 50.740 127.570 51.000 ;
        RECT 135.950 50.740 136.210 51.000 ;
        RECT 139.310 51.110 139.570 51.370 ;
        RECT 138.350 50.370 138.610 50.630 ;
        RECT 20.270 50.000 20.530 50.260 ;
        RECT 32.270 50.000 32.530 50.260 ;
        RECT 35.150 50.000 35.410 50.260 ;
        RECT 36.110 50.000 36.370 50.260 ;
        RECT 48.110 50.000 48.370 50.260 ;
        RECT 35.630 49.630 35.890 49.890 ;
        RECT 74.990 50.000 75.250 50.260 ;
        RECT 94.190 49.630 94.450 49.890 ;
        RECT 45.230 47.780 45.490 48.040 ;
        RECT 72.110 47.780 72.370 48.040 ;
        RECT 61.550 47.410 61.810 47.670 ;
        RECT 66.350 47.410 66.610 47.670 ;
        RECT 97.550 47.410 97.810 47.670 ;
        RECT 12.590 47.040 12.850 47.300 ;
        RECT 21.710 47.040 21.970 47.300 ;
        RECT 26.030 46.670 26.290 46.930 ;
        RECT 29.390 46.670 29.650 46.930 ;
        RECT 52.430 47.040 52.690 47.300 ;
        RECT 35.630 46.670 35.890 46.930 ;
        RECT 44.750 46.670 45.010 46.930 ;
        RECT 20.750 46.300 21.010 46.560 ;
        RECT 28.910 46.300 29.170 46.560 ;
        RECT 30.830 46.300 31.090 46.560 ;
        RECT 42.350 46.300 42.610 46.560 ;
        RECT 42.830 46.300 43.090 46.560 ;
        RECT 52.910 46.670 53.170 46.930 ;
        RECT 54.830 46.670 55.090 46.930 ;
        RECT 60.110 46.670 60.370 46.930 ;
        RECT 43.310 45.930 43.570 46.190 ;
        RECT 58.190 45.930 58.450 46.190 ;
        RECT 59.150 45.930 59.410 46.190 ;
        RECT 66.830 46.670 67.090 46.930 ;
        RECT 89.870 46.670 90.130 46.930 ;
        RECT 101.390 47.040 101.650 47.300 ;
        RECT 100.430 46.670 100.690 46.930 ;
        RECT 66.350 46.300 66.610 46.560 ;
        RECT 65.870 45.930 66.130 46.190 ;
        RECT 91.790 45.930 92.050 46.190 ;
        RECT 48.110 45.560 48.370 45.820 ;
        RECT 83.150 45.560 83.410 45.820 ;
        RECT 87.470 45.560 87.730 45.820 ;
        RECT 95.150 45.560 95.410 45.820 ;
        RECT 97.550 45.930 97.810 46.190 ;
        RECT 98.990 46.300 99.250 46.560 ;
        RECT 102.350 46.300 102.610 46.560 ;
        RECT 103.310 46.300 103.570 46.560 ;
        RECT 112.430 46.670 112.690 46.930 ;
        RECT 117.230 46.670 117.490 46.930 ;
        RECT 128.270 46.300 128.530 46.560 ;
        RECT 101.870 45.930 102.130 46.190 ;
        RECT 117.710 45.930 117.970 46.190 ;
        RECT 136.430 45.930 136.690 46.190 ;
        RECT 100.910 45.560 101.170 45.820 ;
        RECT 136.910 45.560 137.170 45.820 ;
        RECT 50.510 43.710 50.770 43.970 ;
        RECT 96.590 43.710 96.850 43.970 ;
        RECT 98.030 43.710 98.290 43.970 ;
        RECT 15.470 43.340 15.730 43.600 ;
        RECT 22.670 43.340 22.930 43.600 ;
        RECT 54.830 43.340 55.090 43.600 ;
        RECT 13.070 42.970 13.330 43.230 ;
        RECT 20.270 42.970 20.530 43.230 ;
        RECT 21.230 42.970 21.490 43.230 ;
        RECT 15.950 42.600 16.210 42.860 ;
        RECT 17.870 42.600 18.130 42.860 ;
        RECT 29.870 42.970 30.130 43.230 ;
        RECT 30.830 42.970 31.090 43.230 ;
        RECT 38.030 42.970 38.290 43.230 ;
        RECT 40.910 42.970 41.170 43.230 ;
        RECT 54.350 42.970 54.610 43.230 ;
        RECT 59.150 42.970 59.410 43.230 ;
        RECT 22.190 42.600 22.450 42.860 ;
        RECT 23.630 42.600 23.890 42.860 ;
        RECT 33.710 42.600 33.970 42.860 ;
        RECT 28.910 42.230 29.170 42.490 ;
        RECT 29.390 41.860 29.650 42.120 ;
        RECT 56.270 42.600 56.530 42.860 ;
        RECT 58.190 42.600 58.450 42.860 ;
        RECT 59.630 42.600 59.890 42.860 ;
        RECT 76.910 42.970 77.170 43.230 ;
        RECT 64.910 42.600 65.170 42.860 ;
        RECT 66.350 42.600 66.610 42.860 ;
        RECT 66.830 42.230 67.090 42.490 ;
        RECT 72.590 41.860 72.850 42.120 ;
        RECT 87.950 42.970 88.210 43.230 ;
        RECT 94.190 42.970 94.450 43.230 ;
        RECT 100.430 43.340 100.690 43.600 ;
        RECT 110.510 43.340 110.770 43.600 ;
        RECT 97.550 42.970 97.810 43.230 ;
        RECT 85.070 42.600 85.330 42.860 ;
        RECT 91.790 42.600 92.050 42.860 ;
        RECT 95.150 42.600 95.410 42.860 ;
        RECT 98.990 42.600 99.250 42.860 ;
        RECT 106.190 42.600 106.450 42.860 ;
        RECT 121.070 42.970 121.330 43.230 ;
        RECT 127.310 42.970 127.570 43.230 ;
        RECT 127.790 42.970 128.050 43.230 ;
        RECT 120.590 42.600 120.850 42.860 ;
        RECT 121.550 42.600 121.810 42.860 ;
        RECT 133.550 42.600 133.810 42.860 ;
        RECT 94.670 42.230 94.930 42.490 ;
        RECT 138.350 43.340 138.610 43.600 ;
        RECT 103.790 41.860 104.050 42.120 ;
        RECT 22.190 41.490 22.450 41.750 ;
        RECT 26.990 41.490 27.250 41.750 ;
        RECT 56.750 41.490 57.010 41.750 ;
        RECT 79.790 41.490 80.050 41.750 ;
        RECT 96.590 41.490 96.850 41.750 ;
        RECT 103.310 41.490 103.570 41.750 ;
        RECT 138.350 41.490 138.610 41.750 ;
        RECT 15.950 39.640 16.210 39.900 ;
        RECT 13.070 39.270 13.330 39.530 ;
        RECT 33.710 39.640 33.970 39.900 ;
        RECT 40.910 39.640 41.170 39.900 ;
        RECT 74.990 39.640 75.250 39.900 ;
        RECT 25.070 39.270 25.330 39.530 ;
        RECT 54.350 39.270 54.610 39.530 ;
        RECT 81.230 39.640 81.490 39.900 ;
        RECT 83.150 39.640 83.410 39.900 ;
        RECT 100.430 39.640 100.690 39.900 ;
        RECT 124.910 39.640 125.170 39.900 ;
        RECT 129.710 39.640 129.970 39.900 ;
        RECT 136.430 39.640 136.690 39.900 ;
        RECT 89.870 39.270 90.130 39.530 ;
        RECT 95.150 39.270 95.410 39.530 ;
        RECT 97.070 39.270 97.330 39.530 ;
        RECT 99.470 39.270 99.730 39.530 ;
        RECT 130.670 39.270 130.930 39.530 ;
        RECT 21.710 38.900 21.970 39.160 ;
        RECT 19.790 38.530 20.050 38.790 ;
        RECT 28.430 38.530 28.690 38.790 ;
        RECT 31.790 38.530 32.050 38.790 ;
        RECT 33.230 38.530 33.490 38.790 ;
        RECT 34.190 38.900 34.450 39.160 ;
        RECT 45.230 38.900 45.490 39.160 ;
        RECT 25.070 38.160 25.330 38.420 ;
        RECT 26.030 38.160 26.290 38.420 ;
        RECT 29.870 38.160 30.130 38.420 ;
        RECT 36.110 38.160 36.370 38.420 ;
        RECT 44.750 38.160 45.010 38.420 ;
        RECT 48.110 38.530 48.370 38.790 ;
        RECT 38.510 37.790 38.770 38.050 ;
        RECT 50.030 37.790 50.290 38.050 ;
        RECT 26.030 37.420 26.290 37.680 ;
        RECT 29.390 37.420 29.650 37.680 ;
        RECT 33.230 37.420 33.490 37.680 ;
        RECT 40.430 37.420 40.690 37.680 ;
        RECT 59.630 38.530 59.890 38.790 ;
        RECT 57.710 38.160 57.970 38.420 ;
        RECT 68.750 38.530 69.010 38.790 ;
        RECT 86.990 38.530 87.250 38.790 ;
        RECT 64.910 38.160 65.170 38.420 ;
        RECT 85.070 38.160 85.330 38.420 ;
        RECT 97.550 38.900 97.810 39.160 ;
        RECT 98.990 38.900 99.250 39.160 ;
        RECT 101.390 38.900 101.650 39.160 ;
        RECT 98.030 38.530 98.290 38.790 ;
        RECT 102.350 38.530 102.610 38.790 ;
        RECT 100.910 38.160 101.170 38.420 ;
        RECT 136.430 38.900 136.690 39.160 ;
        RECT 138.350 38.900 138.610 39.160 ;
        RECT 112.430 38.530 112.690 38.790 ;
        RECT 124.430 38.530 124.690 38.790 ;
        RECT 108.110 38.160 108.370 38.420 ;
        RECT 123.470 38.160 123.730 38.420 ;
        RECT 129.230 38.530 129.490 38.790 ;
        RECT 135.950 38.530 136.210 38.790 ;
        RECT 101.390 37.790 101.650 38.050 ;
        RECT 122.990 37.790 123.250 38.050 ;
        RECT 57.230 37.420 57.490 37.680 ;
        RECT 99.470 37.420 99.730 37.680 ;
        RECT 57.710 35.570 57.970 35.830 ;
        RECT 98.510 35.570 98.770 35.830 ;
        RECT 103.310 35.570 103.570 35.830 ;
        RECT 21.710 34.830 21.970 35.090 ;
        RECT 29.870 35.200 30.130 35.460 ;
        RECT 60.590 35.200 60.850 35.460 ;
        RECT 111.950 35.570 112.210 35.830 ;
        RECT 123.470 35.570 123.730 35.830 ;
        RECT 26.510 34.830 26.770 35.090 ;
        RECT 23.630 34.460 23.890 34.720 ;
        RECT 35.150 34.830 35.410 35.090 ;
        RECT 28.910 34.460 29.170 34.720 ;
        RECT 32.750 34.460 33.010 34.720 ;
        RECT 42.350 34.460 42.610 34.720 ;
        RECT 25.550 33.720 25.810 33.980 ;
        RECT 9.710 33.350 9.970 33.610 ;
        RECT 15.470 33.350 15.730 33.610 ;
        RECT 20.750 33.350 21.010 33.610 ;
        RECT 35.630 34.090 35.890 34.350 ;
        RECT 54.350 34.830 54.610 35.090 ;
        RECT 66.350 34.830 66.610 35.090 ;
        RECT 78.830 34.830 79.090 35.090 ;
        RECT 44.750 34.460 45.010 34.720 ;
        RECT 51.470 34.460 51.730 34.720 ;
        RECT 59.150 34.460 59.410 34.720 ;
        RECT 81.230 34.460 81.490 34.720 ;
        RECT 86.510 34.460 86.770 34.720 ;
        RECT 94.670 34.830 94.930 35.090 ;
        RECT 98.990 34.460 99.250 34.720 ;
        RECT 100.430 34.460 100.690 34.720 ;
        RECT 63.470 34.090 63.730 34.350 ;
        RECT 64.910 34.090 65.170 34.350 ;
        RECT 106.670 35.200 106.930 35.460 ;
        RECT 124.430 35.570 124.690 35.830 ;
        RECT 118.190 34.830 118.450 35.090 ;
        RECT 124.910 35.200 125.170 35.460 ;
        RECT 126.350 35.570 126.610 35.830 ;
        RECT 129.710 35.570 129.970 35.830 ;
        RECT 136.430 35.570 136.690 35.830 ;
        RECT 110.030 34.460 110.290 34.720 ;
        RECT 110.990 34.460 111.250 34.720 ;
        RECT 127.790 34.460 128.050 34.720 ;
        RECT 106.190 34.090 106.450 34.350 ;
        RECT 136.910 34.830 137.170 35.090 ;
        RECT 118.190 33.720 118.450 33.980 ;
        RECT 120.590 33.720 120.850 33.980 ;
        RECT 35.630 33.350 35.890 33.610 ;
        RECT 57.230 33.350 57.490 33.610 ;
        RECT 86.510 33.350 86.770 33.610 ;
        RECT 103.790 33.350 104.050 33.610 ;
        RECT 106.670 33.350 106.930 33.610 ;
        RECT 110.990 33.350 111.250 33.610 ;
        RECT 111.950 33.350 112.210 33.610 ;
        RECT 122.510 33.350 122.770 33.610 ;
        RECT 29.390 31.500 29.650 31.760 ;
        RECT 31.790 31.500 32.050 31.760 ;
        RECT 42.350 31.500 42.610 31.760 ;
        RECT 79.790 31.500 80.050 31.760 ;
        RECT 95.150 31.500 95.410 31.760 ;
        RECT 22.190 31.130 22.450 31.390 ;
        RECT 54.350 31.130 54.610 31.390 ;
        RECT 59.630 31.130 59.890 31.390 ;
        RECT 9.710 30.760 9.970 31.020 ;
        RECT 25.550 30.760 25.810 31.020 ;
        RECT 20.750 30.020 21.010 30.280 ;
        RECT 26.990 30.020 27.250 30.280 ;
        RECT 32.750 30.390 33.010 30.650 ;
        RECT 35.150 30.390 35.410 30.650 ;
        RECT 37.550 30.760 37.810 31.020 ;
        RECT 29.390 30.020 29.650 30.280 ;
        RECT 33.710 30.020 33.970 30.280 ;
        RECT 36.110 30.020 36.370 30.280 ;
        RECT 42.350 30.390 42.610 30.650 ;
        RECT 51.470 30.760 51.730 31.020 ;
        RECT 55.310 30.390 55.570 30.650 ;
        RECT 59.150 30.390 59.410 30.650 ;
        RECT 34.670 29.650 34.930 29.910 ;
        RECT 60.590 30.020 60.850 30.280 ;
        RECT 65.390 30.020 65.650 30.280 ;
        RECT 82.670 30.390 82.930 30.650 ;
        RECT 83.630 30.390 83.890 30.650 ;
        RECT 80.750 30.020 81.010 30.280 ;
        RECT 98.030 31.130 98.290 31.390 ;
        RECT 105.710 31.130 105.970 31.390 ;
        RECT 97.550 30.760 97.810 31.020 ;
        RECT 101.870 30.760 102.130 31.020 ;
        RECT 110.990 30.760 111.250 31.020 ;
        RECT 94.190 30.390 94.450 30.650 ;
        RECT 100.910 30.390 101.170 30.650 ;
        RECT 48.110 29.650 48.370 29.910 ;
        RECT 62.510 29.650 62.770 29.910 ;
        RECT 95.150 30.020 95.410 30.280 ;
        RECT 98.990 30.020 99.250 30.280 ;
        RECT 93.710 29.650 93.970 29.910 ;
        RECT 99.470 29.650 99.730 29.910 ;
        RECT 103.310 29.650 103.570 29.910 ;
        RECT 105.710 30.020 105.970 30.280 ;
        RECT 108.110 30.390 108.370 30.650 ;
        RECT 111.470 29.650 111.730 29.910 ;
        RECT 21.710 29.280 21.970 29.540 ;
        RECT 29.870 29.280 30.130 29.540 ;
        RECT 33.710 29.280 33.970 29.540 ;
        RECT 47.630 29.280 47.890 29.540 ;
        RECT 72.110 29.280 72.370 29.540 ;
        RECT 86.030 29.280 86.290 29.540 ;
        RECT 105.710 29.280 105.970 29.540 ;
        RECT 121.070 31.130 121.330 31.390 ;
        RECT 137.870 31.130 138.130 31.390 ;
        RECT 115.310 29.650 115.570 29.910 ;
        RECT 121.070 30.020 121.330 30.280 ;
        RECT 122.990 30.390 123.250 30.650 ;
        RECT 123.470 30.020 123.730 30.280 ;
        RECT 116.750 29.650 117.010 29.910 ;
        RECT 136.910 30.020 137.170 30.280 ;
        RECT 127.310 29.650 127.570 29.910 ;
        RECT 117.710 29.280 117.970 29.540 ;
        RECT 125.390 29.280 125.650 29.540 ;
        RECT 21.710 27.430 21.970 27.690 ;
        RECT 19.310 27.060 19.570 27.320 ;
        RECT 26.030 27.060 26.290 27.320 ;
        RECT 19.790 26.320 20.050 26.580 ;
        RECT 26.510 26.690 26.770 26.950 ;
        RECT 33.710 27.430 33.970 27.690 ;
        RECT 32.750 27.060 33.010 27.320 ;
        RECT 43.790 27.060 44.050 27.320 ;
        RECT 38.510 26.690 38.770 26.950 ;
        RECT 22.190 25.950 22.450 26.210 ;
        RECT 24.110 25.950 24.370 26.210 ;
        RECT 27.470 26.320 27.730 26.580 ;
        RECT 36.110 26.320 36.370 26.580 ;
        RECT 39.470 26.320 39.730 26.580 ;
        RECT 40.430 26.320 40.690 26.580 ;
        RECT 56.270 26.320 56.530 26.580 ;
        RECT 58.670 26.320 58.930 26.580 ;
        RECT 35.150 25.950 35.410 26.210 ;
        RECT 35.630 25.950 35.890 26.210 ;
        RECT 65.390 26.320 65.650 26.580 ;
        RECT 103.310 27.430 103.570 27.690 ;
        RECT 106.670 27.430 106.930 27.690 ;
        RECT 111.470 27.430 111.730 27.690 ;
        RECT 68.750 27.060 69.010 27.320 ;
        RECT 96.110 27.060 96.370 27.320 ;
        RECT 111.950 27.060 112.210 27.320 ;
        RECT 124.910 27.430 125.170 27.690 ;
        RECT 68.270 26.690 68.530 26.950 ;
        RECT 86.510 26.690 86.770 26.950 ;
        RECT 76.910 26.320 77.170 26.580 ;
        RECT 82.670 25.950 82.930 26.210 ;
        RECT 94.670 26.320 94.930 26.580 ;
        RECT 97.550 26.690 97.810 26.950 ;
        RECT 103.790 26.690 104.050 26.950 ;
        RECT 108.590 26.690 108.850 26.950 ;
        RECT 99.470 26.320 99.730 26.580 ;
        RECT 115.310 26.320 115.570 26.580 ;
        RECT 116.750 26.320 117.010 26.580 ;
        RECT 118.190 27.060 118.450 27.320 ;
        RECT 127.310 27.060 127.570 27.320 ;
        RECT 122.510 26.690 122.770 26.950 ;
        RECT 123.470 26.690 123.730 26.950 ;
        RECT 118.190 26.320 118.450 26.580 ;
        RECT 130.670 26.690 130.930 26.950 ;
        RECT 93.710 25.950 93.970 26.210 ;
        RECT 19.790 25.580 20.050 25.840 ;
        RECT 20.270 25.210 20.530 25.470 ;
        RECT 64.910 25.580 65.170 25.840 ;
        RECT 110.030 25.580 110.290 25.840 ;
        RECT 34.670 25.210 34.930 25.470 ;
        RECT 86.990 25.210 87.250 25.470 ;
        RECT 129.230 25.210 129.490 25.470 ;
        RECT 20.270 23.360 20.530 23.620 ;
        RECT 67.310 23.360 67.570 23.620 ;
        RECT 78.830 23.360 79.090 23.620 ;
        RECT 86.990 23.360 87.250 23.620 ;
        RECT 94.190 23.360 94.450 23.620 ;
        RECT 117.710 23.360 117.970 23.620 ;
        RECT 136.910 23.360 137.170 23.620 ;
        RECT 35.150 22.990 35.410 23.250 ;
        RECT 42.830 22.990 43.090 23.250 ;
        RECT 64.910 22.990 65.170 23.250 ;
        RECT 66.830 22.990 67.090 23.250 ;
        RECT 81.230 22.990 81.490 23.250 ;
        RECT 87.470 22.990 87.730 23.250 ;
        RECT 103.790 22.990 104.050 23.250 ;
        RECT 52.910 22.620 53.170 22.880 ;
        RECT 67.790 22.620 68.050 22.880 ;
        RECT 97.550 22.620 97.810 22.880 ;
        RECT 94.670 22.250 94.930 22.510 ;
        RECT 130.670 22.990 130.930 23.250 ;
        RECT 115.310 22.620 115.570 22.880 ;
        RECT 129.230 22.620 129.490 22.880 ;
        RECT 29.390 21.880 29.650 22.140 ;
        RECT 47.630 21.880 47.890 22.140 ;
        RECT 72.110 21.880 72.370 22.140 ;
        RECT 96.110 21.880 96.370 22.140 ;
        RECT 101.390 21.880 101.650 22.140 ;
        RECT 103.790 21.880 104.050 22.140 ;
        RECT 99.950 21.510 100.210 21.770 ;
        RECT 100.910 21.510 101.170 21.770 ;
        RECT 116.750 22.250 117.010 22.510 ;
        RECT 118.190 22.250 118.450 22.510 ;
        RECT 120.590 22.250 120.850 22.510 ;
        RECT 125.390 21.880 125.650 22.140 ;
        RECT 33.230 21.140 33.490 21.400 ;
        RECT 53.390 21.140 53.650 21.400 ;
        RECT 66.830 21.140 67.090 21.400 ;
        RECT 69.710 21.140 69.970 21.400 ;
        RECT 83.630 21.140 83.890 21.400 ;
        RECT 94.190 21.140 94.450 21.400 ;
        RECT 105.230 21.510 105.490 21.770 ;
        RECT 109.070 21.140 109.330 21.400 ;
        RECT 53.390 19.290 53.650 19.550 ;
        RECT 56.270 19.290 56.530 19.550 ;
        RECT 65.870 19.290 66.130 19.550 ;
        RECT 66.350 19.290 66.610 19.550 ;
        RECT 72.590 19.290 72.850 19.550 ;
        RECT 76.430 19.290 76.690 19.550 ;
        RECT 86.030 19.290 86.290 19.550 ;
        RECT 97.550 19.290 97.810 19.550 ;
        RECT 105.710 19.290 105.970 19.550 ;
        RECT 118.190 19.290 118.450 19.550 ;
        RECT 64.430 18.920 64.690 19.180 ;
        RECT 94.190 18.920 94.450 19.180 ;
        RECT 109.070 18.920 109.330 19.180 ;
        RECT 33.230 18.180 33.490 18.440 ;
        RECT 37.550 18.180 37.810 18.440 ;
        RECT 57.230 18.550 57.490 18.810 ;
        RECT 59.630 18.550 59.890 18.810 ;
        RECT 65.870 18.550 66.130 18.810 ;
        RECT 67.310 18.550 67.570 18.810 ;
        RECT 77.870 18.550 78.130 18.810 ;
        RECT 39.470 18.180 39.730 18.440 ;
        RECT 15.470 17.440 15.730 17.700 ;
        RECT 42.830 17.440 43.090 17.700 ;
        RECT 24.110 17.070 24.370 17.330 ;
        RECT 41.870 17.070 42.130 17.330 ;
        RECT 45.230 17.810 45.490 18.070 ;
        RECT 51.470 18.180 51.730 18.440 ;
        RECT 52.910 18.180 53.170 18.440 ;
        RECT 63.470 18.180 63.730 18.440 ;
        RECT 68.750 18.180 69.010 18.440 ;
        RECT 69.710 18.180 69.970 18.440 ;
        RECT 45.710 17.440 45.970 17.700 ;
        RECT 64.430 17.440 64.690 17.700 ;
        RECT 66.830 17.440 67.090 17.700 ;
        RECT 106.190 17.440 106.450 17.700 ;
        RECT 53.870 17.070 54.130 17.330 ;
        RECT 41.870 15.590 42.130 15.850 ;
        RECT 64.430 15.590 64.690 15.850 ;
      LAYER met2 ;
        RECT 117.230 144.690 117.490 145.010 ;
        RECT 32.750 143.950 33.010 144.270 ;
        RECT 49.550 143.950 49.810 144.270 ;
        RECT 77.870 143.950 78.130 144.270 ;
        RECT 99.470 143.950 99.730 144.270 ;
        RECT 30.830 143.210 31.090 143.530 ;
        RECT 30.890 136.870 31.030 143.210 ;
        RECT 30.830 136.550 31.090 136.870 ;
        RECT 32.810 133.540 32.950 143.950 ;
        RECT 36.590 143.210 36.850 143.530 ;
        RECT 36.650 141.680 36.790 143.210 ;
        RECT 36.590 141.360 36.850 141.680 ;
        RECT 33.710 140.620 33.970 140.940 ;
        RECT 44.270 140.620 44.530 140.940 ;
        RECT 32.750 133.220 33.010 133.540 ;
        RECT 29.390 132.480 29.650 132.800 ;
        RECT 16.910 127.670 17.170 127.990 ;
        RECT 15.470 126.930 15.730 127.250 ;
        RECT 15.530 125.400 15.670 126.930 ;
        RECT 15.470 125.080 15.730 125.400 ;
        RECT 16.970 120.590 17.110 127.670 ;
        RECT 26.030 127.300 26.290 127.620 ;
        RECT 20.270 124.340 20.530 124.660 ;
        RECT 20.330 121.330 20.470 124.340 ;
        RECT 25.070 122.860 25.330 123.180 ;
        RECT 20.270 121.010 20.530 121.330 ;
        RECT 16.910 120.270 17.170 120.590 ;
        RECT 16.970 116.520 17.110 120.270 ;
        RECT 25.130 119.850 25.270 122.860 ;
        RECT 25.070 119.530 25.330 119.850 ;
        RECT 25.550 119.160 25.810 119.480 ;
        RECT 23.150 118.790 23.410 119.110 ;
        RECT 23.210 116.520 23.350 118.790 ;
        RECT 16.910 116.200 17.170 116.520 ;
        RECT 23.150 116.200 23.410 116.520 ;
        RECT 25.070 116.200 25.330 116.520 ;
        RECT 14.030 114.720 14.290 115.040 ;
        RECT 14.090 112.450 14.230 114.720 ;
        RECT 25.130 113.190 25.270 116.200 ;
        RECT 25.070 112.870 25.330 113.190 ;
        RECT 14.030 112.130 14.290 112.450 ;
        RECT 25.610 111.990 25.750 119.160 ;
        RECT 25.130 111.850 25.750 111.990 ;
        RECT 25.130 111.710 25.270 111.850 ;
        RECT 25.070 111.390 25.330 111.710 ;
        RECT 25.130 109.220 25.270 111.390 ;
        RECT 24.170 109.080 25.270 109.220 ;
        RECT 24.170 108.380 24.310 109.080 ;
        RECT 23.150 108.060 23.410 108.380 ;
        RECT 24.110 108.060 24.370 108.380 ;
        RECT 13.070 106.580 13.330 106.900 ;
        RECT 13.130 103.570 13.270 106.580 ;
        RECT 13.070 103.250 13.330 103.570 ;
        RECT 21.230 102.880 21.490 103.200 ;
        RECT 21.290 100.980 21.430 102.880 ;
        RECT 21.230 100.660 21.490 100.980 ;
        RECT 22.190 99.920 22.450 100.240 ;
        RECT 14.510 98.440 14.770 98.760 ;
        RECT 8.750 94.370 9.010 94.690 ;
        RECT 8.810 92.840 8.950 94.370 ;
        RECT 8.750 92.520 9.010 92.840 ;
        RECT 14.570 90.620 14.710 98.440 ;
        RECT 22.250 96.910 22.390 99.920 ;
        RECT 23.210 98.760 23.350 108.060 ;
        RECT 23.150 98.440 23.410 98.760 ;
        RECT 22.190 96.590 22.450 96.910 ;
        RECT 23.210 96.170 23.350 98.440 ;
        RECT 23.150 95.850 23.410 96.170 ;
        RECT 24.170 95.800 24.310 108.060 ;
        RECT 26.090 95.900 26.230 127.300 ;
        RECT 29.450 120.320 29.590 132.480 ;
        RECT 33.770 129.470 33.910 140.620 ;
        RECT 36.110 135.070 36.370 135.390 ;
        RECT 36.170 132.430 36.310 135.070 ;
        RECT 39.470 132.480 39.730 132.800 ;
        RECT 36.110 132.110 36.370 132.430 ;
        RECT 36.590 131.740 36.850 132.060 ;
        RECT 36.650 129.470 36.790 131.740 ;
        RECT 33.710 129.150 33.970 129.470 ;
        RECT 36.590 129.150 36.850 129.470 ;
        RECT 36.650 128.730 36.790 129.150 ;
        RECT 36.590 128.410 36.850 128.730 ;
        RECT 39.530 127.990 39.670 132.480 ;
        RECT 42.830 128.410 43.090 128.730 ;
        RECT 39.470 127.670 39.730 127.990 ;
        RECT 31.790 126.930 32.050 127.250 ;
        RECT 29.870 124.340 30.130 124.660 ;
        RECT 29.930 121.330 30.070 124.340 ;
        RECT 29.870 121.010 30.130 121.330 ;
        RECT 26.990 119.900 27.250 120.220 ;
        RECT 29.450 120.180 30.070 120.320 ;
        RECT 27.050 112.080 27.190 119.900 ;
        RECT 29.390 116.200 29.650 116.520 ;
        RECT 29.450 112.080 29.590 116.200 ;
        RECT 26.510 111.760 26.770 112.080 ;
        RECT 26.990 111.760 27.250 112.080 ;
        RECT 29.390 111.760 29.650 112.080 ;
        RECT 26.570 108.010 26.710 111.760 ;
        RECT 27.050 108.380 27.190 111.760 ;
        RECT 26.990 108.060 27.250 108.380 ;
        RECT 26.510 107.690 26.770 108.010 ;
        RECT 26.570 105.050 26.710 107.690 ;
        RECT 26.510 104.730 26.770 105.050 ;
        RECT 24.110 95.480 24.370 95.800 ;
        RECT 25.610 95.760 26.230 95.900 ;
        RECT 27.050 95.800 27.190 108.060 ;
        RECT 25.610 95.430 25.750 95.760 ;
        RECT 26.990 95.480 27.250 95.800 ;
        RECT 25.550 95.110 25.810 95.430 ;
        RECT 21.710 92.520 21.970 92.840 ;
        RECT 14.510 90.300 14.770 90.620 ;
        RECT 14.570 79.150 14.710 90.300 ;
        RECT 21.770 84.700 21.910 92.520 ;
        RECT 25.610 92.470 25.750 95.110 ;
        RECT 25.550 92.150 25.810 92.470 ;
        RECT 24.110 91.780 24.370 92.100 ;
        RECT 24.170 84.700 24.310 91.780 ;
        RECT 27.050 91.730 27.190 95.480 ;
        RECT 28.430 95.110 28.690 95.430 ;
        RECT 28.490 92.100 28.630 95.110 ;
        RECT 28.430 91.780 28.690 92.100 ;
        RECT 26.990 91.410 27.250 91.730 ;
        RECT 27.050 88.770 27.190 91.410 ;
        RECT 28.490 90.990 28.630 91.780 ;
        RECT 29.390 91.040 29.650 91.360 ;
        RECT 28.430 90.670 28.690 90.990 ;
        RECT 26.990 88.450 27.250 88.770 ;
        RECT 29.450 88.400 29.590 91.040 ;
        RECT 29.390 88.080 29.650 88.400 ;
        RECT 29.390 87.340 29.650 87.660 ;
        RECT 26.030 86.230 26.290 86.550 ;
        RECT 21.710 84.380 21.970 84.700 ;
        RECT 24.110 84.380 24.370 84.700 ;
        RECT 19.310 84.010 19.570 84.330 ;
        RECT 19.790 84.010 20.050 84.330 ;
        RECT 19.370 80.630 19.510 84.010 ;
        RECT 19.310 80.310 19.570 80.630 ;
        RECT 14.510 78.830 14.770 79.150 ;
        RECT 19.850 72.490 19.990 84.010 ;
        RECT 22.670 78.830 22.930 79.150 ;
        RECT 21.710 78.090 21.970 78.410 ;
        RECT 21.770 76.560 21.910 78.090 ;
        RECT 21.710 76.240 21.970 76.560 ;
        RECT 22.730 74.340 22.870 78.830 ;
        RECT 22.670 74.020 22.930 74.340 ;
        RECT 10.670 72.170 10.930 72.490 ;
        RECT 19.790 72.170 20.050 72.490 ;
        RECT 10.730 67.680 10.870 72.170 ;
        RECT 21.710 70.320 21.970 70.640 ;
        RECT 19.310 69.950 19.570 70.270 ;
        RECT 19.370 68.420 19.510 69.950 ;
        RECT 21.220 69.740 21.500 70.110 ;
        RECT 19.310 68.100 19.570 68.420 ;
        RECT 21.290 68.050 21.430 69.740 ;
        RECT 21.230 67.730 21.490 68.050 ;
        RECT 10.670 67.360 10.930 67.680 ;
        RECT 15.470 67.360 15.730 67.680 ;
        RECT 18.830 67.360 19.090 67.680 ;
        RECT 6.350 63.290 6.610 63.610 ;
        RECT 6.410 54.730 6.550 63.290 ;
        RECT 8.750 62.920 9.010 63.240 ;
        RECT 9.230 62.920 9.490 63.240 ;
        RECT 8.810 58.430 8.950 62.920 ;
        RECT 9.290 58.800 9.430 62.920 ;
        RECT 9.230 58.480 9.490 58.800 ;
        RECT 8.750 58.110 9.010 58.430 ;
        RECT 9.290 56.210 9.430 58.480 ;
        RECT 9.230 55.890 9.490 56.210 ;
        RECT 10.730 55.840 10.870 67.360 ;
        RECT 13.070 63.290 13.330 63.610 ;
        RECT 13.130 63.150 13.270 63.290 ;
        RECT 13.130 63.010 14.710 63.150 ;
        RECT 14.030 62.710 14.290 62.870 ;
        RECT 14.020 62.340 14.300 62.710 ;
        RECT 14.570 62.500 14.710 63.010 ;
        RECT 14.510 62.180 14.770 62.500 ;
        RECT 10.670 55.520 10.930 55.840 ;
        RECT 13.070 55.520 13.330 55.840 ;
        RECT 6.350 54.410 6.610 54.730 ;
        RECT 6.820 54.200 7.100 54.570 ;
        RECT 6.830 54.040 7.090 54.200 ;
        RECT 13.130 51.400 13.270 55.520 ;
        RECT 15.530 55.100 15.670 67.360 ;
        RECT 17.390 62.550 17.650 62.870 ;
        RECT 17.450 59.910 17.590 62.550 ;
        RECT 18.890 62.130 19.030 67.360 ;
        RECT 19.310 66.250 19.570 66.570 ;
        RECT 19.370 63.610 19.510 66.250 ;
        RECT 21.770 66.200 21.910 70.320 ;
        RECT 21.710 65.880 21.970 66.200 ;
        RECT 19.310 63.290 19.570 63.610 ;
        RECT 18.830 61.810 19.090 62.130 ;
        RECT 17.390 59.590 17.650 59.910 ;
        RECT 15.470 54.780 15.730 55.100 ;
        RECT 18.350 54.780 18.610 55.100 ;
        RECT 18.410 52.140 18.550 54.780 ;
        RECT 18.890 53.900 19.030 61.810 ;
        RECT 19.310 59.590 19.570 59.910 ;
        RECT 19.370 56.210 19.510 59.590 ;
        RECT 19.310 55.890 19.570 56.210 ;
        RECT 19.310 53.900 19.570 53.990 ;
        RECT 18.890 53.760 19.570 53.900 ;
        RECT 19.310 53.670 19.570 53.760 ;
        RECT 18.350 51.820 18.610 52.140 ;
        RECT 13.070 51.080 13.330 51.400 ;
        RECT 17.870 51.080 18.130 51.400 ;
        RECT 12.590 50.340 12.850 50.660 ;
        RECT 12.650 47.330 12.790 50.340 ;
        RECT 12.590 47.010 12.850 47.330 ;
        RECT 15.470 43.310 15.730 43.630 ;
        RECT 13.070 42.940 13.330 43.260 ;
        RECT 13.130 39.560 13.270 42.940 ;
        RECT 13.070 39.240 13.330 39.560 ;
        RECT 15.530 33.640 15.670 43.310 ;
        RECT 17.930 42.890 18.070 51.080 ;
        RECT 15.950 42.570 16.210 42.890 ;
        RECT 17.870 42.570 18.130 42.890 ;
        RECT 16.010 39.930 16.150 42.570 ;
        RECT 15.950 39.610 16.210 39.930 ;
        RECT 9.710 33.320 9.970 33.640 ;
        RECT 15.470 33.320 15.730 33.640 ;
        RECT 9.770 31.050 9.910 33.320 ;
        RECT 9.710 30.730 9.970 31.050 ;
        RECT 15.530 17.730 15.670 33.320 ;
        RECT 19.370 27.350 19.510 53.670 ;
        RECT 22.190 51.450 22.450 51.770 ;
        RECT 20.750 51.080 21.010 51.400 ;
        RECT 21.710 51.080 21.970 51.400 ;
        RECT 20.270 49.970 20.530 50.290 ;
        RECT 20.330 43.260 20.470 49.970 ;
        RECT 20.810 46.590 20.950 51.080 ;
        RECT 21.770 50.870 21.910 51.080 ;
        RECT 21.700 50.500 21.980 50.870 ;
        RECT 21.710 47.010 21.970 47.330 ;
        RECT 20.750 46.270 21.010 46.590 ;
        RECT 20.270 42.940 20.530 43.260 ;
        RECT 21.230 42.940 21.490 43.260 ;
        RECT 21.290 42.730 21.430 42.940 ;
        RECT 21.220 42.360 21.500 42.730 ;
        RECT 21.770 39.190 21.910 47.010 ;
        RECT 22.250 42.890 22.390 51.450 ;
        RECT 22.730 43.630 22.870 74.020 ;
        RECT 26.090 67.310 26.230 86.230 ;
        RECT 29.450 80.630 29.590 87.340 ;
        RECT 29.930 83.960 30.070 120.180 ;
        RECT 31.850 119.850 31.990 126.930 ;
        RECT 38.030 124.710 38.290 125.030 ;
        RECT 38.090 121.330 38.230 124.710 ;
        RECT 41.390 124.340 41.650 124.660 ;
        RECT 41.450 123.180 41.590 124.340 ;
        RECT 42.890 124.290 43.030 128.410 ;
        RECT 44.330 125.400 44.470 140.620 ;
        RECT 49.610 136.500 49.750 143.950 ;
        RECT 64.910 143.580 65.170 143.900 ;
        RECT 50.030 143.210 50.290 143.530 ;
        RECT 50.090 141.680 50.230 143.210 ;
        RECT 64.970 141.680 65.110 143.580 ;
        RECT 70.670 143.210 70.930 143.530 ;
        RECT 50.030 141.360 50.290 141.680 ;
        RECT 64.910 141.360 65.170 141.680 ;
        RECT 66.350 139.140 66.610 139.460 ;
        RECT 66.410 137.610 66.550 139.140 ;
        RECT 66.350 137.290 66.610 137.610 ;
        RECT 49.550 136.180 49.810 136.500 ;
        RECT 47.630 127.300 47.890 127.620 ;
        RECT 44.270 125.080 44.530 125.400 ;
        RECT 47.690 124.660 47.830 127.300 ;
        RECT 47.630 124.340 47.890 124.660 ;
        RECT 42.830 123.970 43.090 124.290 ;
        RECT 41.390 122.860 41.650 123.180 ;
        RECT 38.030 121.010 38.290 121.330 ;
        RECT 33.710 120.640 33.970 120.960 ;
        RECT 31.790 119.530 32.050 119.850 ;
        RECT 31.790 108.060 32.050 108.380 ;
        RECT 32.270 108.060 32.530 108.380 ;
        RECT 31.850 100.610 31.990 108.060 ;
        RECT 32.330 105.050 32.470 108.060 ;
        RECT 32.270 104.730 32.530 105.050 ;
        RECT 31.790 100.290 32.050 100.610 ;
        RECT 33.770 100.240 33.910 120.640 ;
        RECT 40.910 120.270 41.170 120.590 ;
        RECT 37.550 115.460 37.810 115.780 ;
        RECT 37.610 110.970 37.750 115.460 ;
        RECT 37.550 110.650 37.810 110.970 ;
        RECT 37.610 105.050 37.750 110.650 ;
        RECT 37.550 104.730 37.810 105.050 ;
        RECT 40.970 103.570 41.110 120.270 ;
        RECT 41.450 120.220 41.590 122.860 ;
        RECT 41.390 119.900 41.650 120.220 ;
        RECT 42.890 115.780 43.030 123.970 ;
        RECT 47.690 116.890 47.830 124.340 ;
        RECT 49.610 121.330 49.750 136.180 ;
        RECT 58.190 126.930 58.450 127.250 ;
        RECT 58.250 125.400 58.390 126.930 ;
        RECT 58.190 125.080 58.450 125.400 ;
        RECT 57.710 122.860 57.970 123.180 ;
        RECT 49.550 121.010 49.810 121.330 ;
        RECT 57.770 120.960 57.910 122.860 ;
        RECT 57.710 120.640 57.970 120.960 ;
        RECT 47.630 116.570 47.890 116.890 ;
        RECT 52.430 116.570 52.690 116.890 ;
        RECT 43.790 116.200 44.050 116.520 ;
        RECT 42.830 115.460 43.090 115.780 ;
        RECT 43.850 103.940 43.990 116.200 ;
        RECT 52.490 112.080 52.630 116.570 ;
        RECT 57.770 116.150 57.910 120.640 ;
        RECT 62.510 119.530 62.770 119.850 ;
        RECT 60.590 118.790 60.850 119.110 ;
        RECT 60.650 117.260 60.790 118.790 ;
        RECT 60.590 116.940 60.850 117.260 ;
        RECT 61.550 116.200 61.810 116.520 ;
        RECT 56.750 115.830 57.010 116.150 ;
        RECT 57.710 115.830 57.970 116.150 ;
        RECT 52.910 115.090 53.170 115.410 ;
        RECT 52.430 111.760 52.690 112.080 ;
        RECT 44.750 111.020 45.010 111.340 ;
        RECT 44.810 103.940 44.950 111.020 ;
        RECT 52.430 110.650 52.690 110.970 ;
        RECT 52.490 103.940 52.630 110.650 ;
        RECT 52.970 109.120 53.110 115.090 ;
        RECT 52.910 108.800 53.170 109.120 ;
        RECT 55.310 106.580 55.570 106.900 ;
        RECT 43.790 103.620 44.050 103.940 ;
        RECT 44.750 103.620 45.010 103.940 ;
        RECT 52.430 103.620 52.690 103.940 ;
        RECT 40.910 103.250 41.170 103.570 ;
        RECT 43.310 100.290 43.570 100.610 ;
        RECT 33.710 99.920 33.970 100.240 ;
        RECT 30.350 98.440 30.610 98.760 ;
        RECT 30.410 96.540 30.550 98.440 ;
        RECT 33.770 96.910 33.910 99.920 ;
        RECT 33.710 96.590 33.970 96.910 ;
        RECT 30.350 96.220 30.610 96.540 ;
        RECT 43.370 95.800 43.510 100.290 ;
        RECT 43.850 96.910 43.990 103.620 ;
        RECT 52.490 100.890 52.630 103.620 ;
        RECT 54.350 103.250 54.610 103.570 ;
        RECT 52.490 100.750 53.110 100.890 ;
        RECT 52.430 99.920 52.690 100.240 ;
        RECT 43.790 96.590 44.050 96.910 ;
        RECT 52.490 95.800 52.630 99.920 ;
        RECT 52.970 95.800 53.110 100.750 ;
        RECT 53.870 100.290 54.130 100.610 ;
        RECT 43.310 95.480 43.570 95.800 ;
        RECT 52.430 95.480 52.690 95.800 ;
        RECT 52.910 95.480 53.170 95.800 ;
        RECT 36.590 95.110 36.850 95.430 ;
        RECT 36.110 94.370 36.370 94.690 ;
        RECT 36.170 92.840 36.310 94.370 ;
        RECT 36.110 92.520 36.370 92.840 ;
        RECT 36.650 92.200 36.790 95.110 ;
        RECT 52.910 94.740 53.170 95.060 ;
        RECT 36.170 92.060 36.790 92.200 ;
        RECT 35.150 91.040 35.410 91.360 ;
        RECT 34.670 90.300 34.930 90.620 ;
        RECT 33.710 87.710 33.970 88.030 ;
        RECT 31.790 86.970 32.050 87.290 ;
        RECT 29.870 83.640 30.130 83.960 ;
        RECT 31.850 83.590 31.990 86.970 ;
        RECT 32.270 84.010 32.530 84.330 ;
        RECT 31.790 83.270 32.050 83.590 ;
        RECT 31.310 82.530 31.570 82.850 ;
        RECT 30.830 82.160 31.090 82.480 ;
        RECT 29.390 80.310 29.650 80.630 ;
        RECT 30.890 79.150 31.030 82.160 ;
        RECT 31.370 79.150 31.510 82.530 ;
        RECT 30.830 78.830 31.090 79.150 ;
        RECT 31.310 78.830 31.570 79.150 ;
        RECT 31.790 75.870 32.050 76.190 ;
        RECT 29.390 75.130 29.650 75.450 ;
        RECT 26.510 70.690 26.770 71.010 ;
        RECT 26.030 66.990 26.290 67.310 ;
        RECT 26.570 63.980 26.710 70.690 ;
        RECT 26.990 67.360 27.250 67.680 ;
        RECT 26.510 63.660 26.770 63.980 ;
        RECT 23.150 62.920 23.410 63.240 ;
        RECT 23.210 55.010 23.350 62.920 ;
        RECT 23.630 59.960 23.890 60.280 ;
        RECT 23.690 55.470 23.830 59.960 ;
        RECT 25.070 57.740 25.330 58.060 ;
        RECT 26.510 57.740 26.770 58.060 ;
        RECT 23.630 55.150 23.890 55.470 ;
        RECT 24.110 55.010 24.370 55.100 ;
        RECT 23.210 54.870 24.370 55.010 ;
        RECT 24.110 54.780 24.370 54.870 ;
        RECT 23.150 54.570 23.410 54.730 ;
        RECT 23.140 54.200 23.420 54.570 ;
        RECT 23.150 51.310 23.410 51.400 ;
        RECT 24.110 51.310 24.370 51.400 ;
        RECT 23.150 51.170 24.370 51.310 ;
        RECT 23.150 51.080 23.410 51.170 ;
        RECT 24.110 51.080 24.370 51.170 ;
        RECT 22.670 43.310 22.930 43.630 ;
        RECT 22.190 42.570 22.450 42.890 ;
        RECT 23.630 42.570 23.890 42.890 ;
        RECT 25.130 42.730 25.270 57.740 ;
        RECT 26.030 55.150 26.290 55.470 ;
        RECT 26.090 51.770 26.230 55.150 ;
        RECT 26.030 51.450 26.290 51.770 ;
        RECT 26.570 51.400 26.710 57.740 ;
        RECT 27.050 55.840 27.190 67.360 ;
        RECT 29.450 60.280 29.590 75.130 ;
        RECT 29.870 71.430 30.130 71.750 ;
        RECT 29.930 62.870 30.070 71.430 ;
        RECT 30.350 71.060 30.610 71.380 ;
        RECT 29.870 62.550 30.130 62.870 ;
        RECT 29.390 59.960 29.650 60.280 ;
        RECT 29.870 59.220 30.130 59.540 ;
        RECT 26.990 55.520 27.250 55.840 ;
        RECT 29.930 55.100 30.070 59.220 ;
        RECT 30.410 58.800 30.550 71.060 ;
        RECT 30.830 70.320 31.090 70.640 ;
        RECT 31.310 70.320 31.570 70.640 ;
        RECT 30.350 58.480 30.610 58.800 ;
        RECT 29.870 54.780 30.130 55.100 ;
        RECT 30.890 51.400 31.030 70.320 ;
        RECT 31.370 70.110 31.510 70.320 ;
        RECT 31.300 69.740 31.580 70.110 ;
        RECT 31.850 55.100 31.990 75.870 ;
        RECT 31.790 54.780 32.050 55.100 ;
        RECT 26.510 51.080 26.770 51.400 ;
        RECT 30.830 51.080 31.090 51.400 ;
        RECT 32.330 50.290 32.470 84.010 ;
        RECT 33.770 83.320 33.910 87.710 ;
        RECT 34.730 86.920 34.870 90.300 ;
        RECT 35.210 86.920 35.350 91.040 ;
        RECT 34.670 86.600 34.930 86.920 ;
        RECT 35.150 86.600 35.410 86.920 ;
        RECT 34.730 83.960 34.870 86.600 ;
        RECT 34.670 83.640 34.930 83.960 ;
        RECT 35.210 83.590 35.350 86.600 ;
        RECT 33.770 83.180 34.390 83.320 ;
        RECT 35.150 83.270 35.410 83.590 ;
        RECT 32.750 70.690 33.010 71.010 ;
        RECT 32.810 67.310 32.950 70.690 ;
        RECT 32.750 66.990 33.010 67.310 ;
        RECT 33.230 58.110 33.490 58.430 ;
        RECT 33.290 51.400 33.430 58.110 ;
        RECT 33.230 51.080 33.490 51.400 ;
        RECT 32.270 49.970 32.530 50.290 ;
        RECT 26.030 46.640 26.290 46.960 ;
        RECT 29.390 46.640 29.650 46.960 ;
        RECT 22.190 41.460 22.450 41.780 ;
        RECT 22.250 39.770 22.390 41.460 ;
        RECT 22.180 39.400 22.460 39.770 ;
        RECT 21.710 38.870 21.970 39.190 ;
        RECT 19.790 38.500 20.050 38.820 ;
        RECT 19.310 27.030 19.570 27.350 ;
        RECT 19.850 26.610 19.990 38.500 ;
        RECT 21.710 34.800 21.970 35.120 ;
        RECT 20.750 33.320 21.010 33.640 ;
        RECT 20.810 30.310 20.950 33.320 ;
        RECT 20.750 29.990 21.010 30.310 ;
        RECT 21.770 29.570 21.910 34.800 ;
        RECT 23.690 34.750 23.830 42.570 ;
        RECT 25.060 42.360 25.340 42.730 ;
        RECT 24.100 39.400 24.380 39.770 ;
        RECT 23.630 34.430 23.890 34.750 ;
        RECT 22.190 31.100 22.450 31.420 ;
        RECT 21.710 29.250 21.970 29.570 ;
        RECT 21.770 27.720 21.910 29.250 ;
        RECT 21.710 27.400 21.970 27.720 ;
        RECT 19.790 26.290 20.050 26.610 ;
        RECT 19.850 25.870 19.990 26.290 ;
        RECT 22.250 26.240 22.390 31.100 ;
        RECT 24.170 26.240 24.310 39.400 ;
        RECT 25.070 39.240 25.330 39.560 ;
        RECT 25.130 38.450 25.270 39.240 ;
        RECT 26.090 38.450 26.230 46.640 ;
        RECT 28.910 46.270 29.170 46.590 ;
        RECT 28.970 42.520 29.110 46.270 ;
        RECT 28.910 42.200 29.170 42.520 ;
        RECT 29.450 42.150 29.590 46.640 ;
        RECT 30.830 46.270 31.090 46.590 ;
        RECT 30.890 43.260 31.030 46.270 ;
        RECT 29.870 42.940 30.130 43.260 ;
        RECT 30.830 42.940 31.090 43.260 ;
        RECT 29.390 41.830 29.650 42.150 ;
        RECT 26.990 41.460 27.250 41.780 ;
        RECT 25.070 38.130 25.330 38.450 ;
        RECT 26.030 38.130 26.290 38.450 ;
        RECT 26.090 37.710 26.230 38.130 ;
        RECT 26.030 37.390 26.290 37.710 ;
        RECT 25.550 33.690 25.810 34.010 ;
        RECT 25.610 31.050 25.750 33.690 ;
        RECT 25.550 30.730 25.810 31.050 ;
        RECT 26.090 27.350 26.230 37.390 ;
        RECT 26.510 34.800 26.770 35.120 ;
        RECT 26.030 27.030 26.290 27.350 ;
        RECT 26.570 26.980 26.710 34.800 ;
        RECT 27.050 30.310 27.190 41.460 ;
        RECT 29.450 38.920 29.590 41.830 ;
        RECT 28.490 38.820 29.590 38.920 ;
        RECT 28.430 38.780 29.590 38.820 ;
        RECT 28.430 38.500 28.690 38.780 ;
        RECT 28.970 34.750 29.110 38.780 ;
        RECT 29.930 38.450 30.070 42.940 ;
        RECT 33.710 42.570 33.970 42.890 ;
        RECT 33.770 39.930 33.910 42.570 ;
        RECT 33.710 39.610 33.970 39.930 ;
        RECT 31.790 38.500 32.050 38.820 ;
        RECT 33.230 38.500 33.490 38.820 ;
        RECT 29.870 38.130 30.130 38.450 ;
        RECT 29.390 37.390 29.650 37.710 ;
        RECT 28.910 34.430 29.170 34.750 ;
        RECT 29.450 31.790 29.590 37.390 ;
        RECT 29.870 35.170 30.130 35.490 ;
        RECT 29.390 31.470 29.650 31.790 ;
        RECT 26.990 29.990 27.250 30.310 ;
        RECT 29.390 29.990 29.650 30.310 ;
        RECT 26.510 26.660 26.770 26.980 ;
        RECT 27.050 26.520 27.190 29.990 ;
        RECT 27.470 26.520 27.730 26.610 ;
        RECT 27.050 26.380 27.730 26.520 ;
        RECT 27.470 26.290 27.730 26.380 ;
        RECT 22.190 25.920 22.450 26.240 ;
        RECT 24.110 25.920 24.370 26.240 ;
        RECT 19.790 25.550 20.050 25.870 ;
        RECT 20.270 25.180 20.530 25.500 ;
        RECT 20.330 23.650 20.470 25.180 ;
        RECT 20.270 23.330 20.530 23.650 ;
        RECT 15.470 17.410 15.730 17.730 ;
        RECT 24.170 17.360 24.310 25.920 ;
        RECT 29.450 22.170 29.590 29.990 ;
        RECT 29.930 29.570 30.070 35.170 ;
        RECT 31.850 31.790 31.990 38.500 ;
        RECT 33.290 37.710 33.430 38.500 ;
        RECT 33.230 37.390 33.490 37.710 ;
        RECT 32.750 34.430 33.010 34.750 ;
        RECT 31.790 31.470 32.050 31.790 ;
        RECT 32.810 30.680 32.950 34.430 ;
        RECT 32.750 30.360 33.010 30.680 ;
        RECT 29.870 29.250 30.130 29.570 ;
        RECT 32.810 27.350 32.950 30.360 ;
        RECT 33.770 30.310 33.910 39.610 ;
        RECT 34.250 39.190 34.390 83.180 ;
        RECT 36.170 82.480 36.310 92.060 ;
        RECT 49.070 87.340 49.330 87.660 ;
        RECT 36.590 83.640 36.850 83.960 ;
        RECT 45.230 83.640 45.490 83.960 ;
        RECT 35.150 82.160 35.410 82.480 ;
        RECT 36.110 82.160 36.370 82.480 ;
        RECT 35.210 79.890 35.350 82.160 ;
        RECT 35.150 79.570 35.410 79.890 ;
        RECT 36.170 72.490 36.310 82.160 ;
        RECT 36.650 75.450 36.790 83.640 ;
        RECT 44.270 83.270 44.530 83.590 ;
        RECT 43.790 75.870 44.050 76.190 ;
        RECT 36.590 75.130 36.850 75.450 ;
        RECT 43.310 75.130 43.570 75.450 ;
        RECT 36.110 72.170 36.370 72.490 ;
        RECT 42.830 67.730 43.090 68.050 ;
        RECT 35.630 67.360 35.890 67.680 ;
        RECT 36.590 67.360 36.850 67.680 ;
        RECT 38.990 67.360 39.250 67.680 ;
        RECT 35.690 67.040 35.830 67.360 ;
        RECT 35.690 66.900 36.310 67.040 ;
        RECT 36.170 62.130 36.310 66.900 ;
        RECT 36.110 61.810 36.370 62.130 ;
        RECT 36.650 54.730 36.790 67.360 ;
        RECT 38.030 62.920 38.290 63.240 ;
        RECT 38.090 59.910 38.230 62.920 ;
        RECT 38.510 61.810 38.770 62.130 ;
        RECT 38.030 59.590 38.290 59.910 ;
        RECT 36.590 54.410 36.850 54.730 ;
        RECT 36.580 50.500 36.860 50.870 ;
        RECT 36.590 50.340 36.850 50.500 ;
        RECT 35.150 50.200 35.410 50.290 ;
        RECT 36.110 50.200 36.370 50.290 ;
        RECT 35.150 50.060 36.370 50.200 ;
        RECT 35.150 49.970 35.410 50.060 ;
        RECT 36.110 49.970 36.370 50.060 ;
        RECT 35.630 49.600 35.890 49.920 ;
        RECT 35.690 46.960 35.830 49.600 ;
        RECT 35.630 46.640 35.890 46.960 ;
        RECT 38.090 43.260 38.230 59.590 ;
        RECT 38.570 55.100 38.710 61.810 ;
        RECT 38.510 54.780 38.770 55.100 ;
        RECT 39.050 53.990 39.190 67.360 ;
        RECT 42.890 67.310 43.030 67.730 ;
        RECT 42.830 66.990 43.090 67.310 ;
        RECT 39.460 62.340 39.740 62.710 ;
        RECT 39.530 62.130 39.670 62.340 ;
        RECT 39.470 61.810 39.730 62.130 ;
        RECT 42.830 58.480 43.090 58.800 ;
        RECT 42.350 55.890 42.610 56.210 ;
        RECT 38.990 53.670 39.250 53.990 ;
        RECT 39.470 53.670 39.730 53.990 ;
        RECT 39.530 51.770 39.670 53.670 ;
        RECT 39.470 51.450 39.730 51.770 ;
        RECT 42.410 46.590 42.550 55.890 ;
        RECT 42.890 54.730 43.030 58.480 ;
        RECT 42.830 54.410 43.090 54.730 ;
        RECT 42.890 51.030 43.030 54.410 ;
        RECT 42.830 50.710 43.090 51.030 ;
        RECT 42.890 46.590 43.030 50.710 ;
        RECT 42.350 46.270 42.610 46.590 ;
        RECT 42.830 46.270 43.090 46.590 ;
        RECT 38.030 42.940 38.290 43.260 ;
        RECT 40.910 42.940 41.170 43.260 ;
        RECT 35.140 42.360 35.420 42.730 ;
        RECT 34.190 38.870 34.450 39.190 ;
        RECT 35.210 35.120 35.350 42.360 ;
        RECT 40.970 39.930 41.110 42.940 ;
        RECT 40.910 39.610 41.170 39.930 ;
        RECT 36.110 38.130 36.370 38.450 ;
        RECT 35.150 34.800 35.410 35.120 ;
        RECT 35.630 34.060 35.890 34.380 ;
        RECT 35.690 33.640 35.830 34.060 ;
        RECT 35.630 33.320 35.890 33.640 ;
        RECT 35.150 30.360 35.410 30.680 ;
        RECT 33.710 29.990 33.970 30.310 ;
        RECT 34.670 29.620 34.930 29.940 ;
        RECT 33.710 29.250 33.970 29.570 ;
        RECT 33.770 27.720 33.910 29.250 ;
        RECT 33.710 27.400 33.970 27.720 ;
        RECT 32.750 27.030 33.010 27.350 ;
        RECT 34.730 25.500 34.870 29.620 ;
        RECT 35.210 26.240 35.350 30.360 ;
        RECT 35.690 26.240 35.830 33.320 ;
        RECT 36.170 30.310 36.310 38.130 ;
        RECT 38.510 37.760 38.770 38.080 ;
        RECT 37.550 30.730 37.810 31.050 ;
        RECT 36.110 29.990 36.370 30.310 ;
        RECT 36.170 26.610 36.310 29.990 ;
        RECT 36.110 26.290 36.370 26.610 ;
        RECT 35.150 25.920 35.410 26.240 ;
        RECT 35.630 25.920 35.890 26.240 ;
        RECT 34.670 25.180 34.930 25.500 ;
        RECT 35.210 23.280 35.350 25.920 ;
        RECT 35.150 22.960 35.410 23.280 ;
        RECT 29.390 21.850 29.650 22.170 ;
        RECT 33.230 21.110 33.490 21.430 ;
        RECT 33.290 18.470 33.430 21.110 ;
        RECT 37.610 18.470 37.750 30.730 ;
        RECT 38.570 26.980 38.710 37.760 ;
        RECT 40.430 37.390 40.690 37.710 ;
        RECT 38.510 26.660 38.770 26.980 ;
        RECT 40.490 26.610 40.630 37.390 ;
        RECT 42.410 35.030 42.550 46.270 ;
        RECT 43.370 46.220 43.510 75.130 ;
        RECT 43.850 71.380 43.990 75.870 ;
        RECT 43.790 71.060 44.050 71.380 ;
        RECT 43.790 55.150 44.050 55.470 ;
        RECT 43.310 45.900 43.570 46.220 ;
        RECT 42.410 34.890 43.030 35.030 ;
        RECT 42.350 34.430 42.610 34.750 ;
        RECT 42.410 31.790 42.550 34.430 ;
        RECT 42.350 31.470 42.610 31.790 ;
        RECT 42.410 30.680 42.550 31.470 ;
        RECT 42.350 30.360 42.610 30.680 ;
        RECT 39.470 26.290 39.730 26.610 ;
        RECT 40.430 26.290 40.690 26.610 ;
        RECT 39.530 18.470 39.670 26.290 ;
        RECT 42.890 23.280 43.030 34.890 ;
        RECT 43.850 27.350 43.990 55.150 ;
        RECT 44.330 54.730 44.470 83.270 ;
        RECT 44.750 75.500 45.010 75.820 ;
        RECT 44.270 54.410 44.530 54.730 ;
        RECT 44.810 46.960 44.950 75.500 ;
        RECT 45.290 71.750 45.430 83.640 ;
        RECT 45.710 78.090 45.970 78.410 ;
        RECT 45.770 76.560 45.910 78.090 ;
        RECT 45.710 76.240 45.970 76.560 ;
        RECT 47.630 75.500 47.890 75.820 ;
        RECT 47.690 72.120 47.830 75.500 ;
        RECT 47.630 71.800 47.890 72.120 ;
        RECT 49.130 71.750 49.270 87.340 ;
        RECT 52.970 87.290 53.110 94.740 ;
        RECT 53.390 91.780 53.650 92.100 ;
        RECT 53.450 88.770 53.590 91.780 ;
        RECT 53.390 88.450 53.650 88.770 ;
        RECT 53.930 87.660 54.070 100.290 ;
        RECT 54.410 99.500 54.550 103.250 ;
        RECT 54.350 99.180 54.610 99.500 ;
        RECT 54.830 98.440 55.090 98.760 ;
        RECT 54.890 96.910 55.030 98.440 ;
        RECT 54.830 96.590 55.090 96.910 ;
        RECT 55.370 96.750 55.510 106.580 ;
        RECT 56.810 100.240 56.950 115.830 ;
        RECT 61.070 115.460 61.330 115.780 ;
        RECT 61.130 108.750 61.270 115.460 ;
        RECT 61.070 108.430 61.330 108.750 ;
        RECT 61.610 107.270 61.750 116.200 ;
        RECT 62.030 111.020 62.290 111.340 ;
        RECT 61.550 106.950 61.810 107.270 ;
        RECT 61.610 105.050 61.750 106.950 ;
        RECT 61.550 104.730 61.810 105.050 ;
        RECT 57.230 102.880 57.490 103.200 ;
        RECT 58.190 102.880 58.450 103.200 ;
        RECT 56.750 99.920 57.010 100.240 ;
        RECT 55.300 96.380 55.580 96.750 ;
        RECT 56.810 96.540 56.950 99.920 ;
        RECT 57.290 99.500 57.430 102.880 ;
        RECT 57.710 99.550 57.970 99.870 ;
        RECT 57.230 99.180 57.490 99.500 ;
        RECT 55.370 87.660 55.510 96.380 ;
        RECT 56.750 96.220 57.010 96.540 ;
        RECT 57.770 95.800 57.910 99.550 ;
        RECT 58.250 99.130 58.390 102.880 ;
        RECT 62.090 100.240 62.230 111.020 ;
        RECT 61.070 99.920 61.330 100.240 ;
        RECT 62.030 99.920 62.290 100.240 ;
        RECT 58.190 98.810 58.450 99.130 ;
        RECT 61.130 96.170 61.270 99.920 ;
        RECT 62.570 99.870 62.710 119.530 ;
        RECT 64.910 115.090 65.170 115.410 ;
        RECT 64.430 111.390 64.690 111.710 ;
        RECT 62.510 99.550 62.770 99.870 ;
        RECT 64.490 96.540 64.630 111.390 ;
        RECT 64.430 96.220 64.690 96.540 ;
        RECT 61.070 95.850 61.330 96.170 ;
        RECT 57.710 95.480 57.970 95.800 ;
        RECT 57.230 94.740 57.490 95.060 ;
        RECT 53.870 87.340 54.130 87.660 ;
        RECT 55.310 87.340 55.570 87.660 ;
        RECT 52.910 86.970 53.170 87.290 ;
        RECT 49.550 84.380 49.810 84.700 ;
        RECT 49.610 83.130 49.750 84.380 ;
        RECT 49.610 82.990 50.710 83.130 ;
        RECT 50.570 82.850 50.710 82.990 ;
        RECT 50.510 82.530 50.770 82.850 ;
        RECT 55.790 74.020 56.050 74.340 ;
        RECT 45.230 71.430 45.490 71.750 ;
        RECT 46.670 71.430 46.930 71.750 ;
        RECT 49.070 71.430 49.330 71.750 ;
        RECT 46.730 62.500 46.870 71.430 ;
        RECT 54.350 71.060 54.610 71.380 ;
        RECT 48.110 70.690 48.370 71.010 ;
        RECT 47.630 69.950 47.890 70.270 ;
        RECT 46.670 62.180 46.930 62.500 ;
        RECT 46.670 58.850 46.930 59.170 ;
        RECT 45.230 55.520 45.490 55.840 ;
        RECT 45.290 48.070 45.430 55.520 ;
        RECT 46.730 54.360 46.870 58.850 ;
        RECT 47.690 54.730 47.830 69.950 ;
        RECT 47.630 54.410 47.890 54.730 ;
        RECT 46.670 54.040 46.930 54.360 ;
        RECT 48.170 50.290 48.310 70.690 ;
        RECT 49.550 70.320 49.810 70.640 ;
        RECT 49.610 55.470 49.750 70.320 ;
        RECT 53.870 67.730 54.130 68.050 ;
        RECT 50.030 66.990 50.290 67.310 ;
        RECT 49.550 55.150 49.810 55.470 ;
        RECT 49.610 51.030 49.750 55.150 ;
        RECT 50.090 51.770 50.230 66.990 ;
        RECT 53.390 66.250 53.650 66.570 ;
        RECT 50.510 65.880 50.770 66.200 ;
        RECT 50.570 63.610 50.710 65.880 ;
        RECT 50.510 63.290 50.770 63.610 ;
        RECT 53.450 59.910 53.590 66.250 ;
        RECT 52.430 59.590 52.690 59.910 ;
        RECT 53.390 59.590 53.650 59.910 ;
        RECT 51.950 58.480 52.210 58.800 ;
        RECT 52.010 55.100 52.150 58.480 ;
        RECT 51.950 54.780 52.210 55.100 ;
        RECT 50.030 51.450 50.290 51.770 ;
        RECT 49.550 50.710 49.810 51.030 ;
        RECT 52.490 50.660 52.630 59.590 ;
        RECT 52.910 54.780 53.170 55.100 ;
        RECT 52.430 50.340 52.690 50.660 ;
        RECT 48.110 49.970 48.370 50.290 ;
        RECT 45.230 47.750 45.490 48.070 ;
        RECT 44.750 46.640 45.010 46.960 ;
        RECT 45.290 39.470 45.430 47.750 ;
        RECT 48.170 45.850 48.310 49.970 ;
        RECT 52.430 47.010 52.690 47.330 ;
        RECT 48.110 45.530 48.370 45.850 ;
        RECT 50.510 43.910 50.770 44.000 ;
        RECT 52.490 43.910 52.630 47.010 ;
        RECT 52.970 46.960 53.110 54.780 ;
        RECT 53.450 47.240 53.590 59.590 ;
        RECT 53.930 59.170 54.070 67.730 ;
        RECT 54.410 59.170 54.550 71.060 ;
        RECT 55.850 64.350 55.990 74.020 ;
        RECT 57.290 72.120 57.430 94.740 ;
        RECT 62.030 94.370 62.290 94.690 ;
        RECT 62.090 92.470 62.230 94.370 ;
        RECT 62.030 92.150 62.290 92.470 ;
        RECT 57.710 91.780 57.970 92.100 ;
        RECT 57.770 88.770 57.910 91.780 ;
        RECT 63.950 91.040 64.210 91.360 ;
        RECT 64.010 88.770 64.150 91.040 ;
        RECT 64.490 88.770 64.630 96.220 ;
        RECT 57.710 88.450 57.970 88.770 ;
        RECT 63.950 88.450 64.210 88.770 ;
        RECT 64.430 88.450 64.690 88.770 ;
        RECT 59.150 87.340 59.410 87.660 ;
        RECT 58.190 75.130 58.450 75.450 ;
        RECT 57.230 71.800 57.490 72.120 ;
        RECT 58.250 68.050 58.390 75.130 ;
        RECT 58.190 67.730 58.450 68.050 ;
        RECT 57.710 67.360 57.970 67.680 ;
        RECT 55.790 64.030 56.050 64.350 ;
        RECT 57.230 62.180 57.490 62.500 ;
        RECT 53.870 58.850 54.130 59.170 ;
        RECT 54.350 58.850 54.610 59.170 ;
        RECT 56.750 58.850 57.010 59.170 ;
        RECT 55.310 57.740 55.570 58.060 ;
        RECT 53.450 47.100 54.070 47.240 ;
        RECT 52.910 46.640 53.170 46.960 ;
        RECT 50.510 43.770 52.630 43.910 ;
        RECT 50.510 43.680 50.770 43.770 ;
        RECT 45.290 39.330 45.910 39.470 ;
        RECT 45.230 38.870 45.490 39.190 ;
        RECT 44.750 38.130 45.010 38.450 ;
        RECT 44.810 34.750 44.950 38.130 ;
        RECT 44.750 34.430 45.010 34.750 ;
        RECT 43.790 27.030 44.050 27.350 ;
        RECT 42.830 22.960 43.090 23.280 ;
        RECT 33.230 18.150 33.490 18.470 ;
        RECT 37.550 18.150 37.810 18.470 ;
        RECT 39.470 18.150 39.730 18.470 ;
        RECT 42.890 17.730 43.030 22.960 ;
        RECT 45.290 18.100 45.430 38.870 ;
        RECT 45.230 17.780 45.490 18.100 ;
        RECT 45.770 17.730 45.910 39.330 ;
        RECT 48.110 38.500 48.370 38.820 ;
        RECT 48.170 29.940 48.310 38.500 ;
        RECT 50.030 37.760 50.290 38.080 ;
        RECT 48.110 29.620 48.370 29.940 ;
        RECT 47.630 29.250 47.890 29.570 ;
        RECT 47.690 22.170 47.830 29.250 ;
        RECT 47.630 21.850 47.890 22.170 ;
        RECT 50.090 18.750 50.230 37.760 ;
        RECT 51.470 34.430 51.730 34.750 ;
        RECT 51.530 31.050 51.670 34.430 ;
        RECT 51.470 30.730 51.730 31.050 ;
        RECT 52.910 22.590 53.170 22.910 ;
        RECT 50.090 18.610 51.670 18.750 ;
        RECT 51.530 18.470 51.670 18.610 ;
        RECT 52.970 18.470 53.110 22.590 ;
        RECT 53.390 21.110 53.650 21.430 ;
        RECT 53.450 19.580 53.590 21.110 ;
        RECT 53.390 19.260 53.650 19.580 ;
        RECT 51.470 18.150 51.730 18.470 ;
        RECT 52.910 18.150 53.170 18.470 ;
        RECT 42.830 17.410 43.090 17.730 ;
        RECT 45.710 17.410 45.970 17.730 ;
        RECT 53.930 17.360 54.070 47.100 ;
        RECT 54.830 46.640 55.090 46.960 ;
        RECT 54.890 43.630 55.030 46.640 ;
        RECT 54.830 43.310 55.090 43.630 ;
        RECT 54.350 42.940 54.610 43.260 ;
        RECT 54.410 39.560 54.550 42.940 ;
        RECT 54.350 39.240 54.610 39.560 ;
        RECT 54.350 34.800 54.610 35.120 ;
        RECT 54.410 31.420 54.550 34.800 ;
        RECT 54.350 31.100 54.610 31.420 ;
        RECT 55.370 30.680 55.510 57.740 ;
        RECT 56.270 54.040 56.530 54.360 ;
        RECT 56.330 42.890 56.470 54.040 ;
        RECT 56.270 42.570 56.530 42.890 ;
        RECT 56.810 41.780 56.950 58.850 ;
        RECT 56.750 41.460 57.010 41.780 ;
        RECT 57.290 37.710 57.430 62.180 ;
        RECT 57.770 62.130 57.910 67.360 ;
        RECT 57.710 61.810 57.970 62.130 ;
        RECT 58.670 55.520 58.930 55.840 ;
        RECT 57.710 55.150 57.970 55.470 ;
        RECT 57.770 54.360 57.910 55.150 ;
        RECT 58.730 55.100 58.870 55.520 ;
        RECT 58.670 54.780 58.930 55.100 ;
        RECT 57.710 54.040 57.970 54.360 ;
        RECT 58.670 50.340 58.930 50.660 ;
        RECT 58.190 45.900 58.450 46.220 ;
        RECT 58.250 42.890 58.390 45.900 ;
        RECT 58.190 42.570 58.450 42.890 ;
        RECT 57.710 38.130 57.970 38.450 ;
        RECT 57.230 37.390 57.490 37.710 ;
        RECT 57.290 33.640 57.430 37.390 ;
        RECT 57.770 35.860 57.910 38.130 ;
        RECT 57.710 35.540 57.970 35.860 ;
        RECT 57.230 33.320 57.490 33.640 ;
        RECT 55.310 30.360 55.570 30.680 ;
        RECT 56.270 26.290 56.530 26.610 ;
        RECT 56.330 19.580 56.470 26.290 ;
        RECT 56.270 19.260 56.530 19.580 ;
        RECT 57.290 18.840 57.430 33.320 ;
        RECT 58.730 26.610 58.870 50.340 ;
        RECT 59.210 46.220 59.350 87.340 ;
        RECT 60.110 86.970 60.370 87.290 ;
        RECT 59.630 83.270 59.890 83.590 ;
        RECT 59.690 70.270 59.830 83.270 ;
        RECT 60.170 80.630 60.310 86.970 ;
        RECT 64.970 83.320 65.110 115.090 ;
        RECT 66.410 112.080 66.550 137.290 ;
        RECT 70.730 136.870 70.870 143.210 ;
        RECT 77.930 140.940 78.070 143.950 ;
        RECT 86.030 143.210 86.290 143.530 ;
        RECT 98.510 143.210 98.770 143.530 ;
        RECT 86.090 141.680 86.230 143.210 ;
        RECT 86.030 141.360 86.290 141.680 ;
        RECT 98.570 141.310 98.710 143.210 ;
        RECT 98.510 140.990 98.770 141.310 ;
        RECT 77.870 140.620 78.130 140.940 ;
        RECT 86.990 140.620 87.250 140.940 ;
        RECT 78.350 139.510 78.610 139.830 ;
        RECT 74.990 139.140 75.250 139.460 ;
        RECT 70.670 136.550 70.930 136.870 ;
        RECT 75.050 120.960 75.190 139.140 ;
        RECT 78.410 136.500 78.550 139.510 ;
        RECT 87.050 136.870 87.190 140.620 ;
        RECT 99.530 139.830 99.670 143.950 ;
        RECT 106.670 143.210 106.930 143.530 ;
        RECT 106.730 141.310 106.870 143.210 ;
        RECT 106.670 140.990 106.930 141.310 ;
        RECT 101.390 140.620 101.650 140.940 ;
        RECT 99.470 139.510 99.730 139.830 ;
        RECT 93.710 139.140 93.970 139.460 ;
        RECT 86.990 136.550 87.250 136.870 ;
        RECT 93.770 136.500 93.910 139.140 ;
        RECT 99.530 137.240 99.670 139.510 ;
        RECT 100.910 139.140 101.170 139.460 ;
        RECT 99.470 136.920 99.730 137.240 ;
        RECT 100.970 136.500 101.110 139.140 ;
        RECT 101.450 136.870 101.590 140.620 ;
        RECT 101.390 136.550 101.650 136.870 ;
        RECT 110.990 136.550 111.250 136.870 ;
        RECT 78.350 136.180 78.610 136.500 ;
        RECT 93.710 136.180 93.970 136.500 ;
        RECT 100.910 136.180 101.170 136.500 ;
        RECT 102.830 136.180 103.090 136.500 ;
        RECT 77.390 135.810 77.650 136.130 ;
        RECT 85.070 135.810 85.330 136.130 ;
        RECT 76.430 131.000 76.690 131.320 ;
        RECT 75.470 127.670 75.730 127.990 ;
        RECT 75.530 124.290 75.670 127.670 ;
        RECT 76.490 124.290 76.630 131.000 ;
        RECT 77.450 125.400 77.590 135.810 ;
        RECT 79.310 132.110 79.570 132.430 ;
        RECT 80.270 132.110 80.530 132.430 ;
        RECT 79.370 128.360 79.510 132.110 ;
        RECT 79.310 128.040 79.570 128.360 ;
        RECT 80.330 127.250 80.470 132.110 ;
        RECT 83.630 131.370 83.890 131.690 ;
        RECT 81.230 131.000 81.490 131.320 ;
        RECT 80.270 126.930 80.530 127.250 ;
        RECT 77.390 125.080 77.650 125.400 ;
        RECT 81.290 124.660 81.430 131.000 ;
        RECT 83.690 128.360 83.830 131.370 ;
        RECT 83.630 128.040 83.890 128.360 ;
        RECT 83.150 127.670 83.410 127.990 ;
        RECT 81.230 124.340 81.490 124.660 ;
        RECT 75.470 123.970 75.730 124.290 ;
        RECT 76.430 123.970 76.690 124.290 ;
        RECT 74.990 120.640 75.250 120.960 ;
        RECT 68.750 120.270 69.010 120.590 ;
        RECT 66.350 111.760 66.610 112.080 ;
        RECT 65.390 111.020 65.650 111.340 ;
        RECT 65.450 108.010 65.590 111.020 ;
        RECT 65.390 107.690 65.650 108.010 ;
        RECT 65.390 102.880 65.650 103.200 ;
        RECT 65.450 100.980 65.590 102.880 ;
        RECT 65.390 100.660 65.650 100.980 ;
        RECT 66.410 96.910 66.550 111.760 ;
        RECT 68.810 99.870 68.950 120.270 ;
        RECT 71.630 118.790 71.890 119.110 ;
        RECT 71.690 116.890 71.830 118.790 ;
        RECT 71.630 116.570 71.890 116.890 ;
        RECT 72.110 115.460 72.370 115.780 ;
        RECT 71.630 115.090 71.890 115.410 ;
        RECT 69.230 108.430 69.490 108.750 ;
        RECT 68.750 99.550 69.010 99.870 ;
        RECT 67.310 99.180 67.570 99.500 ;
        RECT 67.370 96.910 67.510 99.180 ;
        RECT 69.290 98.760 69.430 108.430 ;
        RECT 69.230 98.440 69.490 98.760 ;
        RECT 66.350 96.590 66.610 96.910 ;
        RECT 67.310 96.590 67.570 96.910 ;
        RECT 71.150 90.300 71.410 90.620 ;
        RECT 71.210 86.920 71.350 90.300 ;
        RECT 71.150 86.600 71.410 86.920 ;
        RECT 64.970 83.180 65.590 83.320 ;
        RECT 64.910 82.160 65.170 82.480 ;
        RECT 60.110 80.310 60.370 80.630 ;
        RECT 60.170 75.820 60.310 80.310 ;
        RECT 60.110 75.500 60.370 75.820 ;
        RECT 64.430 71.060 64.690 71.380 ;
        RECT 61.550 70.320 61.810 70.640 ;
        RECT 59.630 69.950 59.890 70.270 ;
        RECT 61.610 67.310 61.750 70.320 ;
        RECT 61.550 66.990 61.810 67.310 ;
        RECT 64.490 58.800 64.630 71.060 ;
        RECT 64.970 60.280 65.110 82.160 ;
        RECT 65.450 76.560 65.590 83.180 ;
        RECT 70.670 79.200 70.930 79.520 ;
        RECT 70.190 78.830 70.450 79.150 ;
        RECT 65.390 76.240 65.650 76.560 ;
        RECT 68.270 70.690 68.530 71.010 ;
        RECT 68.330 64.350 68.470 70.690 ;
        RECT 69.710 68.100 69.970 68.420 ;
        RECT 69.770 64.350 69.910 68.100 ;
        RECT 70.250 64.350 70.390 78.830 ;
        RECT 70.730 71.010 70.870 79.200 ;
        RECT 71.690 79.150 71.830 115.090 ;
        RECT 72.170 113.190 72.310 115.460 ;
        RECT 72.110 112.870 72.370 113.190 ;
        RECT 74.990 111.760 75.250 112.080 ;
        RECT 72.110 106.580 72.370 106.900 ;
        RECT 72.170 104.040 72.310 106.580 ;
        RECT 72.170 103.900 72.790 104.040 ;
        RECT 72.650 99.870 72.790 103.900 ;
        RECT 75.050 100.610 75.190 111.760 ;
        RECT 74.990 100.290 75.250 100.610 ;
        RECT 75.530 100.240 75.670 123.970 ;
        RECT 78.350 119.900 78.610 120.220 ;
        RECT 79.790 119.900 80.050 120.220 ;
        RECT 76.430 102.880 76.690 103.200 ;
        RECT 75.470 99.920 75.730 100.240 ;
        RECT 72.590 99.550 72.850 99.870 ;
        RECT 72.110 95.110 72.370 95.430 ;
        RECT 72.170 91.730 72.310 95.110 ;
        RECT 72.110 91.410 72.370 91.730 ;
        RECT 72.110 84.010 72.370 84.330 ;
        RECT 72.170 80.260 72.310 84.010 ;
        RECT 72.110 79.940 72.370 80.260 ;
        RECT 72.650 79.620 72.790 99.550 ;
        RECT 76.490 96.910 76.630 102.880 ;
        RECT 78.410 100.980 78.550 119.900 ;
        RECT 78.830 119.530 79.090 119.850 ;
        RECT 78.350 100.660 78.610 100.980 ;
        RECT 76.430 96.590 76.690 96.910 ;
        RECT 78.890 95.060 79.030 119.530 ;
        RECT 79.850 117.360 79.990 119.900 ;
        RECT 81.710 118.790 81.970 119.110 ;
        RECT 79.850 117.220 80.470 117.360 ;
        RECT 79.310 110.650 79.570 110.970 ;
        RECT 79.370 108.380 79.510 110.650 ;
        RECT 79.310 108.060 79.570 108.380 ;
        RECT 79.790 106.580 80.050 106.900 ;
        RECT 79.850 103.570 79.990 106.580 ;
        RECT 79.790 103.250 80.050 103.570 ;
        RECT 79.310 95.110 79.570 95.430 ;
        RECT 78.830 94.740 79.090 95.060 ;
        RECT 79.370 92.100 79.510 95.110 ;
        RECT 79.310 91.780 79.570 92.100 ;
        RECT 79.790 91.410 80.050 91.730 ;
        RECT 74.990 86.230 75.250 86.550 ;
        RECT 79.850 86.280 79.990 91.410 ;
        RECT 80.330 86.920 80.470 117.220 ;
        RECT 80.750 111.020 81.010 111.340 ;
        RECT 80.810 108.010 80.950 111.020 ;
        RECT 81.770 108.010 81.910 118.790 ;
        RECT 82.670 116.200 82.930 116.520 ;
        RECT 82.730 113.190 82.870 116.200 ;
        RECT 82.670 112.870 82.930 113.190 ;
        RECT 82.190 111.390 82.450 111.710 ;
        RECT 80.750 107.690 81.010 108.010 ;
        RECT 81.710 107.690 81.970 108.010 ;
        RECT 82.250 103.570 82.390 111.390 ;
        RECT 82.670 108.060 82.930 108.380 ;
        RECT 82.190 103.250 82.450 103.570 ;
        RECT 81.230 100.660 81.490 100.980 ;
        RECT 81.290 95.060 81.430 100.660 ;
        RECT 81.230 94.740 81.490 95.060 ;
        RECT 80.270 86.600 80.530 86.920 ;
        RECT 75.050 84.330 75.190 86.230 ;
        RECT 79.850 86.140 80.470 86.280 ;
        RECT 74.990 84.010 75.250 84.330 ;
        RECT 79.310 84.010 79.570 84.330 ;
        RECT 72.170 79.480 72.790 79.620 ;
        RECT 71.630 78.830 71.890 79.150 ;
        RECT 71.150 75.870 71.410 76.190 ;
        RECT 70.670 70.690 70.930 71.010 ;
        RECT 68.270 64.030 68.530 64.350 ;
        RECT 69.710 64.030 69.970 64.350 ;
        RECT 70.190 64.030 70.450 64.350 ;
        RECT 71.210 62.500 71.350 75.870 ;
        RECT 71.630 63.660 71.890 63.980 ;
        RECT 71.690 62.870 71.830 63.660 ;
        RECT 72.170 63.240 72.310 79.480 ;
        RECT 72.590 78.460 72.850 78.780 ;
        RECT 72.650 76.190 72.790 78.460 ;
        RECT 72.590 75.870 72.850 76.190 ;
        RECT 79.370 75.820 79.510 84.010 ;
        RECT 79.790 82.160 80.050 82.480 ;
        RECT 79.850 80.630 79.990 82.160 ;
        RECT 79.790 80.310 80.050 80.630 ;
        RECT 79.310 75.500 79.570 75.820 ;
        RECT 79.370 74.340 79.510 75.500 ;
        RECT 79.310 74.020 79.570 74.340 ;
        RECT 74.990 71.060 75.250 71.380 ;
        RECT 79.310 71.060 79.570 71.380 ;
        RECT 75.050 67.310 75.190 71.060 ;
        RECT 76.910 70.690 77.170 71.010 ;
        RECT 76.970 67.680 77.110 70.690 ;
        RECT 79.370 68.420 79.510 71.060 ;
        RECT 79.310 68.100 79.570 68.420 ;
        RECT 80.330 68.050 80.470 86.140 ;
        RECT 82.730 76.190 82.870 108.060 ;
        RECT 83.210 100.980 83.350 127.670 ;
        RECT 83.690 109.120 83.830 128.040 ;
        RECT 85.130 115.780 85.270 135.810 ;
        RECT 93.770 132.800 93.910 136.180 ;
        RECT 94.190 135.810 94.450 136.130 ;
        RECT 93.710 132.480 93.970 132.800 ;
        RECT 87.950 132.110 88.210 132.430 ;
        RECT 88.010 129.470 88.150 132.110 ;
        RECT 87.950 129.150 88.210 129.470 ;
        RECT 94.250 125.400 94.390 135.810 ;
        RECT 99.950 132.160 100.210 132.430 ;
        RECT 99.950 132.110 100.630 132.160 ;
        RECT 100.010 132.020 100.630 132.110 ;
        RECT 100.490 128.360 100.630 132.020 ;
        RECT 100.970 128.730 101.110 136.180 ;
        RECT 101.870 135.810 102.130 136.130 ;
        RECT 101.930 133.540 102.070 135.810 ;
        RECT 102.350 135.440 102.610 135.760 ;
        RECT 101.870 133.220 102.130 133.540 ;
        RECT 102.410 132.800 102.550 135.440 ;
        RECT 101.390 132.480 101.650 132.800 ;
        RECT 102.350 132.480 102.610 132.800 ;
        RECT 101.450 129.470 101.590 132.480 ;
        RECT 101.390 129.150 101.650 129.470 ;
        RECT 100.910 128.410 101.170 128.730 ;
        RECT 95.150 128.040 95.410 128.360 ;
        RECT 100.430 128.040 100.690 128.360 ;
        RECT 94.190 125.080 94.450 125.400 ;
        RECT 89.870 124.340 90.130 124.660 ;
        RECT 88.430 121.010 88.690 121.330 ;
        RECT 86.030 120.640 86.290 120.960 ;
        RECT 85.550 119.530 85.810 119.850 ;
        RECT 85.070 115.460 85.330 115.780 ;
        RECT 85.130 111.340 85.270 115.460 ;
        RECT 85.070 111.020 85.330 111.340 ;
        RECT 83.630 108.800 83.890 109.120 ;
        RECT 85.070 108.800 85.330 109.120 ;
        RECT 85.130 107.640 85.270 108.800 ;
        RECT 85.610 108.010 85.750 119.530 ;
        RECT 86.090 117.260 86.230 120.640 ;
        RECT 86.030 116.940 86.290 117.260 ;
        RECT 86.090 112.450 86.230 116.940 ;
        RECT 88.490 116.890 88.630 121.010 ;
        RECT 89.930 119.480 90.070 124.340 ;
        RECT 95.210 124.290 95.350 128.040 ;
        RECT 98.030 124.340 98.290 124.660 ;
        RECT 95.150 123.970 95.410 124.290 ;
        RECT 97.550 123.970 97.810 124.290 ;
        RECT 94.670 120.270 94.930 120.590 ;
        RECT 94.190 119.530 94.450 119.850 ;
        RECT 89.870 119.160 90.130 119.480 ;
        RECT 93.710 119.160 93.970 119.480 ;
        RECT 88.430 116.570 88.690 116.890 ;
        RECT 89.930 116.520 90.070 119.160 ;
        RECT 89.870 116.200 90.130 116.520 ;
        RECT 87.950 114.720 88.210 115.040 ;
        RECT 86.030 112.130 86.290 112.450 ;
        RECT 86.510 111.390 86.770 111.710 ;
        RECT 85.550 107.690 85.810 108.010 ;
        RECT 86.030 107.690 86.290 108.010 ;
        RECT 85.070 107.320 85.330 107.640 ;
        RECT 85.130 103.940 85.270 107.320 ;
        RECT 85.610 105.050 85.750 107.690 ;
        RECT 85.550 104.730 85.810 105.050 ;
        RECT 85.070 103.620 85.330 103.940 ;
        RECT 85.550 103.250 85.810 103.570 ;
        RECT 83.150 100.660 83.410 100.980 ;
        RECT 84.110 94.370 84.370 94.690 ;
        RECT 84.170 78.780 84.310 94.370 ;
        RECT 85.610 91.730 85.750 103.250 ;
        RECT 86.090 96.540 86.230 107.690 ;
        RECT 86.570 107.270 86.710 111.390 ;
        RECT 88.010 108.380 88.150 114.720 ;
        RECT 87.950 108.060 88.210 108.380 ;
        RECT 86.510 106.950 86.770 107.270 ;
        RECT 86.030 96.220 86.290 96.540 ;
        RECT 86.980 96.380 87.260 96.750 ;
        RECT 89.930 96.540 90.070 116.200 ;
        RECT 93.770 113.190 93.910 119.160 ;
        RECT 93.710 112.870 93.970 113.190 ;
        RECT 91.790 111.390 92.050 111.710 ;
        RECT 91.850 108.750 91.990 111.390 ;
        RECT 91.790 108.430 92.050 108.750 ;
        RECT 94.250 103.940 94.390 119.530 ;
        RECT 94.730 108.010 94.870 120.270 ;
        RECT 95.210 119.850 95.350 123.970 ;
        RECT 97.610 119.850 97.750 123.970 ;
        RECT 95.150 119.530 95.410 119.850 ;
        RECT 97.550 119.530 97.810 119.850 ;
        RECT 95.150 118.790 95.410 119.110 ;
        RECT 95.210 116.150 95.350 118.790 ;
        RECT 95.150 115.830 95.410 116.150 ;
        RECT 96.110 115.830 96.370 116.150 ;
        RECT 96.170 111.710 96.310 115.830 ;
        RECT 97.610 115.410 97.750 119.530 ;
        RECT 97.550 115.090 97.810 115.410 ;
        RECT 96.110 111.390 96.370 111.710 ;
        RECT 94.670 107.690 94.930 108.010 ;
        RECT 98.090 105.050 98.230 124.340 ;
        RECT 100.490 124.290 100.630 128.040 ;
        RECT 100.910 127.670 101.170 127.990 ;
        RECT 100.430 123.970 100.690 124.290 ;
        RECT 100.430 111.760 100.690 112.080 ;
        RECT 100.490 108.010 100.630 111.760 ;
        RECT 100.430 107.690 100.690 108.010 ;
        RECT 98.030 104.730 98.290 105.050 ;
        RECT 92.750 103.620 93.010 103.940 ;
        RECT 94.190 103.620 94.450 103.940 ;
        RECT 87.050 96.170 87.190 96.380 ;
        RECT 89.870 96.220 90.130 96.540 ;
        RECT 86.990 95.850 87.250 96.170 ;
        RECT 90.350 95.480 90.610 95.800 ;
        RECT 86.510 95.110 86.770 95.430 ;
        RECT 85.550 91.410 85.810 91.730 ;
        RECT 86.570 88.770 86.710 95.110 ;
        RECT 87.950 94.740 88.210 95.060 ;
        RECT 86.510 88.450 86.770 88.770 ;
        RECT 88.010 87.660 88.150 94.740 ;
        RECT 90.410 92.470 90.550 95.480 ;
        RECT 92.810 92.840 92.950 103.620 ;
        RECT 93.230 99.180 93.490 99.500 ;
        RECT 93.290 95.800 93.430 99.180 ;
        RECT 100.490 99.130 100.630 107.690 ;
        RECT 100.970 100.610 101.110 127.670 ;
        RECT 101.390 124.340 101.650 124.660 ;
        RECT 101.870 124.340 102.130 124.660 ;
        RECT 101.450 116.150 101.590 124.340 ;
        RECT 101.930 120.960 102.070 124.340 ;
        RECT 101.870 120.640 102.130 120.960 ;
        RECT 101.930 116.520 102.070 120.640 ;
        RECT 102.410 120.590 102.550 132.480 ;
        RECT 102.890 132.430 103.030 136.180 ;
        RECT 107.630 135.070 107.890 135.390 ;
        RECT 107.690 133.540 107.830 135.070 ;
        RECT 107.630 133.220 107.890 133.540 ;
        RECT 111.050 132.430 111.190 136.550 ;
        RECT 117.290 136.130 117.430 144.690 ;
        RECT 111.470 135.810 111.730 136.130 ;
        RECT 117.230 135.810 117.490 136.130 ;
        RECT 118.670 135.810 118.930 136.130 ;
        RECT 102.830 132.110 103.090 132.430 ;
        RECT 103.310 132.110 103.570 132.430 ;
        RECT 107.630 132.110 107.890 132.430 ;
        RECT 110.990 132.110 111.250 132.430 ;
        RECT 103.370 128.360 103.510 132.110 ;
        RECT 103.310 128.040 103.570 128.360 ;
        RECT 107.690 125.030 107.830 132.110 ;
        RECT 111.050 129.470 111.190 132.110 ;
        RECT 110.990 129.150 111.250 129.470 ;
        RECT 107.630 124.710 107.890 125.030 ;
        RECT 103.790 123.970 104.050 124.290 ;
        RECT 104.750 123.970 105.010 124.290 ;
        RECT 103.850 121.330 103.990 123.970 ;
        RECT 103.790 121.010 104.050 121.330 ;
        RECT 102.350 120.270 102.610 120.590 ;
        RECT 104.810 116.520 104.950 123.970 ;
        RECT 108.110 122.860 108.370 123.180 ;
        RECT 106.670 119.900 106.930 120.220 ;
        RECT 107.150 119.900 107.410 120.220 ;
        RECT 106.730 117.260 106.870 119.900 ;
        RECT 106.670 116.940 106.930 117.260 ;
        RECT 101.870 116.200 102.130 116.520 ;
        RECT 104.750 116.200 105.010 116.520 ;
        RECT 101.390 115.830 101.650 116.150 ;
        RECT 107.210 112.450 107.350 119.900 ;
        RECT 108.170 119.480 108.310 122.860 ;
        RECT 108.110 119.160 108.370 119.480 ;
        RECT 108.590 118.790 108.850 119.110 ;
        RECT 108.650 116.150 108.790 118.790 ;
        RECT 111.050 116.520 111.190 129.150 ;
        RECT 110.990 116.200 111.250 116.520 ;
        RECT 108.590 116.060 108.850 116.150 ;
        RECT 108.590 115.920 109.270 116.060 ;
        RECT 108.590 115.830 108.850 115.920 ;
        RECT 107.150 112.130 107.410 112.450 ;
        RECT 105.710 111.020 105.970 111.340 ;
        RECT 102.350 107.690 102.610 108.010 ;
        RECT 103.310 107.690 103.570 108.010 ;
        RECT 102.410 103.570 102.550 107.690 ;
        RECT 101.390 103.250 101.650 103.570 ;
        RECT 102.350 103.250 102.610 103.570 ;
        RECT 100.910 100.290 101.170 100.610 ;
        RECT 101.450 100.240 101.590 103.250 ;
        RECT 102.410 100.610 102.550 103.250 ;
        RECT 102.350 100.290 102.610 100.610 ;
        RECT 101.390 99.920 101.650 100.240 ;
        RECT 101.450 99.600 101.590 99.920 ;
        RECT 100.970 99.460 101.590 99.600 ;
        RECT 101.870 99.550 102.130 99.870 ;
        RECT 100.430 98.810 100.690 99.130 ;
        RECT 93.230 95.480 93.490 95.800 ;
        RECT 100.970 95.060 101.110 99.460 ;
        RECT 101.390 96.590 101.650 96.910 ;
        RECT 93.230 94.740 93.490 95.060 ;
        RECT 100.910 94.740 101.170 95.060 ;
        RECT 92.750 92.520 93.010 92.840 ;
        RECT 90.350 92.150 90.610 92.470 ;
        RECT 92.270 91.410 92.530 91.730 ;
        RECT 92.750 91.410 93.010 91.730 ;
        RECT 86.510 87.340 86.770 87.660 ;
        RECT 87.950 87.340 88.210 87.660 ;
        RECT 86.570 84.330 86.710 87.340 ;
        RECT 92.330 87.290 92.470 91.410 ;
        RECT 92.270 86.970 92.530 87.290 ;
        RECT 86.510 84.010 86.770 84.330 ;
        RECT 84.590 83.640 84.850 83.960 ;
        RECT 84.110 78.460 84.370 78.780 ;
        RECT 84.650 78.410 84.790 83.640 ;
        RECT 91.790 83.270 92.050 83.590 ;
        RECT 85.070 82.900 85.330 83.220 ;
        RECT 85.130 79.520 85.270 82.900 ;
        RECT 91.850 82.850 91.990 83.270 ;
        RECT 91.790 82.530 92.050 82.850 ;
        RECT 90.830 82.160 91.090 82.480 ;
        RECT 85.070 79.200 85.330 79.520 ;
        RECT 84.590 78.090 84.850 78.410 ;
        RECT 82.670 75.870 82.930 76.190 ;
        RECT 84.650 75.820 84.790 78.090 ;
        RECT 84.590 75.500 84.850 75.820 ;
        RECT 90.890 75.450 91.030 82.160 ;
        RECT 91.850 79.520 91.990 82.530 ;
        RECT 91.790 79.200 92.050 79.520 ;
        RECT 91.850 78.780 91.990 79.200 ;
        RECT 91.790 78.460 92.050 78.780 ;
        RECT 85.070 75.130 85.330 75.450 ;
        RECT 85.550 75.130 85.810 75.450 ;
        RECT 90.830 75.130 91.090 75.450 ;
        RECT 85.130 72.490 85.270 75.130 ;
        RECT 85.070 72.170 85.330 72.490 ;
        RECT 84.110 70.320 84.370 70.640 ;
        RECT 82.670 68.100 82.930 68.420 ;
        RECT 80.270 67.730 80.530 68.050 ;
        RECT 76.910 67.360 77.170 67.680 ;
        RECT 74.990 66.990 75.250 67.310 ;
        RECT 75.470 66.620 75.730 66.940 ;
        RECT 72.110 62.920 72.370 63.240 ;
        RECT 75.530 62.870 75.670 66.620 ;
        RECT 80.330 66.570 80.470 67.730 ;
        RECT 80.270 66.250 80.530 66.570 ;
        RECT 82.730 64.350 82.870 68.100 ;
        RECT 84.170 67.680 84.310 70.320 ;
        RECT 85.610 68.420 85.750 75.130 ;
        RECT 90.830 74.020 91.090 74.340 ;
        RECT 86.990 71.060 87.250 71.380 ;
        RECT 85.550 68.100 85.810 68.420 ;
        RECT 84.110 67.360 84.370 67.680 ;
        RECT 87.050 64.350 87.190 71.060 ;
        RECT 90.890 68.050 91.030 74.020 ;
        RECT 91.850 70.640 91.990 78.460 ;
        RECT 91.790 70.320 92.050 70.640 ;
        RECT 90.830 67.730 91.090 68.050 ;
        RECT 82.670 64.030 82.930 64.350 ;
        RECT 86.990 64.030 87.250 64.350 ;
        RECT 87.950 62.920 88.210 63.240 ;
        RECT 71.630 62.550 71.890 62.870 ;
        RECT 75.470 62.550 75.730 62.870 ;
        RECT 87.470 62.550 87.730 62.870 ;
        RECT 71.150 62.180 71.410 62.500 ;
        RECT 71.690 60.280 71.830 62.550 ;
        RECT 72.110 62.180 72.370 62.500 ;
        RECT 86.990 62.180 87.250 62.500 ;
        RECT 64.910 59.960 65.170 60.280 ;
        RECT 71.630 59.960 71.890 60.280 ;
        RECT 64.430 58.480 64.690 58.800 ;
        RECT 61.070 58.110 61.330 58.430 ;
        RECT 60.110 51.450 60.370 51.770 ;
        RECT 60.170 46.960 60.310 51.450 ;
        RECT 61.130 51.400 61.270 58.110 ;
        RECT 67.790 54.410 68.050 54.730 ;
        RECT 61.070 51.080 61.330 51.400 ;
        RECT 61.550 50.710 61.810 51.030 ;
        RECT 61.610 47.700 61.750 50.710 ;
        RECT 61.550 47.380 61.810 47.700 ;
        RECT 66.350 47.380 66.610 47.700 ;
        RECT 60.110 46.640 60.370 46.960 ;
        RECT 66.410 46.590 66.550 47.380 ;
        RECT 66.830 46.640 67.090 46.960 ;
        RECT 66.350 46.270 66.610 46.590 ;
        RECT 59.150 45.900 59.410 46.220 ;
        RECT 65.870 45.900 66.130 46.220 ;
        RECT 59.150 42.940 59.410 43.260 ;
        RECT 59.210 34.750 59.350 42.940 ;
        RECT 59.630 42.570 59.890 42.890 ;
        RECT 64.910 42.570 65.170 42.890 ;
        RECT 59.690 38.820 59.830 42.570 ;
        RECT 59.630 38.500 59.890 38.820 ;
        RECT 64.970 38.450 65.110 42.570 ;
        RECT 64.910 38.130 65.170 38.450 ;
        RECT 60.590 35.170 60.850 35.490 ;
        RECT 59.150 34.430 59.410 34.750 ;
        RECT 59.210 30.680 59.350 34.430 ;
        RECT 59.630 31.100 59.890 31.420 ;
        RECT 59.150 30.360 59.410 30.680 ;
        RECT 58.670 26.290 58.930 26.610 ;
        RECT 59.690 18.840 59.830 31.100 ;
        RECT 60.650 30.310 60.790 35.170 ;
        RECT 63.470 34.060 63.730 34.380 ;
        RECT 64.910 34.060 65.170 34.380 ;
        RECT 60.590 29.990 60.850 30.310 ;
        RECT 62.500 29.780 62.780 30.150 ;
        RECT 62.510 29.620 62.770 29.780 ;
        RECT 57.230 18.520 57.490 18.840 ;
        RECT 59.630 18.520 59.890 18.840 ;
        RECT 63.530 18.470 63.670 34.060 ;
        RECT 64.970 25.870 65.110 34.060 ;
        RECT 65.390 29.990 65.650 30.310 ;
        RECT 65.450 26.610 65.590 29.990 ;
        RECT 65.390 26.290 65.650 26.610 ;
        RECT 64.910 25.550 65.170 25.870 ;
        RECT 64.910 22.960 65.170 23.280 ;
        RECT 64.430 18.890 64.690 19.210 ;
        RECT 63.470 18.150 63.730 18.470 ;
        RECT 64.490 17.730 64.630 18.890 ;
        RECT 64.430 17.410 64.690 17.730 ;
        RECT 24.110 17.040 24.370 17.360 ;
        RECT 41.870 17.040 42.130 17.360 ;
        RECT 53.870 17.040 54.130 17.360 ;
        RECT 41.930 15.880 42.070 17.040 ;
        RECT 64.970 16.720 65.110 22.960 ;
        RECT 65.930 19.580 66.070 45.900 ;
        RECT 66.410 42.890 66.550 46.270 ;
        RECT 66.350 42.570 66.610 42.890 ;
        RECT 66.890 42.520 67.030 46.640 ;
        RECT 66.830 42.200 67.090 42.520 ;
        RECT 66.350 34.800 66.610 35.120 ;
        RECT 66.410 19.580 66.550 34.800 ;
        RECT 66.890 23.280 67.030 42.200 ;
        RECT 67.310 23.330 67.570 23.650 ;
        RECT 66.830 22.960 67.090 23.280 ;
        RECT 66.830 21.110 67.090 21.430 ;
        RECT 65.870 19.260 66.130 19.580 ;
        RECT 66.350 19.260 66.610 19.580 ;
        RECT 65.930 18.840 66.070 19.260 ;
        RECT 65.870 18.520 66.130 18.840 ;
        RECT 66.890 17.730 67.030 21.110 ;
        RECT 67.370 18.840 67.510 23.330 ;
        RECT 67.850 22.910 67.990 54.410 ;
        RECT 68.270 50.710 68.530 51.030 ;
        RECT 68.330 26.980 68.470 50.710 ;
        RECT 72.170 48.070 72.310 62.180 ;
        RECT 77.870 61.810 78.130 62.130 ;
        RECT 76.430 59.220 76.690 59.540 ;
        RECT 75.950 55.890 76.210 56.210 ;
        RECT 72.590 51.450 72.850 51.770 ;
        RECT 72.110 47.750 72.370 48.070 ;
        RECT 72.170 41.140 72.310 47.750 ;
        RECT 72.650 42.150 72.790 51.450 ;
        RECT 76.010 51.400 76.150 55.890 ;
        RECT 75.950 51.080 76.210 51.400 ;
        RECT 74.990 50.710 75.250 51.030 ;
        RECT 75.050 50.290 75.190 50.710 ;
        RECT 74.990 49.970 75.250 50.290 ;
        RECT 72.590 41.830 72.850 42.150 ;
        RECT 72.170 41.000 72.790 41.140 ;
        RECT 68.750 38.500 69.010 38.820 ;
        RECT 68.810 27.350 68.950 38.500 ;
        RECT 69.220 29.780 69.500 30.150 ;
        RECT 68.750 27.030 69.010 27.350 ;
        RECT 68.270 26.660 68.530 26.980 ;
        RECT 67.790 22.590 68.050 22.910 ;
        RECT 67.310 18.520 67.570 18.840 ;
        RECT 68.750 18.380 69.010 18.470 ;
        RECT 69.290 18.380 69.430 29.780 ;
        RECT 72.110 29.250 72.370 29.570 ;
        RECT 72.170 22.170 72.310 29.250 ;
        RECT 72.110 21.850 72.370 22.170 ;
        RECT 69.710 21.110 69.970 21.430 ;
        RECT 69.770 18.470 69.910 21.110 ;
        RECT 72.650 19.580 72.790 41.000 ;
        RECT 75.050 39.930 75.190 49.970 ;
        RECT 74.990 39.610 75.250 39.930 ;
        RECT 76.490 19.580 76.630 59.220 ;
        RECT 76.910 42.940 77.170 43.260 ;
        RECT 76.970 26.610 77.110 42.940 ;
        RECT 76.910 26.290 77.170 26.610 ;
        RECT 72.590 19.260 72.850 19.580 ;
        RECT 76.430 19.260 76.690 19.580 ;
        RECT 77.930 18.840 78.070 61.810 ;
        RECT 87.050 55.100 87.190 62.180 ;
        RECT 86.990 54.780 87.250 55.100 ;
        RECT 82.670 54.410 82.930 54.730 ;
        RECT 78.830 53.670 79.090 53.990 ;
        RECT 78.890 51.770 79.030 53.670 ;
        RECT 82.730 52.140 82.870 54.410 ;
        RECT 82.670 51.820 82.930 52.140 ;
        RECT 78.830 51.450 79.090 51.770 ;
        RECT 81.230 50.340 81.490 50.660 ;
        RECT 79.790 41.460 80.050 41.780 ;
        RECT 78.830 34.800 79.090 35.120 ;
        RECT 78.890 23.650 79.030 34.800 ;
        RECT 79.850 31.790 79.990 41.460 ;
        RECT 81.290 39.930 81.430 50.340 ;
        RECT 83.150 45.530 83.410 45.850 ;
        RECT 83.210 39.930 83.350 45.530 ;
        RECT 85.070 42.570 85.330 42.890 ;
        RECT 81.230 39.610 81.490 39.930 ;
        RECT 83.150 39.610 83.410 39.930 ;
        RECT 81.290 34.750 81.430 39.610 ;
        RECT 85.130 38.450 85.270 42.570 ;
        RECT 87.050 38.820 87.190 54.780 ;
        RECT 87.530 54.360 87.670 62.550 ;
        RECT 88.010 59.540 88.150 62.920 ;
        RECT 87.950 59.220 88.210 59.540 ;
        RECT 90.890 56.210 91.030 67.730 ;
        RECT 92.810 66.940 92.950 91.410 ;
        RECT 93.290 70.270 93.430 94.740 ;
        RECT 97.550 91.780 97.810 92.100 ;
        RECT 97.610 87.660 97.750 91.780 ;
        RECT 98.990 87.710 99.250 88.030 ;
        RECT 97.550 87.340 97.810 87.660 ;
        RECT 95.150 79.940 95.410 80.260 ;
        RECT 95.210 79.520 95.350 79.940 ;
        RECT 95.150 79.200 95.410 79.520 ;
        RECT 95.210 75.920 95.350 79.200 ;
        RECT 95.210 75.820 96.790 75.920 ;
        RECT 93.710 75.500 93.970 75.820 ;
        RECT 95.210 75.780 96.850 75.820 ;
        RECT 96.590 75.500 96.850 75.780 ;
        RECT 93.770 72.490 93.910 75.500 ;
        RECT 99.050 75.450 99.190 87.710 ;
        RECT 100.430 86.970 100.690 87.290 ;
        RECT 100.490 79.520 100.630 86.970 ;
        RECT 101.450 83.960 101.590 96.590 ;
        RECT 101.930 92.840 102.070 99.550 ;
        RECT 103.370 96.910 103.510 107.690 ;
        RECT 105.770 103.570 105.910 111.020 ;
        RECT 107.210 109.120 107.350 112.130 ;
        RECT 107.150 108.800 107.410 109.120 ;
        RECT 108.590 108.430 108.850 108.750 ;
        RECT 105.710 103.250 105.970 103.570 ;
        RECT 104.270 99.920 104.530 100.240 ;
        RECT 107.630 99.920 107.890 100.240 ;
        RECT 104.330 96.910 104.470 99.920 ;
        RECT 103.310 96.590 103.570 96.910 ;
        RECT 104.270 96.590 104.530 96.910 ;
        RECT 107.690 95.430 107.830 99.920 ;
        RECT 108.650 95.800 108.790 108.430 ;
        RECT 109.130 108.380 109.270 115.920 ;
        RECT 110.030 114.720 110.290 115.040 ;
        RECT 110.090 112.080 110.230 114.720 ;
        RECT 110.030 111.760 110.290 112.080 ;
        RECT 109.070 108.060 109.330 108.380 ;
        RECT 109.130 106.900 109.270 108.060 ;
        RECT 109.070 106.580 109.330 106.900 ;
        RECT 109.550 103.620 109.810 103.940 ;
        RECT 108.110 95.480 108.370 95.800 ;
        RECT 108.590 95.480 108.850 95.800 ;
        RECT 107.630 95.110 107.890 95.430 ;
        RECT 101.870 92.520 102.130 92.840 ;
        RECT 107.150 92.520 107.410 92.840 ;
        RECT 102.350 91.780 102.610 92.100 ;
        RECT 101.390 83.640 101.650 83.960 ;
        RECT 101.390 79.940 101.650 80.260 ;
        RECT 100.430 79.200 100.690 79.520 ;
        RECT 101.450 76.190 101.590 79.940 ;
        RECT 102.410 78.780 102.550 91.780 ;
        RECT 107.210 88.770 107.350 92.520 ;
        RECT 107.150 88.450 107.410 88.770 ;
        RECT 103.310 87.340 103.570 87.660 ;
        RECT 103.370 80.630 103.510 87.340 ;
        RECT 104.270 86.230 104.530 86.550 ;
        RECT 103.310 80.310 103.570 80.630 ;
        RECT 104.330 79.890 104.470 86.230 ;
        RECT 107.690 84.700 107.830 95.110 ;
        RECT 108.170 91.730 108.310 95.480 ;
        RECT 109.610 95.060 109.750 103.620 ;
        RECT 111.530 103.570 111.670 135.810 ;
        RECT 118.190 135.070 118.450 135.390 ;
        RECT 118.250 133.540 118.390 135.070 ;
        RECT 118.190 133.220 118.450 133.540 ;
        RECT 118.730 132.900 118.870 135.810 ;
        RECT 118.250 132.760 118.870 132.900 ;
        RECT 118.250 127.990 118.390 132.760 ;
        RECT 118.190 127.670 118.450 127.990 ;
        RECT 111.950 126.930 112.210 127.250 ;
        RECT 112.010 125.030 112.150 126.930 ;
        RECT 111.950 124.710 112.210 125.030 ;
        RECT 114.830 124.340 115.090 124.660 ;
        RECT 112.910 123.230 113.170 123.550 ;
        RECT 111.950 116.570 112.210 116.890 ;
        RECT 111.470 103.250 111.730 103.570 ;
        RECT 110.990 100.290 111.250 100.610 ;
        RECT 109.550 94.740 109.810 95.060 ;
        RECT 111.050 92.840 111.190 100.290 ;
        RECT 110.990 92.520 111.250 92.840 ;
        RECT 108.110 91.410 108.370 91.730 ;
        RECT 110.510 91.040 110.770 91.360 ;
        RECT 110.570 87.660 110.710 91.040 ;
        RECT 110.510 87.340 110.770 87.660 ;
        RECT 107.630 84.380 107.890 84.700 ;
        RECT 112.010 84.330 112.150 116.570 ;
        RECT 112.970 111.710 113.110 123.230 ;
        RECT 114.890 121.330 115.030 124.340 ;
        RECT 114.830 121.010 115.090 121.330 ;
        RECT 118.250 115.040 118.390 127.670 ;
        RECT 118.670 126.930 118.930 127.250 ;
        RECT 118.730 125.400 118.870 126.930 ;
        RECT 118.670 125.080 118.930 125.400 ;
        RECT 124.430 116.200 124.690 116.520 ;
        RECT 117.230 114.720 117.490 115.040 ;
        RECT 118.190 114.720 118.450 115.040 ;
        RECT 112.910 111.390 113.170 111.710 ;
        RECT 117.290 111.340 117.430 114.720 ;
        RECT 117.230 111.020 117.490 111.340 ;
        RECT 118.250 109.120 118.390 114.720 ;
        RECT 124.490 113.190 124.630 116.200 ;
        RECT 124.430 112.870 124.690 113.190 ;
        RECT 113.870 108.800 114.130 109.120 ;
        RECT 118.190 108.800 118.450 109.120 ;
        RECT 113.930 100.240 114.070 108.800 ;
        RECT 123.950 108.430 124.210 108.750 ;
        RECT 117.710 106.580 117.970 106.900 ;
        RECT 117.770 104.310 117.910 106.580 ;
        RECT 117.710 103.990 117.970 104.310 ;
        RECT 117.230 103.620 117.490 103.940 ;
        RECT 113.870 99.920 114.130 100.240 ;
        RECT 116.750 99.180 117.010 99.500 ;
        RECT 116.810 96.910 116.950 99.180 ;
        RECT 117.290 99.130 117.430 103.620 ;
        RECT 117.230 98.810 117.490 99.130 ;
        RECT 117.290 96.910 117.430 98.810 ;
        RECT 116.750 96.590 117.010 96.910 ;
        RECT 117.230 96.590 117.490 96.910 ;
        RECT 117.770 92.100 117.910 103.990 ;
        RECT 118.190 99.920 118.450 100.240 ;
        RECT 117.710 91.780 117.970 92.100 ;
        RECT 118.250 88.770 118.390 99.920 ;
        RECT 124.010 99.870 124.150 108.430 ;
        RECT 125.390 103.620 125.650 103.940 ;
        RECT 124.910 102.880 125.170 103.200 ;
        RECT 123.950 99.550 124.210 99.870 ;
        RECT 123.950 95.480 124.210 95.800 ;
        RECT 124.010 92.470 124.150 95.480 ;
        RECT 123.950 92.150 124.210 92.470 ;
        RECT 124.970 91.730 125.110 102.880 ;
        RECT 125.450 100.240 125.590 103.620 ;
        RECT 125.390 99.920 125.650 100.240 ;
        RECT 132.110 94.740 132.370 95.060 ;
        RECT 124.910 91.410 125.170 91.730 ;
        RECT 120.590 90.670 120.850 90.990 ;
        RECT 118.190 88.450 118.450 88.770 ;
        RECT 120.650 87.290 120.790 90.670 ;
        RECT 120.590 86.970 120.850 87.290 ;
        RECT 113.390 86.230 113.650 86.550 ;
        RECT 113.450 84.700 113.590 86.230 ;
        RECT 113.390 84.380 113.650 84.700 ;
        RECT 111.950 84.010 112.210 84.330 ;
        RECT 114.830 84.010 115.090 84.330 ;
        RECT 114.890 80.630 115.030 84.010 ;
        RECT 114.830 80.310 115.090 80.630 ;
        RECT 116.270 80.310 116.530 80.630 ;
        RECT 104.270 79.570 104.530 79.890 ;
        RECT 102.350 78.460 102.610 78.780 ;
        RECT 101.390 75.870 101.650 76.190 ;
        RECT 98.990 75.130 99.250 75.450 ;
        RECT 100.430 75.130 100.690 75.450 ;
        RECT 93.710 72.170 93.970 72.490 ;
        RECT 100.490 72.330 100.630 75.130 ;
        RECT 102.410 75.080 102.550 78.460 ;
        RECT 104.330 76.190 104.470 79.570 ;
        RECT 116.330 79.520 116.470 80.310 ;
        RECT 116.270 79.200 116.530 79.520 ;
        RECT 107.150 78.460 107.410 78.780 ;
        RECT 104.270 75.870 104.530 76.190 ;
        RECT 102.350 74.760 102.610 75.080 ;
        RECT 100.420 71.960 100.700 72.330 ;
        RECT 102.350 72.170 102.610 72.490 ;
        RECT 101.390 71.060 101.650 71.380 ;
        RECT 99.950 70.690 100.210 71.010 ;
        RECT 98.510 70.320 98.770 70.640 ;
        RECT 93.230 69.950 93.490 70.270 ;
        RECT 97.550 68.100 97.810 68.420 ;
        RECT 94.670 67.360 94.930 67.680 ;
        RECT 92.750 66.620 93.010 66.940 ;
        RECT 90.830 55.890 91.090 56.210 ;
        RECT 87.950 54.410 88.210 54.730 ;
        RECT 90.350 54.410 90.610 54.730 ;
        RECT 87.470 54.040 87.730 54.360 ;
        RECT 87.530 45.850 87.670 54.040 ;
        RECT 87.470 45.530 87.730 45.850 ;
        RECT 86.990 38.500 87.250 38.820 ;
        RECT 85.070 38.130 85.330 38.450 ;
        RECT 81.230 34.430 81.490 34.750 ;
        RECT 86.510 34.430 86.770 34.750 ;
        RECT 79.790 31.470 80.050 31.790 ;
        RECT 80.750 30.150 81.010 30.310 ;
        RECT 80.740 29.780 81.020 30.150 ;
        RECT 78.830 23.330 79.090 23.650 ;
        RECT 81.290 23.280 81.430 34.430 ;
        RECT 86.570 33.640 86.710 34.430 ;
        RECT 86.510 33.320 86.770 33.640 ;
        RECT 82.670 30.360 82.930 30.680 ;
        RECT 83.630 30.360 83.890 30.680 ;
        RECT 82.730 26.240 82.870 30.360 ;
        RECT 83.690 30.150 83.830 30.360 ;
        RECT 83.620 29.780 83.900 30.150 ;
        RECT 82.670 25.920 82.930 26.240 ;
        RECT 81.230 22.960 81.490 23.280 ;
        RECT 83.690 21.430 83.830 29.780 ;
        RECT 86.030 29.250 86.290 29.570 ;
        RECT 83.630 21.110 83.890 21.430 ;
        RECT 86.090 19.580 86.230 29.250 ;
        RECT 86.570 26.980 86.710 33.320 ;
        RECT 86.510 26.660 86.770 26.980 ;
        RECT 87.050 25.500 87.190 38.500 ;
        RECT 86.990 25.180 87.250 25.500 ;
        RECT 87.050 23.650 87.190 25.180 ;
        RECT 86.990 23.330 87.250 23.650 ;
        RECT 87.530 23.280 87.670 45.530 ;
        RECT 88.010 43.260 88.150 54.410 ;
        RECT 90.410 51.770 90.550 54.410 ;
        RECT 90.350 51.450 90.610 51.770 ;
        RECT 94.190 49.600 94.450 49.920 ;
        RECT 89.870 46.640 90.130 46.960 ;
        RECT 87.950 42.940 88.210 43.260 ;
        RECT 89.930 39.560 90.070 46.640 ;
        RECT 91.790 45.900 92.050 46.220 ;
        RECT 91.850 42.890 91.990 45.900 ;
        RECT 94.250 43.260 94.390 49.600 ;
        RECT 94.190 42.940 94.450 43.260 ;
        RECT 91.790 42.570 92.050 42.890 ;
        RECT 94.730 42.520 94.870 67.360 ;
        RECT 95.150 66.620 95.410 66.940 ;
        RECT 95.210 63.240 95.350 66.620 ;
        RECT 95.150 62.920 95.410 63.240 ;
        RECT 95.210 59.170 95.350 62.920 ;
        RECT 95.150 58.850 95.410 59.170 ;
        RECT 95.210 51.030 95.350 58.850 ;
        RECT 97.610 56.210 97.750 68.100 ;
        RECT 98.030 62.180 98.290 62.500 ;
        RECT 97.550 55.890 97.810 56.210 ;
        RECT 98.090 54.730 98.230 62.180 ;
        RECT 98.570 62.130 98.710 70.320 ;
        RECT 99.470 62.550 99.730 62.870 ;
        RECT 98.510 61.810 98.770 62.130 ;
        RECT 98.030 54.410 98.290 54.730 ;
        RECT 98.030 53.670 98.290 53.990 ;
        RECT 95.150 50.710 95.410 51.030 ;
        RECT 97.550 47.380 97.810 47.700 ;
        RECT 97.610 46.220 97.750 47.380 ;
        RECT 97.550 45.900 97.810 46.220 ;
        RECT 95.150 45.530 95.410 45.850 ;
        RECT 95.210 42.890 95.350 45.530 ;
        RECT 97.610 44.100 97.750 45.900 ;
        RECT 96.590 43.680 96.850 44.000 ;
        RECT 97.130 43.960 97.750 44.100 ;
        RECT 98.090 44.000 98.230 53.670 ;
        RECT 95.150 42.570 95.410 42.890 ;
        RECT 94.670 42.200 94.930 42.520 ;
        RECT 96.650 41.780 96.790 43.680 ;
        RECT 96.590 41.460 96.850 41.780 ;
        RECT 97.130 39.560 97.270 43.960 ;
        RECT 98.030 43.680 98.290 44.000 ;
        RECT 97.550 42.940 97.810 43.260 ;
        RECT 97.610 42.620 97.750 42.940 ;
        RECT 97.610 42.480 98.230 42.620 ;
        RECT 89.870 39.240 90.130 39.560 ;
        RECT 95.150 39.240 95.410 39.560 ;
        RECT 97.070 39.240 97.330 39.560 ;
        RECT 94.670 35.030 94.930 35.120 ;
        RECT 93.770 34.890 94.930 35.030 ;
        RECT 93.770 29.940 93.910 34.890 ;
        RECT 94.670 34.800 94.930 34.890 ;
        RECT 95.210 31.790 95.350 39.240 ;
        RECT 97.550 38.870 97.810 39.190 ;
        RECT 95.150 31.470 95.410 31.790 ;
        RECT 94.190 30.360 94.450 30.680 ;
        RECT 93.710 29.620 93.970 29.940 ;
        RECT 93.770 26.240 93.910 29.620 ;
        RECT 93.710 25.920 93.970 26.240 ;
        RECT 94.250 23.650 94.390 30.360 ;
        RECT 95.210 30.310 95.350 31.470 ;
        RECT 97.610 31.050 97.750 38.870 ;
        RECT 98.090 38.820 98.230 42.480 ;
        RECT 98.030 38.500 98.290 38.820 ;
        RECT 98.090 31.420 98.230 38.500 ;
        RECT 98.570 35.860 98.710 61.810 ;
        RECT 99.530 54.360 99.670 62.550 ;
        RECT 99.470 54.040 99.730 54.360 ;
        RECT 98.990 46.270 99.250 46.590 ;
        RECT 99.050 42.890 99.190 46.270 ;
        RECT 98.990 42.570 99.250 42.890 ;
        RECT 99.050 39.190 99.190 42.570 ;
        RECT 99.530 39.560 99.670 54.040 ;
        RECT 100.010 53.990 100.150 70.690 ;
        RECT 100.910 65.880 101.170 66.200 ;
        RECT 100.970 64.350 101.110 65.880 ;
        RECT 100.910 64.030 101.170 64.350 ;
        RECT 100.430 62.550 100.690 62.870 ;
        RECT 99.950 53.670 100.210 53.990 ;
        RECT 99.950 51.080 100.210 51.400 ;
        RECT 99.470 39.240 99.730 39.560 ;
        RECT 98.990 38.870 99.250 39.190 ;
        RECT 99.470 37.390 99.730 37.710 ;
        RECT 98.510 35.540 98.770 35.860 ;
        RECT 98.990 34.430 99.250 34.750 ;
        RECT 98.030 31.100 98.290 31.420 ;
        RECT 97.550 30.730 97.810 31.050 ;
        RECT 99.050 30.310 99.190 34.430 ;
        RECT 95.150 30.150 95.410 30.310 ;
        RECT 95.140 29.780 95.420 30.150 ;
        RECT 98.990 29.990 99.250 30.310 ;
        RECT 99.530 29.940 99.670 37.390 ;
        RECT 99.470 29.620 99.730 29.940 ;
        RECT 96.110 27.030 96.370 27.350 ;
        RECT 94.670 26.290 94.930 26.610 ;
        RECT 94.190 23.330 94.450 23.650 ;
        RECT 87.470 22.960 87.730 23.280 ;
        RECT 94.730 22.540 94.870 26.290 ;
        RECT 94.670 22.220 94.930 22.540 ;
        RECT 96.170 22.170 96.310 27.030 ;
        RECT 97.550 26.660 97.810 26.980 ;
        RECT 97.610 22.910 97.750 26.660 ;
        RECT 99.530 26.610 99.670 29.620 ;
        RECT 99.470 26.290 99.730 26.610 ;
        RECT 97.550 22.590 97.810 22.910 ;
        RECT 96.110 21.850 96.370 22.170 ;
        RECT 94.190 21.110 94.450 21.430 ;
        RECT 86.030 19.260 86.290 19.580 ;
        RECT 94.250 19.210 94.390 21.110 ;
        RECT 97.610 19.580 97.750 22.590 ;
        RECT 100.010 21.800 100.150 51.080 ;
        RECT 100.490 46.960 100.630 62.550 ;
        RECT 100.970 55.100 101.110 64.030 ;
        RECT 100.910 54.780 101.170 55.100 ;
        RECT 100.970 51.770 101.110 54.780 ;
        RECT 100.910 51.450 101.170 51.770 ;
        RECT 101.450 47.330 101.590 71.060 ;
        RECT 101.870 70.690 102.130 71.010 ;
        RECT 101.930 59.170 102.070 70.690 ;
        RECT 101.870 58.850 102.130 59.170 ;
        RECT 101.390 47.010 101.650 47.330 ;
        RECT 100.430 46.640 100.690 46.960 ;
        RECT 100.910 45.530 101.170 45.850 ;
        RECT 100.430 43.310 100.690 43.630 ;
        RECT 100.490 39.930 100.630 43.310 ;
        RECT 100.430 39.610 100.690 39.930 ;
        RECT 100.490 34.750 100.630 39.610 ;
        RECT 100.970 38.450 101.110 45.530 ;
        RECT 101.450 39.190 101.590 47.010 ;
        RECT 102.410 46.590 102.550 72.170 ;
        RECT 106.660 71.960 106.940 72.330 ;
        RECT 106.670 71.800 106.930 71.960 ;
        RECT 103.310 71.430 103.570 71.750 ;
        RECT 105.710 71.480 105.970 71.750 ;
        RECT 105.710 71.430 106.870 71.480 ;
        RECT 102.830 70.690 103.090 71.010 ;
        RECT 102.890 68.050 103.030 70.690 ;
        RECT 102.830 67.730 103.090 68.050 ;
        RECT 103.370 46.590 103.510 71.430 ;
        RECT 105.770 71.340 106.870 71.430 ;
        RECT 106.730 70.270 106.870 71.340 ;
        RECT 106.670 69.950 106.930 70.270 ;
        RECT 107.210 68.050 107.350 78.460 ;
        RECT 108.110 78.090 108.370 78.410 ;
        RECT 114.830 78.090 115.090 78.410 ;
        RECT 119.150 78.090 119.410 78.410 ;
        RECT 108.170 75.820 108.310 78.090 ;
        RECT 114.890 76.560 115.030 78.090 ;
        RECT 119.210 76.560 119.350 78.090 ;
        RECT 114.830 76.240 115.090 76.560 ;
        RECT 119.150 76.240 119.410 76.560 ;
        RECT 108.110 75.500 108.370 75.820 ;
        RECT 110.030 75.500 110.290 75.820 ;
        RECT 116.750 75.500 117.010 75.820 ;
        RECT 108.590 71.060 108.850 71.380 ;
        RECT 108.650 68.420 108.790 71.060 ;
        RECT 108.590 68.100 108.850 68.420 ;
        RECT 107.150 67.730 107.410 68.050 ;
        RECT 107.150 61.810 107.410 62.130 ;
        RECT 107.210 60.280 107.350 61.810 ;
        RECT 107.150 59.960 107.410 60.280 ;
        RECT 105.230 59.220 105.490 59.540 ;
        RECT 102.350 46.270 102.610 46.590 ;
        RECT 103.310 46.270 103.570 46.590 ;
        RECT 101.870 45.900 102.130 46.220 ;
        RECT 101.390 38.870 101.650 39.190 ;
        RECT 100.910 38.130 101.170 38.450 ;
        RECT 101.390 37.760 101.650 38.080 ;
        RECT 100.430 34.430 100.690 34.750 ;
        RECT 100.910 30.360 101.170 30.680 ;
        RECT 100.970 21.800 101.110 30.360 ;
        RECT 101.450 22.170 101.590 37.760 ;
        RECT 101.930 31.050 102.070 45.900 ;
        RECT 102.410 38.820 102.550 46.270 ;
        RECT 103.370 41.780 103.510 46.270 ;
        RECT 103.790 41.830 104.050 42.150 ;
        RECT 103.310 41.460 103.570 41.780 ;
        RECT 102.350 38.500 102.610 38.820 ;
        RECT 103.370 35.860 103.510 41.460 ;
        RECT 103.310 35.540 103.570 35.860 ;
        RECT 101.870 30.730 102.130 31.050 ;
        RECT 103.370 29.940 103.510 35.540 ;
        RECT 103.850 33.640 103.990 41.830 ;
        RECT 103.790 33.320 104.050 33.640 ;
        RECT 103.310 29.620 103.570 29.940 ;
        RECT 103.370 27.720 103.510 29.620 ;
        RECT 103.310 27.400 103.570 27.720 ;
        RECT 103.850 26.980 103.990 33.320 ;
        RECT 103.790 26.660 104.050 26.980 ;
        RECT 103.790 22.960 104.050 23.280 ;
        RECT 103.850 22.170 103.990 22.960 ;
        RECT 101.390 21.850 101.650 22.170 ;
        RECT 103.790 21.850 104.050 22.170 ;
        RECT 105.290 21.800 105.430 59.220 ;
        RECT 108.590 54.780 108.850 55.100 ;
        RECT 108.650 51.400 108.790 54.780 ;
        RECT 110.090 54.730 110.230 75.500 ;
        RECT 116.810 75.080 116.950 75.500 ;
        RECT 116.270 74.760 116.530 75.080 ;
        RECT 116.750 74.760 117.010 75.080 ;
        RECT 113.390 71.060 113.650 71.380 ;
        RECT 112.910 70.690 113.170 71.010 ;
        RECT 110.990 68.100 111.250 68.420 ;
        RECT 110.030 54.410 110.290 54.730 ;
        RECT 108.590 51.080 108.850 51.400 ;
        RECT 106.190 42.570 106.450 42.890 ;
        RECT 106.250 34.380 106.390 42.570 ;
        RECT 108.110 38.130 108.370 38.450 ;
        RECT 106.670 35.170 106.930 35.490 ;
        RECT 106.190 34.060 106.450 34.380 ;
        RECT 105.710 31.100 105.970 31.420 ;
        RECT 105.770 30.310 105.910 31.100 ;
        RECT 105.710 30.150 105.970 30.310 ;
        RECT 105.700 29.780 105.980 30.150 ;
        RECT 105.710 29.250 105.970 29.570 ;
        RECT 99.950 21.480 100.210 21.800 ;
        RECT 100.910 21.480 101.170 21.800 ;
        RECT 105.230 21.480 105.490 21.800 ;
        RECT 105.770 19.580 105.910 29.250 ;
        RECT 97.550 19.260 97.810 19.580 ;
        RECT 105.710 19.260 105.970 19.580 ;
        RECT 94.190 18.890 94.450 19.210 ;
        RECT 77.870 18.520 78.130 18.840 ;
        RECT 68.750 18.240 69.430 18.380 ;
        RECT 68.750 18.150 69.010 18.240 ;
        RECT 69.710 18.150 69.970 18.470 ;
        RECT 106.250 17.730 106.390 34.060 ;
        RECT 106.730 33.640 106.870 35.170 ;
        RECT 106.670 33.320 106.930 33.640 ;
        RECT 108.170 30.680 108.310 38.130 ;
        RECT 108.110 30.360 108.370 30.680 ;
        RECT 106.660 29.780 106.940 30.150 ;
        RECT 106.730 27.720 106.870 29.780 ;
        RECT 106.670 27.400 106.930 27.720 ;
        RECT 108.650 26.980 108.790 51.080 ;
        RECT 110.510 50.710 110.770 51.030 ;
        RECT 110.570 43.630 110.710 50.710 ;
        RECT 110.510 43.310 110.770 43.630 ;
        RECT 111.050 34.750 111.190 68.100 ;
        RECT 111.950 66.250 112.210 66.570 ;
        RECT 112.010 35.860 112.150 66.250 ;
        RECT 112.970 62.500 113.110 70.690 ;
        RECT 113.450 68.420 113.590 71.060 ;
        RECT 115.790 70.690 116.050 71.010 ;
        RECT 113.390 68.100 113.650 68.420 ;
        RECT 115.310 67.360 115.570 67.680 ;
        RECT 112.910 62.180 113.170 62.500 ;
        RECT 115.370 59.170 115.510 67.360 ;
        RECT 115.310 58.850 115.570 59.170 ;
        RECT 112.430 46.640 112.690 46.960 ;
        RECT 112.490 38.820 112.630 46.640 ;
        RECT 115.850 39.770 115.990 70.690 ;
        RECT 116.330 51.770 116.470 74.760 ;
        RECT 120.650 71.010 120.790 86.970 ;
        RECT 130.670 79.570 130.930 79.890 ;
        RECT 123.470 78.090 123.730 78.410 ;
        RECT 123.530 76.190 123.670 78.090 ;
        RECT 123.470 75.870 123.730 76.190 ;
        RECT 130.730 72.120 130.870 79.570 ;
        RECT 130.670 71.800 130.930 72.120 ;
        RECT 120.590 70.690 120.850 71.010 ;
        RECT 117.230 69.950 117.490 70.270 ;
        RECT 118.190 69.950 118.450 70.270 ;
        RECT 117.290 67.680 117.430 69.950 ;
        RECT 117.230 67.360 117.490 67.680 ;
        RECT 116.750 66.990 117.010 67.310 ;
        RECT 116.810 54.360 116.950 66.990 ;
        RECT 118.250 62.500 118.390 69.950 ;
        RECT 130.730 68.420 130.870 71.800 ;
        RECT 130.670 68.100 130.930 68.420 ;
        RECT 129.710 66.250 129.970 66.570 ;
        RECT 124.910 65.880 125.170 66.200 ;
        RECT 129.230 65.880 129.490 66.200 ;
        RECT 118.190 62.180 118.450 62.500 ;
        RECT 121.550 59.590 121.810 59.910 ;
        RECT 117.230 59.220 117.490 59.540 ;
        RECT 120.590 59.220 120.850 59.540 ;
        RECT 116.750 54.040 117.010 54.360 ;
        RECT 116.270 51.450 116.530 51.770 ;
        RECT 117.290 46.960 117.430 59.220 ;
        RECT 118.190 58.480 118.450 58.800 ;
        RECT 118.250 55.200 118.390 58.480 ;
        RECT 117.710 54.780 117.970 55.100 ;
        RECT 118.250 55.060 118.870 55.200 ;
        RECT 117.230 46.640 117.490 46.960 ;
        RECT 117.770 46.220 117.910 54.780 ;
        RECT 118.190 54.040 118.450 54.360 ;
        RECT 118.250 51.030 118.390 54.040 ;
        RECT 118.190 50.710 118.450 51.030 ;
        RECT 118.730 50.020 118.870 55.060 ;
        RECT 118.250 49.880 118.870 50.020 ;
        RECT 117.710 45.900 117.970 46.220 ;
        RECT 115.780 39.400 116.060 39.770 ;
        RECT 112.430 38.500 112.690 38.820 ;
        RECT 111.950 35.540 112.210 35.860 ;
        RECT 118.250 35.120 118.390 49.880 ;
        RECT 120.650 42.890 120.790 59.220 ;
        RECT 121.070 54.780 121.330 55.100 ;
        RECT 121.130 43.260 121.270 54.780 ;
        RECT 121.070 42.940 121.330 43.260 ;
        RECT 121.610 42.890 121.750 59.590 ;
        RECT 123.470 59.220 123.730 59.540 ;
        RECT 122.510 58.850 122.770 59.170 ;
        RECT 122.570 54.730 122.710 58.850 ;
        RECT 123.530 55.470 123.670 59.220 ;
        RECT 123.470 55.150 123.730 55.470 ;
        RECT 122.510 54.410 122.770 54.730 ;
        RECT 120.590 42.570 120.850 42.890 ;
        RECT 121.550 42.570 121.810 42.890 ;
        RECT 124.970 39.930 125.110 65.880 ;
        RECT 129.290 55.100 129.430 65.880 ;
        RECT 129.230 54.780 129.490 55.100 ;
        RECT 128.270 51.080 128.530 51.400 ;
        RECT 129.230 51.080 129.490 51.400 ;
        RECT 126.350 50.710 126.610 51.030 ;
        RECT 127.310 50.710 127.570 51.030 ;
        RECT 124.910 39.610 125.170 39.930 ;
        RECT 124.430 38.500 124.690 38.820 ;
        RECT 123.470 38.130 123.730 38.450 ;
        RECT 122.990 37.760 123.250 38.080 ;
        RECT 118.190 34.800 118.450 35.120 ;
        RECT 110.030 34.430 110.290 34.750 ;
        RECT 110.990 34.430 111.250 34.750 ;
        RECT 108.590 26.660 108.850 26.980 ;
        RECT 110.090 25.870 110.230 34.430 ;
        RECT 118.190 33.690 118.450 34.010 ;
        RECT 120.590 33.690 120.850 34.010 ;
        RECT 110.990 33.320 111.250 33.640 ;
        RECT 111.950 33.320 112.210 33.640 ;
        RECT 111.050 31.050 111.190 33.320 ;
        RECT 110.990 30.730 111.250 31.050 ;
        RECT 111.470 29.620 111.730 29.940 ;
        RECT 111.530 27.720 111.670 29.620 ;
        RECT 111.470 27.400 111.730 27.720 ;
        RECT 112.010 27.350 112.150 33.320 ;
        RECT 115.310 29.620 115.570 29.940 ;
        RECT 116.750 29.620 117.010 29.940 ;
        RECT 111.950 27.030 112.210 27.350 ;
        RECT 115.370 26.610 115.510 29.620 ;
        RECT 116.810 26.610 116.950 29.620 ;
        RECT 117.710 29.250 117.970 29.570 ;
        RECT 115.310 26.290 115.570 26.610 ;
        RECT 116.750 26.290 117.010 26.610 ;
        RECT 110.030 25.550 110.290 25.870 ;
        RECT 115.370 22.910 115.510 26.290 ;
        RECT 115.310 22.590 115.570 22.910 ;
        RECT 116.810 22.540 116.950 26.290 ;
        RECT 117.770 23.650 117.910 29.250 ;
        RECT 118.250 27.350 118.390 33.690 ;
        RECT 118.190 27.030 118.450 27.350 ;
        RECT 118.190 26.290 118.450 26.610 ;
        RECT 117.710 23.330 117.970 23.650 ;
        RECT 118.250 22.540 118.390 26.290 ;
        RECT 120.650 22.540 120.790 33.690 ;
        RECT 122.510 33.320 122.770 33.640 ;
        RECT 121.070 31.100 121.330 31.420 ;
        RECT 121.130 30.310 121.270 31.100 ;
        RECT 121.070 30.150 121.330 30.310 ;
        RECT 121.060 29.780 121.340 30.150 ;
        RECT 122.570 26.980 122.710 33.320 ;
        RECT 123.050 30.680 123.190 37.760 ;
        RECT 123.530 35.860 123.670 38.130 ;
        RECT 124.490 35.860 124.630 38.500 ;
        RECT 126.410 35.860 126.550 50.710 ;
        RECT 127.370 43.260 127.510 50.710 ;
        RECT 128.330 46.590 128.470 51.080 ;
        RECT 128.270 46.270 128.530 46.590 ;
        RECT 127.310 42.940 127.570 43.260 ;
        RECT 127.790 42.940 128.050 43.260 ;
        RECT 123.470 35.540 123.730 35.860 ;
        RECT 124.430 35.540 124.690 35.860 ;
        RECT 126.350 35.540 126.610 35.860 ;
        RECT 124.910 35.170 125.170 35.490 ;
        RECT 122.990 30.360 123.250 30.680 ;
        RECT 123.470 29.990 123.730 30.310 ;
        RECT 123.530 26.980 123.670 29.990 ;
        RECT 124.970 27.720 125.110 35.170 ;
        RECT 127.850 34.750 127.990 42.940 ;
        RECT 129.290 38.820 129.430 51.080 ;
        RECT 129.770 39.930 129.910 66.250 ;
        RECT 130.190 58.850 130.450 59.170 ;
        RECT 130.250 54.730 130.390 58.850 ;
        RECT 130.190 54.410 130.450 54.730 ;
        RECT 129.710 39.610 129.970 39.930 ;
        RECT 129.230 38.500 129.490 38.820 ;
        RECT 129.770 35.860 129.910 39.610 ;
        RECT 130.730 39.560 130.870 68.100 ;
        RECT 132.170 67.680 132.310 94.740 ;
        RECT 137.390 74.760 137.650 75.080 ;
        RECT 133.070 70.320 133.330 70.640 ;
        RECT 132.110 67.360 132.370 67.680 ;
        RECT 133.130 55.940 133.270 70.320 ;
        RECT 134.990 69.950 135.250 70.270 ;
        RECT 135.050 62.500 135.190 69.950 ;
        RECT 135.950 67.730 136.210 68.050 ;
        RECT 134.990 62.180 135.250 62.500 ;
        RECT 133.130 55.800 133.750 55.940 ;
        RECT 133.070 54.780 133.330 55.100 ;
        RECT 133.130 51.770 133.270 54.780 ;
        RECT 133.070 51.450 133.330 51.770 ;
        RECT 133.610 42.890 133.750 55.800 ;
        RECT 136.010 55.470 136.150 67.730 ;
        RECT 136.910 61.810 137.170 62.130 ;
        RECT 136.970 56.210 137.110 61.810 ;
        RECT 136.910 55.890 137.170 56.210 ;
        RECT 135.950 55.150 136.210 55.470 ;
        RECT 136.010 51.030 136.150 55.150 ;
        RECT 137.450 54.730 137.590 74.760 ;
        RECT 138.350 67.360 138.610 67.680 ;
        RECT 138.410 64.350 138.550 67.360 ;
        RECT 139.310 66.990 139.570 67.310 ;
        RECT 138.350 64.030 138.610 64.350 ;
        RECT 137.870 54.780 138.130 55.100 ;
        RECT 137.390 54.410 137.650 54.730 ;
        RECT 135.950 50.710 136.210 51.030 ;
        RECT 133.550 42.570 133.810 42.890 ;
        RECT 130.670 39.240 130.930 39.560 ;
        RECT 129.710 35.540 129.970 35.860 ;
        RECT 127.790 34.430 128.050 34.750 ;
        RECT 127.310 29.620 127.570 29.940 ;
        RECT 125.390 29.250 125.650 29.570 ;
        RECT 124.910 27.400 125.170 27.720 ;
        RECT 122.510 26.660 122.770 26.980 ;
        RECT 123.470 26.660 123.730 26.980 ;
        RECT 116.750 22.220 117.010 22.540 ;
        RECT 118.190 22.220 118.450 22.540 ;
        RECT 120.590 22.220 120.850 22.540 ;
        RECT 109.070 21.110 109.330 21.430 ;
        RECT 109.130 19.210 109.270 21.110 ;
        RECT 118.250 19.580 118.390 22.220 ;
        RECT 125.450 22.170 125.590 29.250 ;
        RECT 127.370 27.350 127.510 29.620 ;
        RECT 127.310 27.030 127.570 27.350 ;
        RECT 130.730 26.980 130.870 39.240 ;
        RECT 136.010 38.820 136.150 50.710 ;
        RECT 136.430 45.900 136.690 46.220 ;
        RECT 136.490 39.930 136.630 45.900 ;
        RECT 136.910 45.530 137.170 45.850 ;
        RECT 136.430 39.610 136.690 39.930 ;
        RECT 136.430 38.870 136.690 39.190 ;
        RECT 135.950 38.500 136.210 38.820 ;
        RECT 136.490 35.860 136.630 38.870 ;
        RECT 136.430 35.540 136.690 35.860 ;
        RECT 136.970 35.120 137.110 45.530 ;
        RECT 136.910 34.800 137.170 35.120 ;
        RECT 137.930 31.420 138.070 54.780 ;
        RECT 139.370 51.400 139.510 66.990 ;
        RECT 139.310 51.080 139.570 51.400 ;
        RECT 138.350 50.340 138.610 50.660 ;
        RECT 138.410 43.630 138.550 50.340 ;
        RECT 138.350 43.310 138.610 43.630 ;
        RECT 138.350 41.460 138.610 41.780 ;
        RECT 138.410 39.190 138.550 41.460 ;
        RECT 138.350 38.870 138.610 39.190 ;
        RECT 137.870 31.100 138.130 31.420 ;
        RECT 136.910 29.990 137.170 30.310 ;
        RECT 130.670 26.660 130.930 26.980 ;
        RECT 129.230 25.180 129.490 25.500 ;
        RECT 129.290 22.910 129.430 25.180 ;
        RECT 130.730 23.280 130.870 26.660 ;
        RECT 136.970 23.650 137.110 29.990 ;
        RECT 136.910 23.330 137.170 23.650 ;
        RECT 130.670 22.960 130.930 23.280 ;
        RECT 129.230 22.590 129.490 22.910 ;
        RECT 125.390 21.850 125.650 22.170 ;
        RECT 118.190 19.260 118.450 19.580 ;
        RECT 109.070 18.890 109.330 19.210 ;
        RECT 66.830 17.410 67.090 17.730 ;
        RECT 106.190 17.410 106.450 17.730 ;
        RECT 64.490 16.580 65.110 16.720 ;
        RECT 64.490 15.880 64.630 16.580 ;
        RECT 41.870 15.560 42.130 15.880 ;
        RECT 64.430 15.560 64.690 15.880 ;
      LAYER via2 ;
        RECT 21.220 69.790 21.500 70.070 ;
        RECT 14.020 62.390 14.300 62.670 ;
        RECT 6.820 54.250 7.100 54.530 ;
        RECT 21.700 50.550 21.980 50.830 ;
        RECT 21.220 42.410 21.500 42.690 ;
        RECT 23.140 54.250 23.420 54.530 ;
        RECT 31.300 69.790 31.580 70.070 ;
        RECT 22.180 39.450 22.460 39.730 ;
        RECT 25.060 42.410 25.340 42.690 ;
        RECT 24.100 39.450 24.380 39.730 ;
        RECT 36.580 50.550 36.860 50.830 ;
        RECT 39.460 62.390 39.740 62.670 ;
        RECT 35.140 42.410 35.420 42.690 ;
        RECT 55.300 96.430 55.580 96.710 ;
        RECT 86.980 96.430 87.260 96.710 ;
        RECT 62.500 29.830 62.780 30.110 ;
        RECT 69.220 29.830 69.500 30.110 ;
        RECT 100.420 72.010 100.700 72.290 ;
        RECT 80.740 29.830 81.020 30.110 ;
        RECT 83.620 29.830 83.900 30.110 ;
        RECT 95.140 29.830 95.420 30.110 ;
        RECT 106.660 72.010 106.940 72.290 ;
        RECT 105.700 29.830 105.980 30.110 ;
        RECT 106.660 29.830 106.940 30.110 ;
        RECT 115.780 39.450 116.060 39.730 ;
        RECT 121.060 29.830 121.340 30.110 ;
      LAYER met3 ;
        RECT 55.270 96.720 55.600 96.730 ;
        RECT 86.950 96.720 87.280 96.730 ;
        RECT 55.270 96.420 87.280 96.720 ;
        RECT 55.270 96.400 55.600 96.420 ;
        RECT 86.950 96.400 87.280 96.420 ;
        RECT 100.390 72.300 100.720 72.310 ;
        RECT 106.630 72.300 106.960 72.310 ;
        RECT 100.390 72.000 106.960 72.300 ;
        RECT 100.390 71.980 100.720 72.000 ;
        RECT 106.630 71.980 106.960 72.000 ;
        RECT 21.190 70.080 21.520 70.090 ;
        RECT 31.270 70.080 31.600 70.090 ;
        RECT 21.190 69.780 31.600 70.080 ;
        RECT 21.190 69.760 21.520 69.780 ;
        RECT 31.270 69.760 31.600 69.780 ;
        RECT 13.990 62.680 14.320 62.690 ;
        RECT 39.430 62.680 39.760 62.690 ;
        RECT 13.990 62.380 39.760 62.680 ;
        RECT 13.990 62.360 14.320 62.380 ;
        RECT 39.430 62.360 39.760 62.380 ;
        RECT 6.790 54.540 7.120 54.550 ;
        RECT 23.110 54.540 23.440 54.550 ;
        RECT 6.790 54.240 23.440 54.540 ;
        RECT 6.790 54.220 7.120 54.240 ;
        RECT 23.110 54.220 23.440 54.240 ;
        RECT 21.670 50.840 22.000 50.850 ;
        RECT 36.550 50.840 36.880 50.850 ;
        RECT 21.670 50.540 36.880 50.840 ;
        RECT 21.670 50.520 22.000 50.540 ;
        RECT 36.550 50.520 36.880 50.540 ;
        RECT 21.190 42.700 21.520 42.710 ;
        RECT 25.030 42.700 25.360 42.710 ;
        RECT 35.110 42.700 35.440 42.710 ;
        RECT 21.190 42.400 35.440 42.700 ;
        RECT 21.190 42.380 21.520 42.400 ;
        RECT 25.030 42.380 25.360 42.400 ;
        RECT 35.110 42.380 35.440 42.400 ;
        RECT 22.150 39.740 22.480 39.750 ;
        RECT 24.070 39.740 24.400 39.750 ;
        RECT 115.750 39.740 116.080 39.750 ;
        RECT 22.150 39.440 116.080 39.740 ;
        RECT 22.150 39.420 22.480 39.440 ;
        RECT 24.070 39.420 24.400 39.440 ;
        RECT 115.750 39.420 116.080 39.440 ;
        RECT 62.470 30.120 62.800 30.130 ;
        RECT 69.190 30.120 69.520 30.130 ;
        RECT 80.710 30.120 81.040 30.130 ;
        RECT 62.470 29.820 81.040 30.120 ;
        RECT 62.470 29.800 62.800 29.820 ;
        RECT 69.190 29.800 69.520 29.820 ;
        RECT 80.710 29.800 81.040 29.820 ;
        RECT 83.590 30.120 83.920 30.130 ;
        RECT 95.110 30.120 95.440 30.130 ;
        RECT 83.590 29.820 95.440 30.120 ;
        RECT 83.590 29.800 83.920 29.820 ;
        RECT 95.110 29.800 95.440 29.820 ;
        RECT 105.670 30.120 106.000 30.130 ;
        RECT 106.630 30.120 106.960 30.130 ;
        RECT 121.030 30.120 121.360 30.130 ;
        RECT 105.670 29.820 121.360 30.120 ;
        RECT 105.670 29.800 106.000 29.820 ;
        RECT 106.630 29.800 106.960 29.820 ;
        RECT 121.030 29.800 121.360 29.820 ;
  END
END raven_spi
END LIBRARY

